module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module fs(input [0:0] a, input [0:0] b, input [0:0] bin, output [0:0] fs_xor1, output [0:0] fs_or0);
  wire [0:0] fs_xor0;
  wire [0:0] fs_not0;
  wire [0:0] fs_and0;
  wire [0:0] fs_not1;
  wire [0:0] fs_and1;
  xor_gate xor_gate_fs_xor0(.a(a[0]), .b(b[0]), .out(fs_xor0));
  not_gate not_gate_fs_not0(.a(a[0]), .out(fs_not0));
  and_gate and_gate_fs_and0(.a(fs_not0[0]), .b(b[0]), .out(fs_and0));
  xor_gate xor_gate_fs_xor1(.a(bin[0]), .b(fs_xor0[0]), .out(fs_xor1));
  not_gate not_gate_fs_not1(.a(fs_xor0[0]), .out(fs_not1));
  and_gate and_gate_fs_and1(.a(fs_not1[0]), .b(bin[0]), .out(fs_and1));
  or_gate or_gate_fs_or0(.a(fs_and1[0]), .b(fs_and0[0]), .out(fs_or0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module arrdiv32(input [31:0] a, input [31:0] b, output [31:0] arrdiv32_out);
  wire [0:0] arrdiv32_fs0_xor0;
  wire [0:0] arrdiv32_fs0_and0;
  wire [0:0] arrdiv32_fs1_xor1;
  wire [0:0] arrdiv32_fs1_or0;
  wire [0:0] arrdiv32_fs2_xor1;
  wire [0:0] arrdiv32_fs2_or0;
  wire [0:0] arrdiv32_fs3_xor1;
  wire [0:0] arrdiv32_fs3_or0;
  wire [0:0] arrdiv32_fs4_xor1;
  wire [0:0] arrdiv32_fs4_or0;
  wire [0:0] arrdiv32_fs5_xor1;
  wire [0:0] arrdiv32_fs5_or0;
  wire [0:0] arrdiv32_fs6_xor1;
  wire [0:0] arrdiv32_fs6_or0;
  wire [0:0] arrdiv32_fs7_xor1;
  wire [0:0] arrdiv32_fs7_or0;
  wire [0:0] arrdiv32_fs8_xor1;
  wire [0:0] arrdiv32_fs8_or0;
  wire [0:0] arrdiv32_fs9_xor1;
  wire [0:0] arrdiv32_fs9_or0;
  wire [0:0] arrdiv32_fs10_xor1;
  wire [0:0] arrdiv32_fs10_or0;
  wire [0:0] arrdiv32_fs11_xor1;
  wire [0:0] arrdiv32_fs11_or0;
  wire [0:0] arrdiv32_fs12_xor1;
  wire [0:0] arrdiv32_fs12_or0;
  wire [0:0] arrdiv32_fs13_xor1;
  wire [0:0] arrdiv32_fs13_or0;
  wire [0:0] arrdiv32_fs14_xor1;
  wire [0:0] arrdiv32_fs14_or0;
  wire [0:0] arrdiv32_fs15_xor1;
  wire [0:0] arrdiv32_fs15_or0;
  wire [0:0] arrdiv32_fs16_xor1;
  wire [0:0] arrdiv32_fs16_or0;
  wire [0:0] arrdiv32_fs17_xor1;
  wire [0:0] arrdiv32_fs17_or0;
  wire [0:0] arrdiv32_fs18_xor1;
  wire [0:0] arrdiv32_fs18_or0;
  wire [0:0] arrdiv32_fs19_xor1;
  wire [0:0] arrdiv32_fs19_or0;
  wire [0:0] arrdiv32_fs20_xor1;
  wire [0:0] arrdiv32_fs20_or0;
  wire [0:0] arrdiv32_fs21_xor1;
  wire [0:0] arrdiv32_fs21_or0;
  wire [0:0] arrdiv32_fs22_xor1;
  wire [0:0] arrdiv32_fs22_or0;
  wire [0:0] arrdiv32_fs23_xor1;
  wire [0:0] arrdiv32_fs23_or0;
  wire [0:0] arrdiv32_fs24_xor1;
  wire [0:0] arrdiv32_fs24_or0;
  wire [0:0] arrdiv32_fs25_xor1;
  wire [0:0] arrdiv32_fs25_or0;
  wire [0:0] arrdiv32_fs26_xor1;
  wire [0:0] arrdiv32_fs26_or0;
  wire [0:0] arrdiv32_fs27_xor1;
  wire [0:0] arrdiv32_fs27_or0;
  wire [0:0] arrdiv32_fs28_xor1;
  wire [0:0] arrdiv32_fs28_or0;
  wire [0:0] arrdiv32_fs29_xor1;
  wire [0:0] arrdiv32_fs29_or0;
  wire [0:0] arrdiv32_fs30_xor1;
  wire [0:0] arrdiv32_fs30_or0;
  wire [0:0] arrdiv32_fs31_xor1;
  wire [0:0] arrdiv32_fs31_or0;
  wire [0:0] arrdiv32_mux2to10_xor0;
  wire [0:0] arrdiv32_mux2to11_and1;
  wire [0:0] arrdiv32_mux2to12_and1;
  wire [0:0] arrdiv32_mux2to13_and1;
  wire [0:0] arrdiv32_mux2to14_and1;
  wire [0:0] arrdiv32_mux2to15_and1;
  wire [0:0] arrdiv32_mux2to16_and1;
  wire [0:0] arrdiv32_mux2to17_and1;
  wire [0:0] arrdiv32_mux2to18_and1;
  wire [0:0] arrdiv32_mux2to19_and1;
  wire [0:0] arrdiv32_mux2to110_and1;
  wire [0:0] arrdiv32_mux2to111_and1;
  wire [0:0] arrdiv32_mux2to112_and1;
  wire [0:0] arrdiv32_mux2to113_and1;
  wire [0:0] arrdiv32_mux2to114_and1;
  wire [0:0] arrdiv32_mux2to115_and1;
  wire [0:0] arrdiv32_mux2to116_and1;
  wire [0:0] arrdiv32_mux2to117_and1;
  wire [0:0] arrdiv32_mux2to118_and1;
  wire [0:0] arrdiv32_mux2to119_and1;
  wire [0:0] arrdiv32_mux2to120_and1;
  wire [0:0] arrdiv32_mux2to121_and1;
  wire [0:0] arrdiv32_mux2to122_and1;
  wire [0:0] arrdiv32_mux2to123_and1;
  wire [0:0] arrdiv32_mux2to124_and1;
  wire [0:0] arrdiv32_mux2to125_and1;
  wire [0:0] arrdiv32_mux2to126_and1;
  wire [0:0] arrdiv32_mux2to127_and1;
  wire [0:0] arrdiv32_mux2to128_and1;
  wire [0:0] arrdiv32_mux2to129_and1;
  wire [0:0] arrdiv32_mux2to130_and1;
  wire [0:0] arrdiv32_not0;
  wire [0:0] arrdiv32_fs32_xor0;
  wire [0:0] arrdiv32_fs32_and0;
  wire [0:0] arrdiv32_fs33_xor1;
  wire [0:0] arrdiv32_fs33_or0;
  wire [0:0] arrdiv32_fs34_xor1;
  wire [0:0] arrdiv32_fs34_or0;
  wire [0:0] arrdiv32_fs35_xor1;
  wire [0:0] arrdiv32_fs35_or0;
  wire [0:0] arrdiv32_fs36_xor1;
  wire [0:0] arrdiv32_fs36_or0;
  wire [0:0] arrdiv32_fs37_xor1;
  wire [0:0] arrdiv32_fs37_or0;
  wire [0:0] arrdiv32_fs38_xor1;
  wire [0:0] arrdiv32_fs38_or0;
  wire [0:0] arrdiv32_fs39_xor1;
  wire [0:0] arrdiv32_fs39_or0;
  wire [0:0] arrdiv32_fs40_xor1;
  wire [0:0] arrdiv32_fs40_or0;
  wire [0:0] arrdiv32_fs41_xor1;
  wire [0:0] arrdiv32_fs41_or0;
  wire [0:0] arrdiv32_fs42_xor1;
  wire [0:0] arrdiv32_fs42_or0;
  wire [0:0] arrdiv32_fs43_xor1;
  wire [0:0] arrdiv32_fs43_or0;
  wire [0:0] arrdiv32_fs44_xor1;
  wire [0:0] arrdiv32_fs44_or0;
  wire [0:0] arrdiv32_fs45_xor1;
  wire [0:0] arrdiv32_fs45_or0;
  wire [0:0] arrdiv32_fs46_xor1;
  wire [0:0] arrdiv32_fs46_or0;
  wire [0:0] arrdiv32_fs47_xor1;
  wire [0:0] arrdiv32_fs47_or0;
  wire [0:0] arrdiv32_fs48_xor1;
  wire [0:0] arrdiv32_fs48_or0;
  wire [0:0] arrdiv32_fs49_xor1;
  wire [0:0] arrdiv32_fs49_or0;
  wire [0:0] arrdiv32_fs50_xor1;
  wire [0:0] arrdiv32_fs50_or0;
  wire [0:0] arrdiv32_fs51_xor1;
  wire [0:0] arrdiv32_fs51_or0;
  wire [0:0] arrdiv32_fs52_xor1;
  wire [0:0] arrdiv32_fs52_or0;
  wire [0:0] arrdiv32_fs53_xor1;
  wire [0:0] arrdiv32_fs53_or0;
  wire [0:0] arrdiv32_fs54_xor1;
  wire [0:0] arrdiv32_fs54_or0;
  wire [0:0] arrdiv32_fs55_xor1;
  wire [0:0] arrdiv32_fs55_or0;
  wire [0:0] arrdiv32_fs56_xor1;
  wire [0:0] arrdiv32_fs56_or0;
  wire [0:0] arrdiv32_fs57_xor1;
  wire [0:0] arrdiv32_fs57_or0;
  wire [0:0] arrdiv32_fs58_xor1;
  wire [0:0] arrdiv32_fs58_or0;
  wire [0:0] arrdiv32_fs59_xor1;
  wire [0:0] arrdiv32_fs59_or0;
  wire [0:0] arrdiv32_fs60_xor1;
  wire [0:0] arrdiv32_fs60_or0;
  wire [0:0] arrdiv32_fs61_xor1;
  wire [0:0] arrdiv32_fs61_or0;
  wire [0:0] arrdiv32_fs62_xor1;
  wire [0:0] arrdiv32_fs62_or0;
  wire [0:0] arrdiv32_fs63_xor1;
  wire [0:0] arrdiv32_fs63_or0;
  wire [0:0] arrdiv32_mux2to131_xor0;
  wire [0:0] arrdiv32_mux2to132_xor0;
  wire [0:0] arrdiv32_mux2to133_xor0;
  wire [0:0] arrdiv32_mux2to134_xor0;
  wire [0:0] arrdiv32_mux2to135_xor0;
  wire [0:0] arrdiv32_mux2to136_xor0;
  wire [0:0] arrdiv32_mux2to137_xor0;
  wire [0:0] arrdiv32_mux2to138_xor0;
  wire [0:0] arrdiv32_mux2to139_xor0;
  wire [0:0] arrdiv32_mux2to140_xor0;
  wire [0:0] arrdiv32_mux2to141_xor0;
  wire [0:0] arrdiv32_mux2to142_xor0;
  wire [0:0] arrdiv32_mux2to143_xor0;
  wire [0:0] arrdiv32_mux2to144_xor0;
  wire [0:0] arrdiv32_mux2to145_xor0;
  wire [0:0] arrdiv32_mux2to146_xor0;
  wire [0:0] arrdiv32_mux2to147_xor0;
  wire [0:0] arrdiv32_mux2to148_xor0;
  wire [0:0] arrdiv32_mux2to149_xor0;
  wire [0:0] arrdiv32_mux2to150_xor0;
  wire [0:0] arrdiv32_mux2to151_xor0;
  wire [0:0] arrdiv32_mux2to152_xor0;
  wire [0:0] arrdiv32_mux2to153_xor0;
  wire [0:0] arrdiv32_mux2to154_xor0;
  wire [0:0] arrdiv32_mux2to155_xor0;
  wire [0:0] arrdiv32_mux2to156_xor0;
  wire [0:0] arrdiv32_mux2to157_xor0;
  wire [0:0] arrdiv32_mux2to158_xor0;
  wire [0:0] arrdiv32_mux2to159_xor0;
  wire [0:0] arrdiv32_mux2to160_xor0;
  wire [0:0] arrdiv32_mux2to161_xor0;
  wire [0:0] arrdiv32_not1;
  wire [0:0] arrdiv32_fs64_xor0;
  wire [0:0] arrdiv32_fs64_and0;
  wire [0:0] arrdiv32_fs65_xor1;
  wire [0:0] arrdiv32_fs65_or0;
  wire [0:0] arrdiv32_fs66_xor1;
  wire [0:0] arrdiv32_fs66_or0;
  wire [0:0] arrdiv32_fs67_xor1;
  wire [0:0] arrdiv32_fs67_or0;
  wire [0:0] arrdiv32_fs68_xor1;
  wire [0:0] arrdiv32_fs68_or0;
  wire [0:0] arrdiv32_fs69_xor1;
  wire [0:0] arrdiv32_fs69_or0;
  wire [0:0] arrdiv32_fs70_xor1;
  wire [0:0] arrdiv32_fs70_or0;
  wire [0:0] arrdiv32_fs71_xor1;
  wire [0:0] arrdiv32_fs71_or0;
  wire [0:0] arrdiv32_fs72_xor1;
  wire [0:0] arrdiv32_fs72_or0;
  wire [0:0] arrdiv32_fs73_xor1;
  wire [0:0] arrdiv32_fs73_or0;
  wire [0:0] arrdiv32_fs74_xor1;
  wire [0:0] arrdiv32_fs74_or0;
  wire [0:0] arrdiv32_fs75_xor1;
  wire [0:0] arrdiv32_fs75_or0;
  wire [0:0] arrdiv32_fs76_xor1;
  wire [0:0] arrdiv32_fs76_or0;
  wire [0:0] arrdiv32_fs77_xor1;
  wire [0:0] arrdiv32_fs77_or0;
  wire [0:0] arrdiv32_fs78_xor1;
  wire [0:0] arrdiv32_fs78_or0;
  wire [0:0] arrdiv32_fs79_xor1;
  wire [0:0] arrdiv32_fs79_or0;
  wire [0:0] arrdiv32_fs80_xor1;
  wire [0:0] arrdiv32_fs80_or0;
  wire [0:0] arrdiv32_fs81_xor1;
  wire [0:0] arrdiv32_fs81_or0;
  wire [0:0] arrdiv32_fs82_xor1;
  wire [0:0] arrdiv32_fs82_or0;
  wire [0:0] arrdiv32_fs83_xor1;
  wire [0:0] arrdiv32_fs83_or0;
  wire [0:0] arrdiv32_fs84_xor1;
  wire [0:0] arrdiv32_fs84_or0;
  wire [0:0] arrdiv32_fs85_xor1;
  wire [0:0] arrdiv32_fs85_or0;
  wire [0:0] arrdiv32_fs86_xor1;
  wire [0:0] arrdiv32_fs86_or0;
  wire [0:0] arrdiv32_fs87_xor1;
  wire [0:0] arrdiv32_fs87_or0;
  wire [0:0] arrdiv32_fs88_xor1;
  wire [0:0] arrdiv32_fs88_or0;
  wire [0:0] arrdiv32_fs89_xor1;
  wire [0:0] arrdiv32_fs89_or0;
  wire [0:0] arrdiv32_fs90_xor1;
  wire [0:0] arrdiv32_fs90_or0;
  wire [0:0] arrdiv32_fs91_xor1;
  wire [0:0] arrdiv32_fs91_or0;
  wire [0:0] arrdiv32_fs92_xor1;
  wire [0:0] arrdiv32_fs92_or0;
  wire [0:0] arrdiv32_fs93_xor1;
  wire [0:0] arrdiv32_fs93_or0;
  wire [0:0] arrdiv32_fs94_xor1;
  wire [0:0] arrdiv32_fs94_or0;
  wire [0:0] arrdiv32_fs95_xor1;
  wire [0:0] arrdiv32_fs95_or0;
  wire [0:0] arrdiv32_mux2to162_xor0;
  wire [0:0] arrdiv32_mux2to163_xor0;
  wire [0:0] arrdiv32_mux2to164_xor0;
  wire [0:0] arrdiv32_mux2to165_xor0;
  wire [0:0] arrdiv32_mux2to166_xor0;
  wire [0:0] arrdiv32_mux2to167_xor0;
  wire [0:0] arrdiv32_mux2to168_xor0;
  wire [0:0] arrdiv32_mux2to169_xor0;
  wire [0:0] arrdiv32_mux2to170_xor0;
  wire [0:0] arrdiv32_mux2to171_xor0;
  wire [0:0] arrdiv32_mux2to172_xor0;
  wire [0:0] arrdiv32_mux2to173_xor0;
  wire [0:0] arrdiv32_mux2to174_xor0;
  wire [0:0] arrdiv32_mux2to175_xor0;
  wire [0:0] arrdiv32_mux2to176_xor0;
  wire [0:0] arrdiv32_mux2to177_xor0;
  wire [0:0] arrdiv32_mux2to178_xor0;
  wire [0:0] arrdiv32_mux2to179_xor0;
  wire [0:0] arrdiv32_mux2to180_xor0;
  wire [0:0] arrdiv32_mux2to181_xor0;
  wire [0:0] arrdiv32_mux2to182_xor0;
  wire [0:0] arrdiv32_mux2to183_xor0;
  wire [0:0] arrdiv32_mux2to184_xor0;
  wire [0:0] arrdiv32_mux2to185_xor0;
  wire [0:0] arrdiv32_mux2to186_xor0;
  wire [0:0] arrdiv32_mux2to187_xor0;
  wire [0:0] arrdiv32_mux2to188_xor0;
  wire [0:0] arrdiv32_mux2to189_xor0;
  wire [0:0] arrdiv32_mux2to190_xor0;
  wire [0:0] arrdiv32_mux2to191_xor0;
  wire [0:0] arrdiv32_mux2to192_xor0;
  wire [0:0] arrdiv32_not2;
  wire [0:0] arrdiv32_fs96_xor0;
  wire [0:0] arrdiv32_fs96_and0;
  wire [0:0] arrdiv32_fs97_xor1;
  wire [0:0] arrdiv32_fs97_or0;
  wire [0:0] arrdiv32_fs98_xor1;
  wire [0:0] arrdiv32_fs98_or0;
  wire [0:0] arrdiv32_fs99_xor1;
  wire [0:0] arrdiv32_fs99_or0;
  wire [0:0] arrdiv32_fs100_xor1;
  wire [0:0] arrdiv32_fs100_or0;
  wire [0:0] arrdiv32_fs101_xor1;
  wire [0:0] arrdiv32_fs101_or0;
  wire [0:0] arrdiv32_fs102_xor1;
  wire [0:0] arrdiv32_fs102_or0;
  wire [0:0] arrdiv32_fs103_xor1;
  wire [0:0] arrdiv32_fs103_or0;
  wire [0:0] arrdiv32_fs104_xor1;
  wire [0:0] arrdiv32_fs104_or0;
  wire [0:0] arrdiv32_fs105_xor1;
  wire [0:0] arrdiv32_fs105_or0;
  wire [0:0] arrdiv32_fs106_xor1;
  wire [0:0] arrdiv32_fs106_or0;
  wire [0:0] arrdiv32_fs107_xor1;
  wire [0:0] arrdiv32_fs107_or0;
  wire [0:0] arrdiv32_fs108_xor1;
  wire [0:0] arrdiv32_fs108_or0;
  wire [0:0] arrdiv32_fs109_xor1;
  wire [0:0] arrdiv32_fs109_or0;
  wire [0:0] arrdiv32_fs110_xor1;
  wire [0:0] arrdiv32_fs110_or0;
  wire [0:0] arrdiv32_fs111_xor1;
  wire [0:0] arrdiv32_fs111_or0;
  wire [0:0] arrdiv32_fs112_xor1;
  wire [0:0] arrdiv32_fs112_or0;
  wire [0:0] arrdiv32_fs113_xor1;
  wire [0:0] arrdiv32_fs113_or0;
  wire [0:0] arrdiv32_fs114_xor1;
  wire [0:0] arrdiv32_fs114_or0;
  wire [0:0] arrdiv32_fs115_xor1;
  wire [0:0] arrdiv32_fs115_or0;
  wire [0:0] arrdiv32_fs116_xor1;
  wire [0:0] arrdiv32_fs116_or0;
  wire [0:0] arrdiv32_fs117_xor1;
  wire [0:0] arrdiv32_fs117_or0;
  wire [0:0] arrdiv32_fs118_xor1;
  wire [0:0] arrdiv32_fs118_or0;
  wire [0:0] arrdiv32_fs119_xor1;
  wire [0:0] arrdiv32_fs119_or0;
  wire [0:0] arrdiv32_fs120_xor1;
  wire [0:0] arrdiv32_fs120_or0;
  wire [0:0] arrdiv32_fs121_xor1;
  wire [0:0] arrdiv32_fs121_or0;
  wire [0:0] arrdiv32_fs122_xor1;
  wire [0:0] arrdiv32_fs122_or0;
  wire [0:0] arrdiv32_fs123_xor1;
  wire [0:0] arrdiv32_fs123_or0;
  wire [0:0] arrdiv32_fs124_xor1;
  wire [0:0] arrdiv32_fs124_or0;
  wire [0:0] arrdiv32_fs125_xor1;
  wire [0:0] arrdiv32_fs125_or0;
  wire [0:0] arrdiv32_fs126_xor1;
  wire [0:0] arrdiv32_fs126_or0;
  wire [0:0] arrdiv32_fs127_xor1;
  wire [0:0] arrdiv32_fs127_or0;
  wire [0:0] arrdiv32_mux2to193_xor0;
  wire [0:0] arrdiv32_mux2to194_xor0;
  wire [0:0] arrdiv32_mux2to195_xor0;
  wire [0:0] arrdiv32_mux2to196_xor0;
  wire [0:0] arrdiv32_mux2to197_xor0;
  wire [0:0] arrdiv32_mux2to198_xor0;
  wire [0:0] arrdiv32_mux2to199_xor0;
  wire [0:0] arrdiv32_mux2to1100_xor0;
  wire [0:0] arrdiv32_mux2to1101_xor0;
  wire [0:0] arrdiv32_mux2to1102_xor0;
  wire [0:0] arrdiv32_mux2to1103_xor0;
  wire [0:0] arrdiv32_mux2to1104_xor0;
  wire [0:0] arrdiv32_mux2to1105_xor0;
  wire [0:0] arrdiv32_mux2to1106_xor0;
  wire [0:0] arrdiv32_mux2to1107_xor0;
  wire [0:0] arrdiv32_mux2to1108_xor0;
  wire [0:0] arrdiv32_mux2to1109_xor0;
  wire [0:0] arrdiv32_mux2to1110_xor0;
  wire [0:0] arrdiv32_mux2to1111_xor0;
  wire [0:0] arrdiv32_mux2to1112_xor0;
  wire [0:0] arrdiv32_mux2to1113_xor0;
  wire [0:0] arrdiv32_mux2to1114_xor0;
  wire [0:0] arrdiv32_mux2to1115_xor0;
  wire [0:0] arrdiv32_mux2to1116_xor0;
  wire [0:0] arrdiv32_mux2to1117_xor0;
  wire [0:0] arrdiv32_mux2to1118_xor0;
  wire [0:0] arrdiv32_mux2to1119_xor0;
  wire [0:0] arrdiv32_mux2to1120_xor0;
  wire [0:0] arrdiv32_mux2to1121_xor0;
  wire [0:0] arrdiv32_mux2to1122_xor0;
  wire [0:0] arrdiv32_mux2to1123_xor0;
  wire [0:0] arrdiv32_not3;
  wire [0:0] arrdiv32_fs128_xor0;
  wire [0:0] arrdiv32_fs128_and0;
  wire [0:0] arrdiv32_fs129_xor1;
  wire [0:0] arrdiv32_fs129_or0;
  wire [0:0] arrdiv32_fs130_xor1;
  wire [0:0] arrdiv32_fs130_or0;
  wire [0:0] arrdiv32_fs131_xor1;
  wire [0:0] arrdiv32_fs131_or0;
  wire [0:0] arrdiv32_fs132_xor1;
  wire [0:0] arrdiv32_fs132_or0;
  wire [0:0] arrdiv32_fs133_xor1;
  wire [0:0] arrdiv32_fs133_or0;
  wire [0:0] arrdiv32_fs134_xor1;
  wire [0:0] arrdiv32_fs134_or0;
  wire [0:0] arrdiv32_fs135_xor1;
  wire [0:0] arrdiv32_fs135_or0;
  wire [0:0] arrdiv32_fs136_xor1;
  wire [0:0] arrdiv32_fs136_or0;
  wire [0:0] arrdiv32_fs137_xor1;
  wire [0:0] arrdiv32_fs137_or0;
  wire [0:0] arrdiv32_fs138_xor1;
  wire [0:0] arrdiv32_fs138_or0;
  wire [0:0] arrdiv32_fs139_xor1;
  wire [0:0] arrdiv32_fs139_or0;
  wire [0:0] arrdiv32_fs140_xor1;
  wire [0:0] arrdiv32_fs140_or0;
  wire [0:0] arrdiv32_fs141_xor1;
  wire [0:0] arrdiv32_fs141_or0;
  wire [0:0] arrdiv32_fs142_xor1;
  wire [0:0] arrdiv32_fs142_or0;
  wire [0:0] arrdiv32_fs143_xor1;
  wire [0:0] arrdiv32_fs143_or0;
  wire [0:0] arrdiv32_fs144_xor1;
  wire [0:0] arrdiv32_fs144_or0;
  wire [0:0] arrdiv32_fs145_xor1;
  wire [0:0] arrdiv32_fs145_or0;
  wire [0:0] arrdiv32_fs146_xor1;
  wire [0:0] arrdiv32_fs146_or0;
  wire [0:0] arrdiv32_fs147_xor1;
  wire [0:0] arrdiv32_fs147_or0;
  wire [0:0] arrdiv32_fs148_xor1;
  wire [0:0] arrdiv32_fs148_or0;
  wire [0:0] arrdiv32_fs149_xor1;
  wire [0:0] arrdiv32_fs149_or0;
  wire [0:0] arrdiv32_fs150_xor1;
  wire [0:0] arrdiv32_fs150_or0;
  wire [0:0] arrdiv32_fs151_xor1;
  wire [0:0] arrdiv32_fs151_or0;
  wire [0:0] arrdiv32_fs152_xor1;
  wire [0:0] arrdiv32_fs152_or0;
  wire [0:0] arrdiv32_fs153_xor1;
  wire [0:0] arrdiv32_fs153_or0;
  wire [0:0] arrdiv32_fs154_xor1;
  wire [0:0] arrdiv32_fs154_or0;
  wire [0:0] arrdiv32_fs155_xor1;
  wire [0:0] arrdiv32_fs155_or0;
  wire [0:0] arrdiv32_fs156_xor1;
  wire [0:0] arrdiv32_fs156_or0;
  wire [0:0] arrdiv32_fs157_xor1;
  wire [0:0] arrdiv32_fs157_or0;
  wire [0:0] arrdiv32_fs158_xor1;
  wire [0:0] arrdiv32_fs158_or0;
  wire [0:0] arrdiv32_fs159_xor1;
  wire [0:0] arrdiv32_fs159_or0;
  wire [0:0] arrdiv32_mux2to1124_xor0;
  wire [0:0] arrdiv32_mux2to1125_xor0;
  wire [0:0] arrdiv32_mux2to1126_xor0;
  wire [0:0] arrdiv32_mux2to1127_xor0;
  wire [0:0] arrdiv32_mux2to1128_xor0;
  wire [0:0] arrdiv32_mux2to1129_xor0;
  wire [0:0] arrdiv32_mux2to1130_xor0;
  wire [0:0] arrdiv32_mux2to1131_xor0;
  wire [0:0] arrdiv32_mux2to1132_xor0;
  wire [0:0] arrdiv32_mux2to1133_xor0;
  wire [0:0] arrdiv32_mux2to1134_xor0;
  wire [0:0] arrdiv32_mux2to1135_xor0;
  wire [0:0] arrdiv32_mux2to1136_xor0;
  wire [0:0] arrdiv32_mux2to1137_xor0;
  wire [0:0] arrdiv32_mux2to1138_xor0;
  wire [0:0] arrdiv32_mux2to1139_xor0;
  wire [0:0] arrdiv32_mux2to1140_xor0;
  wire [0:0] arrdiv32_mux2to1141_xor0;
  wire [0:0] arrdiv32_mux2to1142_xor0;
  wire [0:0] arrdiv32_mux2to1143_xor0;
  wire [0:0] arrdiv32_mux2to1144_xor0;
  wire [0:0] arrdiv32_mux2to1145_xor0;
  wire [0:0] arrdiv32_mux2to1146_xor0;
  wire [0:0] arrdiv32_mux2to1147_xor0;
  wire [0:0] arrdiv32_mux2to1148_xor0;
  wire [0:0] arrdiv32_mux2to1149_xor0;
  wire [0:0] arrdiv32_mux2to1150_xor0;
  wire [0:0] arrdiv32_mux2to1151_xor0;
  wire [0:0] arrdiv32_mux2to1152_xor0;
  wire [0:0] arrdiv32_mux2to1153_xor0;
  wire [0:0] arrdiv32_mux2to1154_xor0;
  wire [0:0] arrdiv32_not4;
  wire [0:0] arrdiv32_fs160_xor0;
  wire [0:0] arrdiv32_fs160_and0;
  wire [0:0] arrdiv32_fs161_xor1;
  wire [0:0] arrdiv32_fs161_or0;
  wire [0:0] arrdiv32_fs162_xor1;
  wire [0:0] arrdiv32_fs162_or0;
  wire [0:0] arrdiv32_fs163_xor1;
  wire [0:0] arrdiv32_fs163_or0;
  wire [0:0] arrdiv32_fs164_xor1;
  wire [0:0] arrdiv32_fs164_or0;
  wire [0:0] arrdiv32_fs165_xor1;
  wire [0:0] arrdiv32_fs165_or0;
  wire [0:0] arrdiv32_fs166_xor1;
  wire [0:0] arrdiv32_fs166_or0;
  wire [0:0] arrdiv32_fs167_xor1;
  wire [0:0] arrdiv32_fs167_or0;
  wire [0:0] arrdiv32_fs168_xor1;
  wire [0:0] arrdiv32_fs168_or0;
  wire [0:0] arrdiv32_fs169_xor1;
  wire [0:0] arrdiv32_fs169_or0;
  wire [0:0] arrdiv32_fs170_xor1;
  wire [0:0] arrdiv32_fs170_or0;
  wire [0:0] arrdiv32_fs171_xor1;
  wire [0:0] arrdiv32_fs171_or0;
  wire [0:0] arrdiv32_fs172_xor1;
  wire [0:0] arrdiv32_fs172_or0;
  wire [0:0] arrdiv32_fs173_xor1;
  wire [0:0] arrdiv32_fs173_or0;
  wire [0:0] arrdiv32_fs174_xor1;
  wire [0:0] arrdiv32_fs174_or0;
  wire [0:0] arrdiv32_fs175_xor1;
  wire [0:0] arrdiv32_fs175_or0;
  wire [0:0] arrdiv32_fs176_xor1;
  wire [0:0] arrdiv32_fs176_or0;
  wire [0:0] arrdiv32_fs177_xor1;
  wire [0:0] arrdiv32_fs177_or0;
  wire [0:0] arrdiv32_fs178_xor1;
  wire [0:0] arrdiv32_fs178_or0;
  wire [0:0] arrdiv32_fs179_xor1;
  wire [0:0] arrdiv32_fs179_or0;
  wire [0:0] arrdiv32_fs180_xor1;
  wire [0:0] arrdiv32_fs180_or0;
  wire [0:0] arrdiv32_fs181_xor1;
  wire [0:0] arrdiv32_fs181_or0;
  wire [0:0] arrdiv32_fs182_xor1;
  wire [0:0] arrdiv32_fs182_or0;
  wire [0:0] arrdiv32_fs183_xor1;
  wire [0:0] arrdiv32_fs183_or0;
  wire [0:0] arrdiv32_fs184_xor1;
  wire [0:0] arrdiv32_fs184_or0;
  wire [0:0] arrdiv32_fs185_xor1;
  wire [0:0] arrdiv32_fs185_or0;
  wire [0:0] arrdiv32_fs186_xor1;
  wire [0:0] arrdiv32_fs186_or0;
  wire [0:0] arrdiv32_fs187_xor1;
  wire [0:0] arrdiv32_fs187_or0;
  wire [0:0] arrdiv32_fs188_xor1;
  wire [0:0] arrdiv32_fs188_or0;
  wire [0:0] arrdiv32_fs189_xor1;
  wire [0:0] arrdiv32_fs189_or0;
  wire [0:0] arrdiv32_fs190_xor1;
  wire [0:0] arrdiv32_fs190_or0;
  wire [0:0] arrdiv32_fs191_xor1;
  wire [0:0] arrdiv32_fs191_or0;
  wire [0:0] arrdiv32_mux2to1155_xor0;
  wire [0:0] arrdiv32_mux2to1156_xor0;
  wire [0:0] arrdiv32_mux2to1157_xor0;
  wire [0:0] arrdiv32_mux2to1158_xor0;
  wire [0:0] arrdiv32_mux2to1159_xor0;
  wire [0:0] arrdiv32_mux2to1160_xor0;
  wire [0:0] arrdiv32_mux2to1161_xor0;
  wire [0:0] arrdiv32_mux2to1162_xor0;
  wire [0:0] arrdiv32_mux2to1163_xor0;
  wire [0:0] arrdiv32_mux2to1164_xor0;
  wire [0:0] arrdiv32_mux2to1165_xor0;
  wire [0:0] arrdiv32_mux2to1166_xor0;
  wire [0:0] arrdiv32_mux2to1167_xor0;
  wire [0:0] arrdiv32_mux2to1168_xor0;
  wire [0:0] arrdiv32_mux2to1169_xor0;
  wire [0:0] arrdiv32_mux2to1170_xor0;
  wire [0:0] arrdiv32_mux2to1171_xor0;
  wire [0:0] arrdiv32_mux2to1172_xor0;
  wire [0:0] arrdiv32_mux2to1173_xor0;
  wire [0:0] arrdiv32_mux2to1174_xor0;
  wire [0:0] arrdiv32_mux2to1175_xor0;
  wire [0:0] arrdiv32_mux2to1176_xor0;
  wire [0:0] arrdiv32_mux2to1177_xor0;
  wire [0:0] arrdiv32_mux2to1178_xor0;
  wire [0:0] arrdiv32_mux2to1179_xor0;
  wire [0:0] arrdiv32_mux2to1180_xor0;
  wire [0:0] arrdiv32_mux2to1181_xor0;
  wire [0:0] arrdiv32_mux2to1182_xor0;
  wire [0:0] arrdiv32_mux2to1183_xor0;
  wire [0:0] arrdiv32_mux2to1184_xor0;
  wire [0:0] arrdiv32_mux2to1185_xor0;
  wire [0:0] arrdiv32_not5;
  wire [0:0] arrdiv32_fs192_xor0;
  wire [0:0] arrdiv32_fs192_and0;
  wire [0:0] arrdiv32_fs193_xor1;
  wire [0:0] arrdiv32_fs193_or0;
  wire [0:0] arrdiv32_fs194_xor1;
  wire [0:0] arrdiv32_fs194_or0;
  wire [0:0] arrdiv32_fs195_xor1;
  wire [0:0] arrdiv32_fs195_or0;
  wire [0:0] arrdiv32_fs196_xor1;
  wire [0:0] arrdiv32_fs196_or0;
  wire [0:0] arrdiv32_fs197_xor1;
  wire [0:0] arrdiv32_fs197_or0;
  wire [0:0] arrdiv32_fs198_xor1;
  wire [0:0] arrdiv32_fs198_or0;
  wire [0:0] arrdiv32_fs199_xor1;
  wire [0:0] arrdiv32_fs199_or0;
  wire [0:0] arrdiv32_fs200_xor1;
  wire [0:0] arrdiv32_fs200_or0;
  wire [0:0] arrdiv32_fs201_xor1;
  wire [0:0] arrdiv32_fs201_or0;
  wire [0:0] arrdiv32_fs202_xor1;
  wire [0:0] arrdiv32_fs202_or0;
  wire [0:0] arrdiv32_fs203_xor1;
  wire [0:0] arrdiv32_fs203_or0;
  wire [0:0] arrdiv32_fs204_xor1;
  wire [0:0] arrdiv32_fs204_or0;
  wire [0:0] arrdiv32_fs205_xor1;
  wire [0:0] arrdiv32_fs205_or0;
  wire [0:0] arrdiv32_fs206_xor1;
  wire [0:0] arrdiv32_fs206_or0;
  wire [0:0] arrdiv32_fs207_xor1;
  wire [0:0] arrdiv32_fs207_or0;
  wire [0:0] arrdiv32_fs208_xor1;
  wire [0:0] arrdiv32_fs208_or0;
  wire [0:0] arrdiv32_fs209_xor1;
  wire [0:0] arrdiv32_fs209_or0;
  wire [0:0] arrdiv32_fs210_xor1;
  wire [0:0] arrdiv32_fs210_or0;
  wire [0:0] arrdiv32_fs211_xor1;
  wire [0:0] arrdiv32_fs211_or0;
  wire [0:0] arrdiv32_fs212_xor1;
  wire [0:0] arrdiv32_fs212_or0;
  wire [0:0] arrdiv32_fs213_xor1;
  wire [0:0] arrdiv32_fs213_or0;
  wire [0:0] arrdiv32_fs214_xor1;
  wire [0:0] arrdiv32_fs214_or0;
  wire [0:0] arrdiv32_fs215_xor1;
  wire [0:0] arrdiv32_fs215_or0;
  wire [0:0] arrdiv32_fs216_xor1;
  wire [0:0] arrdiv32_fs216_or0;
  wire [0:0] arrdiv32_fs217_xor1;
  wire [0:0] arrdiv32_fs217_or0;
  wire [0:0] arrdiv32_fs218_xor1;
  wire [0:0] arrdiv32_fs218_or0;
  wire [0:0] arrdiv32_fs219_xor1;
  wire [0:0] arrdiv32_fs219_or0;
  wire [0:0] arrdiv32_fs220_xor1;
  wire [0:0] arrdiv32_fs220_or0;
  wire [0:0] arrdiv32_fs221_xor1;
  wire [0:0] arrdiv32_fs221_or0;
  wire [0:0] arrdiv32_fs222_xor1;
  wire [0:0] arrdiv32_fs222_or0;
  wire [0:0] arrdiv32_fs223_xor1;
  wire [0:0] arrdiv32_fs223_or0;
  wire [0:0] arrdiv32_mux2to1186_xor0;
  wire [0:0] arrdiv32_mux2to1187_xor0;
  wire [0:0] arrdiv32_mux2to1188_xor0;
  wire [0:0] arrdiv32_mux2to1189_xor0;
  wire [0:0] arrdiv32_mux2to1190_xor0;
  wire [0:0] arrdiv32_mux2to1191_xor0;
  wire [0:0] arrdiv32_mux2to1192_xor0;
  wire [0:0] arrdiv32_mux2to1193_xor0;
  wire [0:0] arrdiv32_mux2to1194_xor0;
  wire [0:0] arrdiv32_mux2to1195_xor0;
  wire [0:0] arrdiv32_mux2to1196_xor0;
  wire [0:0] arrdiv32_mux2to1197_xor0;
  wire [0:0] arrdiv32_mux2to1198_xor0;
  wire [0:0] arrdiv32_mux2to1199_xor0;
  wire [0:0] arrdiv32_mux2to1200_xor0;
  wire [0:0] arrdiv32_mux2to1201_xor0;
  wire [0:0] arrdiv32_mux2to1202_xor0;
  wire [0:0] arrdiv32_mux2to1203_xor0;
  wire [0:0] arrdiv32_mux2to1204_xor0;
  wire [0:0] arrdiv32_mux2to1205_xor0;
  wire [0:0] arrdiv32_mux2to1206_xor0;
  wire [0:0] arrdiv32_mux2to1207_xor0;
  wire [0:0] arrdiv32_mux2to1208_xor0;
  wire [0:0] arrdiv32_mux2to1209_xor0;
  wire [0:0] arrdiv32_mux2to1210_xor0;
  wire [0:0] arrdiv32_mux2to1211_xor0;
  wire [0:0] arrdiv32_mux2to1212_xor0;
  wire [0:0] arrdiv32_mux2to1213_xor0;
  wire [0:0] arrdiv32_mux2to1214_xor0;
  wire [0:0] arrdiv32_mux2to1215_xor0;
  wire [0:0] arrdiv32_mux2to1216_xor0;
  wire [0:0] arrdiv32_not6;
  wire [0:0] arrdiv32_fs224_xor0;
  wire [0:0] arrdiv32_fs224_and0;
  wire [0:0] arrdiv32_fs225_xor1;
  wire [0:0] arrdiv32_fs225_or0;
  wire [0:0] arrdiv32_fs226_xor1;
  wire [0:0] arrdiv32_fs226_or0;
  wire [0:0] arrdiv32_fs227_xor1;
  wire [0:0] arrdiv32_fs227_or0;
  wire [0:0] arrdiv32_fs228_xor1;
  wire [0:0] arrdiv32_fs228_or0;
  wire [0:0] arrdiv32_fs229_xor1;
  wire [0:0] arrdiv32_fs229_or0;
  wire [0:0] arrdiv32_fs230_xor1;
  wire [0:0] arrdiv32_fs230_or0;
  wire [0:0] arrdiv32_fs231_xor1;
  wire [0:0] arrdiv32_fs231_or0;
  wire [0:0] arrdiv32_fs232_xor1;
  wire [0:0] arrdiv32_fs232_or0;
  wire [0:0] arrdiv32_fs233_xor1;
  wire [0:0] arrdiv32_fs233_or0;
  wire [0:0] arrdiv32_fs234_xor1;
  wire [0:0] arrdiv32_fs234_or0;
  wire [0:0] arrdiv32_fs235_xor1;
  wire [0:0] arrdiv32_fs235_or0;
  wire [0:0] arrdiv32_fs236_xor1;
  wire [0:0] arrdiv32_fs236_or0;
  wire [0:0] arrdiv32_fs237_xor1;
  wire [0:0] arrdiv32_fs237_or0;
  wire [0:0] arrdiv32_fs238_xor1;
  wire [0:0] arrdiv32_fs238_or0;
  wire [0:0] arrdiv32_fs239_xor1;
  wire [0:0] arrdiv32_fs239_or0;
  wire [0:0] arrdiv32_fs240_xor1;
  wire [0:0] arrdiv32_fs240_or0;
  wire [0:0] arrdiv32_fs241_xor1;
  wire [0:0] arrdiv32_fs241_or0;
  wire [0:0] arrdiv32_fs242_xor1;
  wire [0:0] arrdiv32_fs242_or0;
  wire [0:0] arrdiv32_fs243_xor1;
  wire [0:0] arrdiv32_fs243_or0;
  wire [0:0] arrdiv32_fs244_xor1;
  wire [0:0] arrdiv32_fs244_or0;
  wire [0:0] arrdiv32_fs245_xor1;
  wire [0:0] arrdiv32_fs245_or0;
  wire [0:0] arrdiv32_fs246_xor1;
  wire [0:0] arrdiv32_fs246_or0;
  wire [0:0] arrdiv32_fs247_xor1;
  wire [0:0] arrdiv32_fs247_or0;
  wire [0:0] arrdiv32_fs248_xor1;
  wire [0:0] arrdiv32_fs248_or0;
  wire [0:0] arrdiv32_fs249_xor1;
  wire [0:0] arrdiv32_fs249_or0;
  wire [0:0] arrdiv32_fs250_xor1;
  wire [0:0] arrdiv32_fs250_or0;
  wire [0:0] arrdiv32_fs251_xor1;
  wire [0:0] arrdiv32_fs251_or0;
  wire [0:0] arrdiv32_fs252_xor1;
  wire [0:0] arrdiv32_fs252_or0;
  wire [0:0] arrdiv32_fs253_xor1;
  wire [0:0] arrdiv32_fs253_or0;
  wire [0:0] arrdiv32_fs254_xor1;
  wire [0:0] arrdiv32_fs254_or0;
  wire [0:0] arrdiv32_fs255_xor1;
  wire [0:0] arrdiv32_fs255_or0;
  wire [0:0] arrdiv32_mux2to1217_xor0;
  wire [0:0] arrdiv32_mux2to1218_xor0;
  wire [0:0] arrdiv32_mux2to1219_xor0;
  wire [0:0] arrdiv32_mux2to1220_xor0;
  wire [0:0] arrdiv32_mux2to1221_xor0;
  wire [0:0] arrdiv32_mux2to1222_xor0;
  wire [0:0] arrdiv32_mux2to1223_xor0;
  wire [0:0] arrdiv32_mux2to1224_xor0;
  wire [0:0] arrdiv32_mux2to1225_xor0;
  wire [0:0] arrdiv32_mux2to1226_xor0;
  wire [0:0] arrdiv32_mux2to1227_xor0;
  wire [0:0] arrdiv32_mux2to1228_xor0;
  wire [0:0] arrdiv32_mux2to1229_xor0;
  wire [0:0] arrdiv32_mux2to1230_xor0;
  wire [0:0] arrdiv32_mux2to1231_xor0;
  wire [0:0] arrdiv32_mux2to1232_xor0;
  wire [0:0] arrdiv32_mux2to1233_xor0;
  wire [0:0] arrdiv32_mux2to1234_xor0;
  wire [0:0] arrdiv32_mux2to1235_xor0;
  wire [0:0] arrdiv32_mux2to1236_xor0;
  wire [0:0] arrdiv32_mux2to1237_xor0;
  wire [0:0] arrdiv32_mux2to1238_xor0;
  wire [0:0] arrdiv32_mux2to1239_xor0;
  wire [0:0] arrdiv32_mux2to1240_xor0;
  wire [0:0] arrdiv32_mux2to1241_xor0;
  wire [0:0] arrdiv32_mux2to1242_xor0;
  wire [0:0] arrdiv32_mux2to1243_xor0;
  wire [0:0] arrdiv32_mux2to1244_xor0;
  wire [0:0] arrdiv32_mux2to1245_xor0;
  wire [0:0] arrdiv32_mux2to1246_xor0;
  wire [0:0] arrdiv32_mux2to1247_xor0;
  wire [0:0] arrdiv32_not7;
  wire [0:0] arrdiv32_fs256_xor0;
  wire [0:0] arrdiv32_fs256_and0;
  wire [0:0] arrdiv32_fs257_xor1;
  wire [0:0] arrdiv32_fs257_or0;
  wire [0:0] arrdiv32_fs258_xor1;
  wire [0:0] arrdiv32_fs258_or0;
  wire [0:0] arrdiv32_fs259_xor1;
  wire [0:0] arrdiv32_fs259_or0;
  wire [0:0] arrdiv32_fs260_xor1;
  wire [0:0] arrdiv32_fs260_or0;
  wire [0:0] arrdiv32_fs261_xor1;
  wire [0:0] arrdiv32_fs261_or0;
  wire [0:0] arrdiv32_fs262_xor1;
  wire [0:0] arrdiv32_fs262_or0;
  wire [0:0] arrdiv32_fs263_xor1;
  wire [0:0] arrdiv32_fs263_or0;
  wire [0:0] arrdiv32_fs264_xor1;
  wire [0:0] arrdiv32_fs264_or0;
  wire [0:0] arrdiv32_fs265_xor1;
  wire [0:0] arrdiv32_fs265_or0;
  wire [0:0] arrdiv32_fs266_xor1;
  wire [0:0] arrdiv32_fs266_or0;
  wire [0:0] arrdiv32_fs267_xor1;
  wire [0:0] arrdiv32_fs267_or0;
  wire [0:0] arrdiv32_fs268_xor1;
  wire [0:0] arrdiv32_fs268_or0;
  wire [0:0] arrdiv32_fs269_xor1;
  wire [0:0] arrdiv32_fs269_or0;
  wire [0:0] arrdiv32_fs270_xor1;
  wire [0:0] arrdiv32_fs270_or0;
  wire [0:0] arrdiv32_fs271_xor1;
  wire [0:0] arrdiv32_fs271_or0;
  wire [0:0] arrdiv32_fs272_xor1;
  wire [0:0] arrdiv32_fs272_or0;
  wire [0:0] arrdiv32_fs273_xor1;
  wire [0:0] arrdiv32_fs273_or0;
  wire [0:0] arrdiv32_fs274_xor1;
  wire [0:0] arrdiv32_fs274_or0;
  wire [0:0] arrdiv32_fs275_xor1;
  wire [0:0] arrdiv32_fs275_or0;
  wire [0:0] arrdiv32_fs276_xor1;
  wire [0:0] arrdiv32_fs276_or0;
  wire [0:0] arrdiv32_fs277_xor1;
  wire [0:0] arrdiv32_fs277_or0;
  wire [0:0] arrdiv32_fs278_xor1;
  wire [0:0] arrdiv32_fs278_or0;
  wire [0:0] arrdiv32_fs279_xor1;
  wire [0:0] arrdiv32_fs279_or0;
  wire [0:0] arrdiv32_fs280_xor1;
  wire [0:0] arrdiv32_fs280_or0;
  wire [0:0] arrdiv32_fs281_xor1;
  wire [0:0] arrdiv32_fs281_or0;
  wire [0:0] arrdiv32_fs282_xor1;
  wire [0:0] arrdiv32_fs282_or0;
  wire [0:0] arrdiv32_fs283_xor1;
  wire [0:0] arrdiv32_fs283_or0;
  wire [0:0] arrdiv32_fs284_xor1;
  wire [0:0] arrdiv32_fs284_or0;
  wire [0:0] arrdiv32_fs285_xor1;
  wire [0:0] arrdiv32_fs285_or0;
  wire [0:0] arrdiv32_fs286_xor1;
  wire [0:0] arrdiv32_fs286_or0;
  wire [0:0] arrdiv32_fs287_xor1;
  wire [0:0] arrdiv32_fs287_or0;
  wire [0:0] arrdiv32_mux2to1248_xor0;
  wire [0:0] arrdiv32_mux2to1249_xor0;
  wire [0:0] arrdiv32_mux2to1250_xor0;
  wire [0:0] arrdiv32_mux2to1251_xor0;
  wire [0:0] arrdiv32_mux2to1252_xor0;
  wire [0:0] arrdiv32_mux2to1253_xor0;
  wire [0:0] arrdiv32_mux2to1254_xor0;
  wire [0:0] arrdiv32_mux2to1255_xor0;
  wire [0:0] arrdiv32_mux2to1256_xor0;
  wire [0:0] arrdiv32_mux2to1257_xor0;
  wire [0:0] arrdiv32_mux2to1258_xor0;
  wire [0:0] arrdiv32_mux2to1259_xor0;
  wire [0:0] arrdiv32_mux2to1260_xor0;
  wire [0:0] arrdiv32_mux2to1261_xor0;
  wire [0:0] arrdiv32_mux2to1262_xor0;
  wire [0:0] arrdiv32_mux2to1263_xor0;
  wire [0:0] arrdiv32_mux2to1264_xor0;
  wire [0:0] arrdiv32_mux2to1265_xor0;
  wire [0:0] arrdiv32_mux2to1266_xor0;
  wire [0:0] arrdiv32_mux2to1267_xor0;
  wire [0:0] arrdiv32_mux2to1268_xor0;
  wire [0:0] arrdiv32_mux2to1269_xor0;
  wire [0:0] arrdiv32_mux2to1270_xor0;
  wire [0:0] arrdiv32_mux2to1271_xor0;
  wire [0:0] arrdiv32_mux2to1272_xor0;
  wire [0:0] arrdiv32_mux2to1273_xor0;
  wire [0:0] arrdiv32_mux2to1274_xor0;
  wire [0:0] arrdiv32_mux2to1275_xor0;
  wire [0:0] arrdiv32_mux2to1276_xor0;
  wire [0:0] arrdiv32_mux2to1277_xor0;
  wire [0:0] arrdiv32_mux2to1278_xor0;
  wire [0:0] arrdiv32_not8;
  wire [0:0] arrdiv32_fs288_xor0;
  wire [0:0] arrdiv32_fs288_and0;
  wire [0:0] arrdiv32_fs289_xor1;
  wire [0:0] arrdiv32_fs289_or0;
  wire [0:0] arrdiv32_fs290_xor1;
  wire [0:0] arrdiv32_fs290_or0;
  wire [0:0] arrdiv32_fs291_xor1;
  wire [0:0] arrdiv32_fs291_or0;
  wire [0:0] arrdiv32_fs292_xor1;
  wire [0:0] arrdiv32_fs292_or0;
  wire [0:0] arrdiv32_fs293_xor1;
  wire [0:0] arrdiv32_fs293_or0;
  wire [0:0] arrdiv32_fs294_xor1;
  wire [0:0] arrdiv32_fs294_or0;
  wire [0:0] arrdiv32_fs295_xor1;
  wire [0:0] arrdiv32_fs295_or0;
  wire [0:0] arrdiv32_fs296_xor1;
  wire [0:0] arrdiv32_fs296_or0;
  wire [0:0] arrdiv32_fs297_xor1;
  wire [0:0] arrdiv32_fs297_or0;
  wire [0:0] arrdiv32_fs298_xor1;
  wire [0:0] arrdiv32_fs298_or0;
  wire [0:0] arrdiv32_fs299_xor1;
  wire [0:0] arrdiv32_fs299_or0;
  wire [0:0] arrdiv32_fs300_xor1;
  wire [0:0] arrdiv32_fs300_or0;
  wire [0:0] arrdiv32_fs301_xor1;
  wire [0:0] arrdiv32_fs301_or0;
  wire [0:0] arrdiv32_fs302_xor1;
  wire [0:0] arrdiv32_fs302_or0;
  wire [0:0] arrdiv32_fs303_xor1;
  wire [0:0] arrdiv32_fs303_or0;
  wire [0:0] arrdiv32_fs304_xor1;
  wire [0:0] arrdiv32_fs304_or0;
  wire [0:0] arrdiv32_fs305_xor1;
  wire [0:0] arrdiv32_fs305_or0;
  wire [0:0] arrdiv32_fs306_xor1;
  wire [0:0] arrdiv32_fs306_or0;
  wire [0:0] arrdiv32_fs307_xor1;
  wire [0:0] arrdiv32_fs307_or0;
  wire [0:0] arrdiv32_fs308_xor1;
  wire [0:0] arrdiv32_fs308_or0;
  wire [0:0] arrdiv32_fs309_xor1;
  wire [0:0] arrdiv32_fs309_or0;
  wire [0:0] arrdiv32_fs310_xor1;
  wire [0:0] arrdiv32_fs310_or0;
  wire [0:0] arrdiv32_fs311_xor1;
  wire [0:0] arrdiv32_fs311_or0;
  wire [0:0] arrdiv32_fs312_xor1;
  wire [0:0] arrdiv32_fs312_or0;
  wire [0:0] arrdiv32_fs313_xor1;
  wire [0:0] arrdiv32_fs313_or0;
  wire [0:0] arrdiv32_fs314_xor1;
  wire [0:0] arrdiv32_fs314_or0;
  wire [0:0] arrdiv32_fs315_xor1;
  wire [0:0] arrdiv32_fs315_or0;
  wire [0:0] arrdiv32_fs316_xor1;
  wire [0:0] arrdiv32_fs316_or0;
  wire [0:0] arrdiv32_fs317_xor1;
  wire [0:0] arrdiv32_fs317_or0;
  wire [0:0] arrdiv32_fs318_xor1;
  wire [0:0] arrdiv32_fs318_or0;
  wire [0:0] arrdiv32_fs319_xor1;
  wire [0:0] arrdiv32_fs319_or0;
  wire [0:0] arrdiv32_mux2to1279_xor0;
  wire [0:0] arrdiv32_mux2to1280_xor0;
  wire [0:0] arrdiv32_mux2to1281_xor0;
  wire [0:0] arrdiv32_mux2to1282_xor0;
  wire [0:0] arrdiv32_mux2to1283_xor0;
  wire [0:0] arrdiv32_mux2to1284_xor0;
  wire [0:0] arrdiv32_mux2to1285_xor0;
  wire [0:0] arrdiv32_mux2to1286_xor0;
  wire [0:0] arrdiv32_mux2to1287_xor0;
  wire [0:0] arrdiv32_mux2to1288_xor0;
  wire [0:0] arrdiv32_mux2to1289_xor0;
  wire [0:0] arrdiv32_mux2to1290_xor0;
  wire [0:0] arrdiv32_mux2to1291_xor0;
  wire [0:0] arrdiv32_mux2to1292_xor0;
  wire [0:0] arrdiv32_mux2to1293_xor0;
  wire [0:0] arrdiv32_mux2to1294_xor0;
  wire [0:0] arrdiv32_mux2to1295_xor0;
  wire [0:0] arrdiv32_mux2to1296_xor0;
  wire [0:0] arrdiv32_mux2to1297_xor0;
  wire [0:0] arrdiv32_mux2to1298_xor0;
  wire [0:0] arrdiv32_mux2to1299_xor0;
  wire [0:0] arrdiv32_mux2to1300_xor0;
  wire [0:0] arrdiv32_mux2to1301_xor0;
  wire [0:0] arrdiv32_mux2to1302_xor0;
  wire [0:0] arrdiv32_mux2to1303_xor0;
  wire [0:0] arrdiv32_mux2to1304_xor0;
  wire [0:0] arrdiv32_mux2to1305_xor0;
  wire [0:0] arrdiv32_mux2to1306_xor0;
  wire [0:0] arrdiv32_mux2to1307_xor0;
  wire [0:0] arrdiv32_mux2to1308_xor0;
  wire [0:0] arrdiv32_mux2to1309_xor0;
  wire [0:0] arrdiv32_not9;
  wire [0:0] arrdiv32_fs320_xor0;
  wire [0:0] arrdiv32_fs320_and0;
  wire [0:0] arrdiv32_fs321_xor1;
  wire [0:0] arrdiv32_fs321_or0;
  wire [0:0] arrdiv32_fs322_xor1;
  wire [0:0] arrdiv32_fs322_or0;
  wire [0:0] arrdiv32_fs323_xor1;
  wire [0:0] arrdiv32_fs323_or0;
  wire [0:0] arrdiv32_fs324_xor1;
  wire [0:0] arrdiv32_fs324_or0;
  wire [0:0] arrdiv32_fs325_xor1;
  wire [0:0] arrdiv32_fs325_or0;
  wire [0:0] arrdiv32_fs326_xor1;
  wire [0:0] arrdiv32_fs326_or0;
  wire [0:0] arrdiv32_fs327_xor1;
  wire [0:0] arrdiv32_fs327_or0;
  wire [0:0] arrdiv32_fs328_xor1;
  wire [0:0] arrdiv32_fs328_or0;
  wire [0:0] arrdiv32_fs329_xor1;
  wire [0:0] arrdiv32_fs329_or0;
  wire [0:0] arrdiv32_fs330_xor1;
  wire [0:0] arrdiv32_fs330_or0;
  wire [0:0] arrdiv32_fs331_xor1;
  wire [0:0] arrdiv32_fs331_or0;
  wire [0:0] arrdiv32_fs332_xor1;
  wire [0:0] arrdiv32_fs332_or0;
  wire [0:0] arrdiv32_fs333_xor1;
  wire [0:0] arrdiv32_fs333_or0;
  wire [0:0] arrdiv32_fs334_xor1;
  wire [0:0] arrdiv32_fs334_or0;
  wire [0:0] arrdiv32_fs335_xor1;
  wire [0:0] arrdiv32_fs335_or0;
  wire [0:0] arrdiv32_fs336_xor1;
  wire [0:0] arrdiv32_fs336_or0;
  wire [0:0] arrdiv32_fs337_xor1;
  wire [0:0] arrdiv32_fs337_or0;
  wire [0:0] arrdiv32_fs338_xor1;
  wire [0:0] arrdiv32_fs338_or0;
  wire [0:0] arrdiv32_fs339_xor1;
  wire [0:0] arrdiv32_fs339_or0;
  wire [0:0] arrdiv32_fs340_xor1;
  wire [0:0] arrdiv32_fs340_or0;
  wire [0:0] arrdiv32_fs341_xor1;
  wire [0:0] arrdiv32_fs341_or0;
  wire [0:0] arrdiv32_fs342_xor1;
  wire [0:0] arrdiv32_fs342_or0;
  wire [0:0] arrdiv32_fs343_xor1;
  wire [0:0] arrdiv32_fs343_or0;
  wire [0:0] arrdiv32_fs344_xor1;
  wire [0:0] arrdiv32_fs344_or0;
  wire [0:0] arrdiv32_fs345_xor1;
  wire [0:0] arrdiv32_fs345_or0;
  wire [0:0] arrdiv32_fs346_xor1;
  wire [0:0] arrdiv32_fs346_or0;
  wire [0:0] arrdiv32_fs347_xor1;
  wire [0:0] arrdiv32_fs347_or0;
  wire [0:0] arrdiv32_fs348_xor1;
  wire [0:0] arrdiv32_fs348_or0;
  wire [0:0] arrdiv32_fs349_xor1;
  wire [0:0] arrdiv32_fs349_or0;
  wire [0:0] arrdiv32_fs350_xor1;
  wire [0:0] arrdiv32_fs350_or0;
  wire [0:0] arrdiv32_fs351_xor1;
  wire [0:0] arrdiv32_fs351_or0;
  wire [0:0] arrdiv32_mux2to1310_xor0;
  wire [0:0] arrdiv32_mux2to1311_xor0;
  wire [0:0] arrdiv32_mux2to1312_xor0;
  wire [0:0] arrdiv32_mux2to1313_xor0;
  wire [0:0] arrdiv32_mux2to1314_xor0;
  wire [0:0] arrdiv32_mux2to1315_xor0;
  wire [0:0] arrdiv32_mux2to1316_xor0;
  wire [0:0] arrdiv32_mux2to1317_xor0;
  wire [0:0] arrdiv32_mux2to1318_xor0;
  wire [0:0] arrdiv32_mux2to1319_xor0;
  wire [0:0] arrdiv32_mux2to1320_xor0;
  wire [0:0] arrdiv32_mux2to1321_xor0;
  wire [0:0] arrdiv32_mux2to1322_xor0;
  wire [0:0] arrdiv32_mux2to1323_xor0;
  wire [0:0] arrdiv32_mux2to1324_xor0;
  wire [0:0] arrdiv32_mux2to1325_xor0;
  wire [0:0] arrdiv32_mux2to1326_xor0;
  wire [0:0] arrdiv32_mux2to1327_xor0;
  wire [0:0] arrdiv32_mux2to1328_xor0;
  wire [0:0] arrdiv32_mux2to1329_xor0;
  wire [0:0] arrdiv32_mux2to1330_xor0;
  wire [0:0] arrdiv32_mux2to1331_xor0;
  wire [0:0] arrdiv32_mux2to1332_xor0;
  wire [0:0] arrdiv32_mux2to1333_xor0;
  wire [0:0] arrdiv32_mux2to1334_xor0;
  wire [0:0] arrdiv32_mux2to1335_xor0;
  wire [0:0] arrdiv32_mux2to1336_xor0;
  wire [0:0] arrdiv32_mux2to1337_xor0;
  wire [0:0] arrdiv32_mux2to1338_xor0;
  wire [0:0] arrdiv32_mux2to1339_xor0;
  wire [0:0] arrdiv32_mux2to1340_xor0;
  wire [0:0] arrdiv32_not10;
  wire [0:0] arrdiv32_fs352_xor0;
  wire [0:0] arrdiv32_fs352_and0;
  wire [0:0] arrdiv32_fs353_xor1;
  wire [0:0] arrdiv32_fs353_or0;
  wire [0:0] arrdiv32_fs354_xor1;
  wire [0:0] arrdiv32_fs354_or0;
  wire [0:0] arrdiv32_fs355_xor1;
  wire [0:0] arrdiv32_fs355_or0;
  wire [0:0] arrdiv32_fs356_xor1;
  wire [0:0] arrdiv32_fs356_or0;
  wire [0:0] arrdiv32_fs357_xor1;
  wire [0:0] arrdiv32_fs357_or0;
  wire [0:0] arrdiv32_fs358_xor1;
  wire [0:0] arrdiv32_fs358_or0;
  wire [0:0] arrdiv32_fs359_xor1;
  wire [0:0] arrdiv32_fs359_or0;
  wire [0:0] arrdiv32_fs360_xor1;
  wire [0:0] arrdiv32_fs360_or0;
  wire [0:0] arrdiv32_fs361_xor1;
  wire [0:0] arrdiv32_fs361_or0;
  wire [0:0] arrdiv32_fs362_xor1;
  wire [0:0] arrdiv32_fs362_or0;
  wire [0:0] arrdiv32_fs363_xor1;
  wire [0:0] arrdiv32_fs363_or0;
  wire [0:0] arrdiv32_fs364_xor1;
  wire [0:0] arrdiv32_fs364_or0;
  wire [0:0] arrdiv32_fs365_xor1;
  wire [0:0] arrdiv32_fs365_or0;
  wire [0:0] arrdiv32_fs366_xor1;
  wire [0:0] arrdiv32_fs366_or0;
  wire [0:0] arrdiv32_fs367_xor1;
  wire [0:0] arrdiv32_fs367_or0;
  wire [0:0] arrdiv32_fs368_xor1;
  wire [0:0] arrdiv32_fs368_or0;
  wire [0:0] arrdiv32_fs369_xor1;
  wire [0:0] arrdiv32_fs369_or0;
  wire [0:0] arrdiv32_fs370_xor1;
  wire [0:0] arrdiv32_fs370_or0;
  wire [0:0] arrdiv32_fs371_xor1;
  wire [0:0] arrdiv32_fs371_or0;
  wire [0:0] arrdiv32_fs372_xor1;
  wire [0:0] arrdiv32_fs372_or0;
  wire [0:0] arrdiv32_fs373_xor1;
  wire [0:0] arrdiv32_fs373_or0;
  wire [0:0] arrdiv32_fs374_xor1;
  wire [0:0] arrdiv32_fs374_or0;
  wire [0:0] arrdiv32_fs375_xor1;
  wire [0:0] arrdiv32_fs375_or0;
  wire [0:0] arrdiv32_fs376_xor1;
  wire [0:0] arrdiv32_fs376_or0;
  wire [0:0] arrdiv32_fs377_xor1;
  wire [0:0] arrdiv32_fs377_or0;
  wire [0:0] arrdiv32_fs378_xor1;
  wire [0:0] arrdiv32_fs378_or0;
  wire [0:0] arrdiv32_fs379_xor1;
  wire [0:0] arrdiv32_fs379_or0;
  wire [0:0] arrdiv32_fs380_xor1;
  wire [0:0] arrdiv32_fs380_or0;
  wire [0:0] arrdiv32_fs381_xor1;
  wire [0:0] arrdiv32_fs381_or0;
  wire [0:0] arrdiv32_fs382_xor1;
  wire [0:0] arrdiv32_fs382_or0;
  wire [0:0] arrdiv32_fs383_xor1;
  wire [0:0] arrdiv32_fs383_or0;
  wire [0:0] arrdiv32_mux2to1341_xor0;
  wire [0:0] arrdiv32_mux2to1342_xor0;
  wire [0:0] arrdiv32_mux2to1343_xor0;
  wire [0:0] arrdiv32_mux2to1344_xor0;
  wire [0:0] arrdiv32_mux2to1345_xor0;
  wire [0:0] arrdiv32_mux2to1346_xor0;
  wire [0:0] arrdiv32_mux2to1347_xor0;
  wire [0:0] arrdiv32_mux2to1348_xor0;
  wire [0:0] arrdiv32_mux2to1349_xor0;
  wire [0:0] arrdiv32_mux2to1350_xor0;
  wire [0:0] arrdiv32_mux2to1351_xor0;
  wire [0:0] arrdiv32_mux2to1352_xor0;
  wire [0:0] arrdiv32_mux2to1353_xor0;
  wire [0:0] arrdiv32_mux2to1354_xor0;
  wire [0:0] arrdiv32_mux2to1355_xor0;
  wire [0:0] arrdiv32_mux2to1356_xor0;
  wire [0:0] arrdiv32_mux2to1357_xor0;
  wire [0:0] arrdiv32_mux2to1358_xor0;
  wire [0:0] arrdiv32_mux2to1359_xor0;
  wire [0:0] arrdiv32_mux2to1360_xor0;
  wire [0:0] arrdiv32_mux2to1361_xor0;
  wire [0:0] arrdiv32_mux2to1362_xor0;
  wire [0:0] arrdiv32_mux2to1363_xor0;
  wire [0:0] arrdiv32_mux2to1364_xor0;
  wire [0:0] arrdiv32_mux2to1365_xor0;
  wire [0:0] arrdiv32_mux2to1366_xor0;
  wire [0:0] arrdiv32_mux2to1367_xor0;
  wire [0:0] arrdiv32_mux2to1368_xor0;
  wire [0:0] arrdiv32_mux2to1369_xor0;
  wire [0:0] arrdiv32_mux2to1370_xor0;
  wire [0:0] arrdiv32_mux2to1371_xor0;
  wire [0:0] arrdiv32_not11;
  wire [0:0] arrdiv32_fs384_xor0;
  wire [0:0] arrdiv32_fs384_and0;
  wire [0:0] arrdiv32_fs385_xor1;
  wire [0:0] arrdiv32_fs385_or0;
  wire [0:0] arrdiv32_fs386_xor1;
  wire [0:0] arrdiv32_fs386_or0;
  wire [0:0] arrdiv32_fs387_xor1;
  wire [0:0] arrdiv32_fs387_or0;
  wire [0:0] arrdiv32_fs388_xor1;
  wire [0:0] arrdiv32_fs388_or0;
  wire [0:0] arrdiv32_fs389_xor1;
  wire [0:0] arrdiv32_fs389_or0;
  wire [0:0] arrdiv32_fs390_xor1;
  wire [0:0] arrdiv32_fs390_or0;
  wire [0:0] arrdiv32_fs391_xor1;
  wire [0:0] arrdiv32_fs391_or0;
  wire [0:0] arrdiv32_fs392_xor1;
  wire [0:0] arrdiv32_fs392_or0;
  wire [0:0] arrdiv32_fs393_xor1;
  wire [0:0] arrdiv32_fs393_or0;
  wire [0:0] arrdiv32_fs394_xor1;
  wire [0:0] arrdiv32_fs394_or0;
  wire [0:0] arrdiv32_fs395_xor1;
  wire [0:0] arrdiv32_fs395_or0;
  wire [0:0] arrdiv32_fs396_xor1;
  wire [0:0] arrdiv32_fs396_or0;
  wire [0:0] arrdiv32_fs397_xor1;
  wire [0:0] arrdiv32_fs397_or0;
  wire [0:0] arrdiv32_fs398_xor1;
  wire [0:0] arrdiv32_fs398_or0;
  wire [0:0] arrdiv32_fs399_xor1;
  wire [0:0] arrdiv32_fs399_or0;
  wire [0:0] arrdiv32_fs400_xor1;
  wire [0:0] arrdiv32_fs400_or0;
  wire [0:0] arrdiv32_fs401_xor1;
  wire [0:0] arrdiv32_fs401_or0;
  wire [0:0] arrdiv32_fs402_xor1;
  wire [0:0] arrdiv32_fs402_or0;
  wire [0:0] arrdiv32_fs403_xor1;
  wire [0:0] arrdiv32_fs403_or0;
  wire [0:0] arrdiv32_fs404_xor1;
  wire [0:0] arrdiv32_fs404_or0;
  wire [0:0] arrdiv32_fs405_xor1;
  wire [0:0] arrdiv32_fs405_or0;
  wire [0:0] arrdiv32_fs406_xor1;
  wire [0:0] arrdiv32_fs406_or0;
  wire [0:0] arrdiv32_fs407_xor1;
  wire [0:0] arrdiv32_fs407_or0;
  wire [0:0] arrdiv32_fs408_xor1;
  wire [0:0] arrdiv32_fs408_or0;
  wire [0:0] arrdiv32_fs409_xor1;
  wire [0:0] arrdiv32_fs409_or0;
  wire [0:0] arrdiv32_fs410_xor1;
  wire [0:0] arrdiv32_fs410_or0;
  wire [0:0] arrdiv32_fs411_xor1;
  wire [0:0] arrdiv32_fs411_or0;
  wire [0:0] arrdiv32_fs412_xor1;
  wire [0:0] arrdiv32_fs412_or0;
  wire [0:0] arrdiv32_fs413_xor1;
  wire [0:0] arrdiv32_fs413_or0;
  wire [0:0] arrdiv32_fs414_xor1;
  wire [0:0] arrdiv32_fs414_or0;
  wire [0:0] arrdiv32_fs415_xor1;
  wire [0:0] arrdiv32_fs415_or0;
  wire [0:0] arrdiv32_mux2to1372_xor0;
  wire [0:0] arrdiv32_mux2to1373_xor0;
  wire [0:0] arrdiv32_mux2to1374_xor0;
  wire [0:0] arrdiv32_mux2to1375_xor0;
  wire [0:0] arrdiv32_mux2to1376_xor0;
  wire [0:0] arrdiv32_mux2to1377_xor0;
  wire [0:0] arrdiv32_mux2to1378_xor0;
  wire [0:0] arrdiv32_mux2to1379_xor0;
  wire [0:0] arrdiv32_mux2to1380_xor0;
  wire [0:0] arrdiv32_mux2to1381_xor0;
  wire [0:0] arrdiv32_mux2to1382_xor0;
  wire [0:0] arrdiv32_mux2to1383_xor0;
  wire [0:0] arrdiv32_mux2to1384_xor0;
  wire [0:0] arrdiv32_mux2to1385_xor0;
  wire [0:0] arrdiv32_mux2to1386_xor0;
  wire [0:0] arrdiv32_mux2to1387_xor0;
  wire [0:0] arrdiv32_mux2to1388_xor0;
  wire [0:0] arrdiv32_mux2to1389_xor0;
  wire [0:0] arrdiv32_mux2to1390_xor0;
  wire [0:0] arrdiv32_mux2to1391_xor0;
  wire [0:0] arrdiv32_mux2to1392_xor0;
  wire [0:0] arrdiv32_mux2to1393_xor0;
  wire [0:0] arrdiv32_mux2to1394_xor0;
  wire [0:0] arrdiv32_mux2to1395_xor0;
  wire [0:0] arrdiv32_mux2to1396_xor0;
  wire [0:0] arrdiv32_mux2to1397_xor0;
  wire [0:0] arrdiv32_mux2to1398_xor0;
  wire [0:0] arrdiv32_mux2to1399_xor0;
  wire [0:0] arrdiv32_mux2to1400_xor0;
  wire [0:0] arrdiv32_mux2to1401_xor0;
  wire [0:0] arrdiv32_mux2to1402_xor0;
  wire [0:0] arrdiv32_not12;
  wire [0:0] arrdiv32_fs416_xor0;
  wire [0:0] arrdiv32_fs416_and0;
  wire [0:0] arrdiv32_fs417_xor1;
  wire [0:0] arrdiv32_fs417_or0;
  wire [0:0] arrdiv32_fs418_xor1;
  wire [0:0] arrdiv32_fs418_or0;
  wire [0:0] arrdiv32_fs419_xor1;
  wire [0:0] arrdiv32_fs419_or0;
  wire [0:0] arrdiv32_fs420_xor1;
  wire [0:0] arrdiv32_fs420_or0;
  wire [0:0] arrdiv32_fs421_xor1;
  wire [0:0] arrdiv32_fs421_or0;
  wire [0:0] arrdiv32_fs422_xor1;
  wire [0:0] arrdiv32_fs422_or0;
  wire [0:0] arrdiv32_fs423_xor1;
  wire [0:0] arrdiv32_fs423_or0;
  wire [0:0] arrdiv32_fs424_xor1;
  wire [0:0] arrdiv32_fs424_or0;
  wire [0:0] arrdiv32_fs425_xor1;
  wire [0:0] arrdiv32_fs425_or0;
  wire [0:0] arrdiv32_fs426_xor1;
  wire [0:0] arrdiv32_fs426_or0;
  wire [0:0] arrdiv32_fs427_xor1;
  wire [0:0] arrdiv32_fs427_or0;
  wire [0:0] arrdiv32_fs428_xor1;
  wire [0:0] arrdiv32_fs428_or0;
  wire [0:0] arrdiv32_fs429_xor1;
  wire [0:0] arrdiv32_fs429_or0;
  wire [0:0] arrdiv32_fs430_xor1;
  wire [0:0] arrdiv32_fs430_or0;
  wire [0:0] arrdiv32_fs431_xor1;
  wire [0:0] arrdiv32_fs431_or0;
  wire [0:0] arrdiv32_fs432_xor1;
  wire [0:0] arrdiv32_fs432_or0;
  wire [0:0] arrdiv32_fs433_xor1;
  wire [0:0] arrdiv32_fs433_or0;
  wire [0:0] arrdiv32_fs434_xor1;
  wire [0:0] arrdiv32_fs434_or0;
  wire [0:0] arrdiv32_fs435_xor1;
  wire [0:0] arrdiv32_fs435_or0;
  wire [0:0] arrdiv32_fs436_xor1;
  wire [0:0] arrdiv32_fs436_or0;
  wire [0:0] arrdiv32_fs437_xor1;
  wire [0:0] arrdiv32_fs437_or0;
  wire [0:0] arrdiv32_fs438_xor1;
  wire [0:0] arrdiv32_fs438_or0;
  wire [0:0] arrdiv32_fs439_xor1;
  wire [0:0] arrdiv32_fs439_or0;
  wire [0:0] arrdiv32_fs440_xor1;
  wire [0:0] arrdiv32_fs440_or0;
  wire [0:0] arrdiv32_fs441_xor1;
  wire [0:0] arrdiv32_fs441_or0;
  wire [0:0] arrdiv32_fs442_xor1;
  wire [0:0] arrdiv32_fs442_or0;
  wire [0:0] arrdiv32_fs443_xor1;
  wire [0:0] arrdiv32_fs443_or0;
  wire [0:0] arrdiv32_fs444_xor1;
  wire [0:0] arrdiv32_fs444_or0;
  wire [0:0] arrdiv32_fs445_xor1;
  wire [0:0] arrdiv32_fs445_or0;
  wire [0:0] arrdiv32_fs446_xor1;
  wire [0:0] arrdiv32_fs446_or0;
  wire [0:0] arrdiv32_fs447_xor1;
  wire [0:0] arrdiv32_fs447_or0;
  wire [0:0] arrdiv32_mux2to1403_xor0;
  wire [0:0] arrdiv32_mux2to1404_xor0;
  wire [0:0] arrdiv32_mux2to1405_xor0;
  wire [0:0] arrdiv32_mux2to1406_xor0;
  wire [0:0] arrdiv32_mux2to1407_xor0;
  wire [0:0] arrdiv32_mux2to1408_xor0;
  wire [0:0] arrdiv32_mux2to1409_xor0;
  wire [0:0] arrdiv32_mux2to1410_xor0;
  wire [0:0] arrdiv32_mux2to1411_xor0;
  wire [0:0] arrdiv32_mux2to1412_xor0;
  wire [0:0] arrdiv32_mux2to1413_xor0;
  wire [0:0] arrdiv32_mux2to1414_xor0;
  wire [0:0] arrdiv32_mux2to1415_xor0;
  wire [0:0] arrdiv32_mux2to1416_xor0;
  wire [0:0] arrdiv32_mux2to1417_xor0;
  wire [0:0] arrdiv32_mux2to1418_xor0;
  wire [0:0] arrdiv32_mux2to1419_xor0;
  wire [0:0] arrdiv32_mux2to1420_xor0;
  wire [0:0] arrdiv32_mux2to1421_xor0;
  wire [0:0] arrdiv32_mux2to1422_xor0;
  wire [0:0] arrdiv32_mux2to1423_xor0;
  wire [0:0] arrdiv32_mux2to1424_xor0;
  wire [0:0] arrdiv32_mux2to1425_xor0;
  wire [0:0] arrdiv32_mux2to1426_xor0;
  wire [0:0] arrdiv32_mux2to1427_xor0;
  wire [0:0] arrdiv32_mux2to1428_xor0;
  wire [0:0] arrdiv32_mux2to1429_xor0;
  wire [0:0] arrdiv32_mux2to1430_xor0;
  wire [0:0] arrdiv32_mux2to1431_xor0;
  wire [0:0] arrdiv32_mux2to1432_xor0;
  wire [0:0] arrdiv32_mux2to1433_xor0;
  wire [0:0] arrdiv32_not13;
  wire [0:0] arrdiv32_fs448_xor0;
  wire [0:0] arrdiv32_fs448_and0;
  wire [0:0] arrdiv32_fs449_xor1;
  wire [0:0] arrdiv32_fs449_or0;
  wire [0:0] arrdiv32_fs450_xor1;
  wire [0:0] arrdiv32_fs450_or0;
  wire [0:0] arrdiv32_fs451_xor1;
  wire [0:0] arrdiv32_fs451_or0;
  wire [0:0] arrdiv32_fs452_xor1;
  wire [0:0] arrdiv32_fs452_or0;
  wire [0:0] arrdiv32_fs453_xor1;
  wire [0:0] arrdiv32_fs453_or0;
  wire [0:0] arrdiv32_fs454_xor1;
  wire [0:0] arrdiv32_fs454_or0;
  wire [0:0] arrdiv32_fs455_xor1;
  wire [0:0] arrdiv32_fs455_or0;
  wire [0:0] arrdiv32_fs456_xor1;
  wire [0:0] arrdiv32_fs456_or0;
  wire [0:0] arrdiv32_fs457_xor1;
  wire [0:0] arrdiv32_fs457_or0;
  wire [0:0] arrdiv32_fs458_xor1;
  wire [0:0] arrdiv32_fs458_or0;
  wire [0:0] arrdiv32_fs459_xor1;
  wire [0:0] arrdiv32_fs459_or0;
  wire [0:0] arrdiv32_fs460_xor1;
  wire [0:0] arrdiv32_fs460_or0;
  wire [0:0] arrdiv32_fs461_xor1;
  wire [0:0] arrdiv32_fs461_or0;
  wire [0:0] arrdiv32_fs462_xor1;
  wire [0:0] arrdiv32_fs462_or0;
  wire [0:0] arrdiv32_fs463_xor1;
  wire [0:0] arrdiv32_fs463_or0;
  wire [0:0] arrdiv32_fs464_xor1;
  wire [0:0] arrdiv32_fs464_or0;
  wire [0:0] arrdiv32_fs465_xor1;
  wire [0:0] arrdiv32_fs465_or0;
  wire [0:0] arrdiv32_fs466_xor1;
  wire [0:0] arrdiv32_fs466_or0;
  wire [0:0] arrdiv32_fs467_xor1;
  wire [0:0] arrdiv32_fs467_or0;
  wire [0:0] arrdiv32_fs468_xor1;
  wire [0:0] arrdiv32_fs468_or0;
  wire [0:0] arrdiv32_fs469_xor1;
  wire [0:0] arrdiv32_fs469_or0;
  wire [0:0] arrdiv32_fs470_xor1;
  wire [0:0] arrdiv32_fs470_or0;
  wire [0:0] arrdiv32_fs471_xor1;
  wire [0:0] arrdiv32_fs471_or0;
  wire [0:0] arrdiv32_fs472_xor1;
  wire [0:0] arrdiv32_fs472_or0;
  wire [0:0] arrdiv32_fs473_xor1;
  wire [0:0] arrdiv32_fs473_or0;
  wire [0:0] arrdiv32_fs474_xor1;
  wire [0:0] arrdiv32_fs474_or0;
  wire [0:0] arrdiv32_fs475_xor1;
  wire [0:0] arrdiv32_fs475_or0;
  wire [0:0] arrdiv32_fs476_xor1;
  wire [0:0] arrdiv32_fs476_or0;
  wire [0:0] arrdiv32_fs477_xor1;
  wire [0:0] arrdiv32_fs477_or0;
  wire [0:0] arrdiv32_fs478_xor1;
  wire [0:0] arrdiv32_fs478_or0;
  wire [0:0] arrdiv32_fs479_xor1;
  wire [0:0] arrdiv32_fs479_or0;
  wire [0:0] arrdiv32_mux2to1434_xor0;
  wire [0:0] arrdiv32_mux2to1435_xor0;
  wire [0:0] arrdiv32_mux2to1436_xor0;
  wire [0:0] arrdiv32_mux2to1437_xor0;
  wire [0:0] arrdiv32_mux2to1438_xor0;
  wire [0:0] arrdiv32_mux2to1439_xor0;
  wire [0:0] arrdiv32_mux2to1440_xor0;
  wire [0:0] arrdiv32_mux2to1441_xor0;
  wire [0:0] arrdiv32_mux2to1442_xor0;
  wire [0:0] arrdiv32_mux2to1443_xor0;
  wire [0:0] arrdiv32_mux2to1444_xor0;
  wire [0:0] arrdiv32_mux2to1445_xor0;
  wire [0:0] arrdiv32_mux2to1446_xor0;
  wire [0:0] arrdiv32_mux2to1447_xor0;
  wire [0:0] arrdiv32_mux2to1448_xor0;
  wire [0:0] arrdiv32_mux2to1449_xor0;
  wire [0:0] arrdiv32_mux2to1450_xor0;
  wire [0:0] arrdiv32_mux2to1451_xor0;
  wire [0:0] arrdiv32_mux2to1452_xor0;
  wire [0:0] arrdiv32_mux2to1453_xor0;
  wire [0:0] arrdiv32_mux2to1454_xor0;
  wire [0:0] arrdiv32_mux2to1455_xor0;
  wire [0:0] arrdiv32_mux2to1456_xor0;
  wire [0:0] arrdiv32_mux2to1457_xor0;
  wire [0:0] arrdiv32_mux2to1458_xor0;
  wire [0:0] arrdiv32_mux2to1459_xor0;
  wire [0:0] arrdiv32_mux2to1460_xor0;
  wire [0:0] arrdiv32_mux2to1461_xor0;
  wire [0:0] arrdiv32_mux2to1462_xor0;
  wire [0:0] arrdiv32_mux2to1463_xor0;
  wire [0:0] arrdiv32_mux2to1464_xor0;
  wire [0:0] arrdiv32_not14;
  wire [0:0] arrdiv32_fs480_xor0;
  wire [0:0] arrdiv32_fs480_and0;
  wire [0:0] arrdiv32_fs481_xor1;
  wire [0:0] arrdiv32_fs481_or0;
  wire [0:0] arrdiv32_fs482_xor1;
  wire [0:0] arrdiv32_fs482_or0;
  wire [0:0] arrdiv32_fs483_xor1;
  wire [0:0] arrdiv32_fs483_or0;
  wire [0:0] arrdiv32_fs484_xor1;
  wire [0:0] arrdiv32_fs484_or0;
  wire [0:0] arrdiv32_fs485_xor1;
  wire [0:0] arrdiv32_fs485_or0;
  wire [0:0] arrdiv32_fs486_xor1;
  wire [0:0] arrdiv32_fs486_or0;
  wire [0:0] arrdiv32_fs487_xor1;
  wire [0:0] arrdiv32_fs487_or0;
  wire [0:0] arrdiv32_fs488_xor1;
  wire [0:0] arrdiv32_fs488_or0;
  wire [0:0] arrdiv32_fs489_xor1;
  wire [0:0] arrdiv32_fs489_or0;
  wire [0:0] arrdiv32_fs490_xor1;
  wire [0:0] arrdiv32_fs490_or0;
  wire [0:0] arrdiv32_fs491_xor1;
  wire [0:0] arrdiv32_fs491_or0;
  wire [0:0] arrdiv32_fs492_xor1;
  wire [0:0] arrdiv32_fs492_or0;
  wire [0:0] arrdiv32_fs493_xor1;
  wire [0:0] arrdiv32_fs493_or0;
  wire [0:0] arrdiv32_fs494_xor1;
  wire [0:0] arrdiv32_fs494_or0;
  wire [0:0] arrdiv32_fs495_xor1;
  wire [0:0] arrdiv32_fs495_or0;
  wire [0:0] arrdiv32_fs496_xor1;
  wire [0:0] arrdiv32_fs496_or0;
  wire [0:0] arrdiv32_fs497_xor1;
  wire [0:0] arrdiv32_fs497_or0;
  wire [0:0] arrdiv32_fs498_xor1;
  wire [0:0] arrdiv32_fs498_or0;
  wire [0:0] arrdiv32_fs499_xor1;
  wire [0:0] arrdiv32_fs499_or0;
  wire [0:0] arrdiv32_fs500_xor1;
  wire [0:0] arrdiv32_fs500_or0;
  wire [0:0] arrdiv32_fs501_xor1;
  wire [0:0] arrdiv32_fs501_or0;
  wire [0:0] arrdiv32_fs502_xor1;
  wire [0:0] arrdiv32_fs502_or0;
  wire [0:0] arrdiv32_fs503_xor1;
  wire [0:0] arrdiv32_fs503_or0;
  wire [0:0] arrdiv32_fs504_xor1;
  wire [0:0] arrdiv32_fs504_or0;
  wire [0:0] arrdiv32_fs505_xor1;
  wire [0:0] arrdiv32_fs505_or0;
  wire [0:0] arrdiv32_fs506_xor1;
  wire [0:0] arrdiv32_fs506_or0;
  wire [0:0] arrdiv32_fs507_xor1;
  wire [0:0] arrdiv32_fs507_or0;
  wire [0:0] arrdiv32_fs508_xor1;
  wire [0:0] arrdiv32_fs508_or0;
  wire [0:0] arrdiv32_fs509_xor1;
  wire [0:0] arrdiv32_fs509_or0;
  wire [0:0] arrdiv32_fs510_xor1;
  wire [0:0] arrdiv32_fs510_or0;
  wire [0:0] arrdiv32_fs511_xor1;
  wire [0:0] arrdiv32_fs511_or0;
  wire [0:0] arrdiv32_mux2to1465_xor0;
  wire [0:0] arrdiv32_mux2to1466_xor0;
  wire [0:0] arrdiv32_mux2to1467_xor0;
  wire [0:0] arrdiv32_mux2to1468_xor0;
  wire [0:0] arrdiv32_mux2to1469_xor0;
  wire [0:0] arrdiv32_mux2to1470_xor0;
  wire [0:0] arrdiv32_mux2to1471_xor0;
  wire [0:0] arrdiv32_mux2to1472_xor0;
  wire [0:0] arrdiv32_mux2to1473_xor0;
  wire [0:0] arrdiv32_mux2to1474_xor0;
  wire [0:0] arrdiv32_mux2to1475_xor0;
  wire [0:0] arrdiv32_mux2to1476_xor0;
  wire [0:0] arrdiv32_mux2to1477_xor0;
  wire [0:0] arrdiv32_mux2to1478_xor0;
  wire [0:0] arrdiv32_mux2to1479_xor0;
  wire [0:0] arrdiv32_mux2to1480_xor0;
  wire [0:0] arrdiv32_mux2to1481_xor0;
  wire [0:0] arrdiv32_mux2to1482_xor0;
  wire [0:0] arrdiv32_mux2to1483_xor0;
  wire [0:0] arrdiv32_mux2to1484_xor0;
  wire [0:0] arrdiv32_mux2to1485_xor0;
  wire [0:0] arrdiv32_mux2to1486_xor0;
  wire [0:0] arrdiv32_mux2to1487_xor0;
  wire [0:0] arrdiv32_mux2to1488_xor0;
  wire [0:0] arrdiv32_mux2to1489_xor0;
  wire [0:0] arrdiv32_mux2to1490_xor0;
  wire [0:0] arrdiv32_mux2to1491_xor0;
  wire [0:0] arrdiv32_mux2to1492_xor0;
  wire [0:0] arrdiv32_mux2to1493_xor0;
  wire [0:0] arrdiv32_mux2to1494_xor0;
  wire [0:0] arrdiv32_mux2to1495_xor0;
  wire [0:0] arrdiv32_not15;
  wire [0:0] arrdiv32_fs512_xor0;
  wire [0:0] arrdiv32_fs512_and0;
  wire [0:0] arrdiv32_fs513_xor1;
  wire [0:0] arrdiv32_fs513_or0;
  wire [0:0] arrdiv32_fs514_xor1;
  wire [0:0] arrdiv32_fs514_or0;
  wire [0:0] arrdiv32_fs515_xor1;
  wire [0:0] arrdiv32_fs515_or0;
  wire [0:0] arrdiv32_fs516_xor1;
  wire [0:0] arrdiv32_fs516_or0;
  wire [0:0] arrdiv32_fs517_xor1;
  wire [0:0] arrdiv32_fs517_or0;
  wire [0:0] arrdiv32_fs518_xor1;
  wire [0:0] arrdiv32_fs518_or0;
  wire [0:0] arrdiv32_fs519_xor1;
  wire [0:0] arrdiv32_fs519_or0;
  wire [0:0] arrdiv32_fs520_xor1;
  wire [0:0] arrdiv32_fs520_or0;
  wire [0:0] arrdiv32_fs521_xor1;
  wire [0:0] arrdiv32_fs521_or0;
  wire [0:0] arrdiv32_fs522_xor1;
  wire [0:0] arrdiv32_fs522_or0;
  wire [0:0] arrdiv32_fs523_xor1;
  wire [0:0] arrdiv32_fs523_or0;
  wire [0:0] arrdiv32_fs524_xor1;
  wire [0:0] arrdiv32_fs524_or0;
  wire [0:0] arrdiv32_fs525_xor1;
  wire [0:0] arrdiv32_fs525_or0;
  wire [0:0] arrdiv32_fs526_xor1;
  wire [0:0] arrdiv32_fs526_or0;
  wire [0:0] arrdiv32_fs527_xor1;
  wire [0:0] arrdiv32_fs527_or0;
  wire [0:0] arrdiv32_fs528_xor1;
  wire [0:0] arrdiv32_fs528_or0;
  wire [0:0] arrdiv32_fs529_xor1;
  wire [0:0] arrdiv32_fs529_or0;
  wire [0:0] arrdiv32_fs530_xor1;
  wire [0:0] arrdiv32_fs530_or0;
  wire [0:0] arrdiv32_fs531_xor1;
  wire [0:0] arrdiv32_fs531_or0;
  wire [0:0] arrdiv32_fs532_xor1;
  wire [0:0] arrdiv32_fs532_or0;
  wire [0:0] arrdiv32_fs533_xor1;
  wire [0:0] arrdiv32_fs533_or0;
  wire [0:0] arrdiv32_fs534_xor1;
  wire [0:0] arrdiv32_fs534_or0;
  wire [0:0] arrdiv32_fs535_xor1;
  wire [0:0] arrdiv32_fs535_or0;
  wire [0:0] arrdiv32_fs536_xor1;
  wire [0:0] arrdiv32_fs536_or0;
  wire [0:0] arrdiv32_fs537_xor1;
  wire [0:0] arrdiv32_fs537_or0;
  wire [0:0] arrdiv32_fs538_xor1;
  wire [0:0] arrdiv32_fs538_or0;
  wire [0:0] arrdiv32_fs539_xor1;
  wire [0:0] arrdiv32_fs539_or0;
  wire [0:0] arrdiv32_fs540_xor1;
  wire [0:0] arrdiv32_fs540_or0;
  wire [0:0] arrdiv32_fs541_xor1;
  wire [0:0] arrdiv32_fs541_or0;
  wire [0:0] arrdiv32_fs542_xor1;
  wire [0:0] arrdiv32_fs542_or0;
  wire [0:0] arrdiv32_fs543_xor1;
  wire [0:0] arrdiv32_fs543_or0;
  wire [0:0] arrdiv32_mux2to1496_xor0;
  wire [0:0] arrdiv32_mux2to1497_xor0;
  wire [0:0] arrdiv32_mux2to1498_xor0;
  wire [0:0] arrdiv32_mux2to1499_xor0;
  wire [0:0] arrdiv32_mux2to1500_xor0;
  wire [0:0] arrdiv32_mux2to1501_xor0;
  wire [0:0] arrdiv32_mux2to1502_xor0;
  wire [0:0] arrdiv32_mux2to1503_xor0;
  wire [0:0] arrdiv32_mux2to1504_xor0;
  wire [0:0] arrdiv32_mux2to1505_xor0;
  wire [0:0] arrdiv32_mux2to1506_xor0;
  wire [0:0] arrdiv32_mux2to1507_xor0;
  wire [0:0] arrdiv32_mux2to1508_xor0;
  wire [0:0] arrdiv32_mux2to1509_xor0;
  wire [0:0] arrdiv32_mux2to1510_xor0;
  wire [0:0] arrdiv32_mux2to1511_xor0;
  wire [0:0] arrdiv32_mux2to1512_xor0;
  wire [0:0] arrdiv32_mux2to1513_xor0;
  wire [0:0] arrdiv32_mux2to1514_xor0;
  wire [0:0] arrdiv32_mux2to1515_xor0;
  wire [0:0] arrdiv32_mux2to1516_xor0;
  wire [0:0] arrdiv32_mux2to1517_xor0;
  wire [0:0] arrdiv32_mux2to1518_xor0;
  wire [0:0] arrdiv32_mux2to1519_xor0;
  wire [0:0] arrdiv32_mux2to1520_xor0;
  wire [0:0] arrdiv32_mux2to1521_xor0;
  wire [0:0] arrdiv32_mux2to1522_xor0;
  wire [0:0] arrdiv32_mux2to1523_xor0;
  wire [0:0] arrdiv32_mux2to1524_xor0;
  wire [0:0] arrdiv32_mux2to1525_xor0;
  wire [0:0] arrdiv32_mux2to1526_xor0;
  wire [0:0] arrdiv32_not16;
  wire [0:0] arrdiv32_fs544_xor0;
  wire [0:0] arrdiv32_fs544_and0;
  wire [0:0] arrdiv32_fs545_xor1;
  wire [0:0] arrdiv32_fs545_or0;
  wire [0:0] arrdiv32_fs546_xor1;
  wire [0:0] arrdiv32_fs546_or0;
  wire [0:0] arrdiv32_fs547_xor1;
  wire [0:0] arrdiv32_fs547_or0;
  wire [0:0] arrdiv32_fs548_xor1;
  wire [0:0] arrdiv32_fs548_or0;
  wire [0:0] arrdiv32_fs549_xor1;
  wire [0:0] arrdiv32_fs549_or0;
  wire [0:0] arrdiv32_fs550_xor1;
  wire [0:0] arrdiv32_fs550_or0;
  wire [0:0] arrdiv32_fs551_xor1;
  wire [0:0] arrdiv32_fs551_or0;
  wire [0:0] arrdiv32_fs552_xor1;
  wire [0:0] arrdiv32_fs552_or0;
  wire [0:0] arrdiv32_fs553_xor1;
  wire [0:0] arrdiv32_fs553_or0;
  wire [0:0] arrdiv32_fs554_xor1;
  wire [0:0] arrdiv32_fs554_or0;
  wire [0:0] arrdiv32_fs555_xor1;
  wire [0:0] arrdiv32_fs555_or0;
  wire [0:0] arrdiv32_fs556_xor1;
  wire [0:0] arrdiv32_fs556_or0;
  wire [0:0] arrdiv32_fs557_xor1;
  wire [0:0] arrdiv32_fs557_or0;
  wire [0:0] arrdiv32_fs558_xor1;
  wire [0:0] arrdiv32_fs558_or0;
  wire [0:0] arrdiv32_fs559_xor1;
  wire [0:0] arrdiv32_fs559_or0;
  wire [0:0] arrdiv32_fs560_xor1;
  wire [0:0] arrdiv32_fs560_or0;
  wire [0:0] arrdiv32_fs561_xor1;
  wire [0:0] arrdiv32_fs561_or0;
  wire [0:0] arrdiv32_fs562_xor1;
  wire [0:0] arrdiv32_fs562_or0;
  wire [0:0] arrdiv32_fs563_xor1;
  wire [0:0] arrdiv32_fs563_or0;
  wire [0:0] arrdiv32_fs564_xor1;
  wire [0:0] arrdiv32_fs564_or0;
  wire [0:0] arrdiv32_fs565_xor1;
  wire [0:0] arrdiv32_fs565_or0;
  wire [0:0] arrdiv32_fs566_xor1;
  wire [0:0] arrdiv32_fs566_or0;
  wire [0:0] arrdiv32_fs567_xor1;
  wire [0:0] arrdiv32_fs567_or0;
  wire [0:0] arrdiv32_fs568_xor1;
  wire [0:0] arrdiv32_fs568_or0;
  wire [0:0] arrdiv32_fs569_xor1;
  wire [0:0] arrdiv32_fs569_or0;
  wire [0:0] arrdiv32_fs570_xor1;
  wire [0:0] arrdiv32_fs570_or0;
  wire [0:0] arrdiv32_fs571_xor1;
  wire [0:0] arrdiv32_fs571_or0;
  wire [0:0] arrdiv32_fs572_xor1;
  wire [0:0] arrdiv32_fs572_or0;
  wire [0:0] arrdiv32_fs573_xor1;
  wire [0:0] arrdiv32_fs573_or0;
  wire [0:0] arrdiv32_fs574_xor1;
  wire [0:0] arrdiv32_fs574_or0;
  wire [0:0] arrdiv32_fs575_xor1;
  wire [0:0] arrdiv32_fs575_or0;
  wire [0:0] arrdiv32_mux2to1527_xor0;
  wire [0:0] arrdiv32_mux2to1528_xor0;
  wire [0:0] arrdiv32_mux2to1529_xor0;
  wire [0:0] arrdiv32_mux2to1530_xor0;
  wire [0:0] arrdiv32_mux2to1531_xor0;
  wire [0:0] arrdiv32_mux2to1532_xor0;
  wire [0:0] arrdiv32_mux2to1533_xor0;
  wire [0:0] arrdiv32_mux2to1534_xor0;
  wire [0:0] arrdiv32_mux2to1535_xor0;
  wire [0:0] arrdiv32_mux2to1536_xor0;
  wire [0:0] arrdiv32_mux2to1537_xor0;
  wire [0:0] arrdiv32_mux2to1538_xor0;
  wire [0:0] arrdiv32_mux2to1539_xor0;
  wire [0:0] arrdiv32_mux2to1540_xor0;
  wire [0:0] arrdiv32_mux2to1541_xor0;
  wire [0:0] arrdiv32_mux2to1542_xor0;
  wire [0:0] arrdiv32_mux2to1543_xor0;
  wire [0:0] arrdiv32_mux2to1544_xor0;
  wire [0:0] arrdiv32_mux2to1545_xor0;
  wire [0:0] arrdiv32_mux2to1546_xor0;
  wire [0:0] arrdiv32_mux2to1547_xor0;
  wire [0:0] arrdiv32_mux2to1548_xor0;
  wire [0:0] arrdiv32_mux2to1549_xor0;
  wire [0:0] arrdiv32_mux2to1550_xor0;
  wire [0:0] arrdiv32_mux2to1551_xor0;
  wire [0:0] arrdiv32_mux2to1552_xor0;
  wire [0:0] arrdiv32_mux2to1553_xor0;
  wire [0:0] arrdiv32_mux2to1554_xor0;
  wire [0:0] arrdiv32_mux2to1555_xor0;
  wire [0:0] arrdiv32_mux2to1556_xor0;
  wire [0:0] arrdiv32_mux2to1557_xor0;
  wire [0:0] arrdiv32_not17;
  wire [0:0] arrdiv32_fs576_xor0;
  wire [0:0] arrdiv32_fs576_and0;
  wire [0:0] arrdiv32_fs577_xor1;
  wire [0:0] arrdiv32_fs577_or0;
  wire [0:0] arrdiv32_fs578_xor1;
  wire [0:0] arrdiv32_fs578_or0;
  wire [0:0] arrdiv32_fs579_xor1;
  wire [0:0] arrdiv32_fs579_or0;
  wire [0:0] arrdiv32_fs580_xor1;
  wire [0:0] arrdiv32_fs580_or0;
  wire [0:0] arrdiv32_fs581_xor1;
  wire [0:0] arrdiv32_fs581_or0;
  wire [0:0] arrdiv32_fs582_xor1;
  wire [0:0] arrdiv32_fs582_or0;
  wire [0:0] arrdiv32_fs583_xor1;
  wire [0:0] arrdiv32_fs583_or0;
  wire [0:0] arrdiv32_fs584_xor1;
  wire [0:0] arrdiv32_fs584_or0;
  wire [0:0] arrdiv32_fs585_xor1;
  wire [0:0] arrdiv32_fs585_or0;
  wire [0:0] arrdiv32_fs586_xor1;
  wire [0:0] arrdiv32_fs586_or0;
  wire [0:0] arrdiv32_fs587_xor1;
  wire [0:0] arrdiv32_fs587_or0;
  wire [0:0] arrdiv32_fs588_xor1;
  wire [0:0] arrdiv32_fs588_or0;
  wire [0:0] arrdiv32_fs589_xor1;
  wire [0:0] arrdiv32_fs589_or0;
  wire [0:0] arrdiv32_fs590_xor1;
  wire [0:0] arrdiv32_fs590_or0;
  wire [0:0] arrdiv32_fs591_xor1;
  wire [0:0] arrdiv32_fs591_or0;
  wire [0:0] arrdiv32_fs592_xor1;
  wire [0:0] arrdiv32_fs592_or0;
  wire [0:0] arrdiv32_fs593_xor1;
  wire [0:0] arrdiv32_fs593_or0;
  wire [0:0] arrdiv32_fs594_xor1;
  wire [0:0] arrdiv32_fs594_or0;
  wire [0:0] arrdiv32_fs595_xor1;
  wire [0:0] arrdiv32_fs595_or0;
  wire [0:0] arrdiv32_fs596_xor1;
  wire [0:0] arrdiv32_fs596_or0;
  wire [0:0] arrdiv32_fs597_xor1;
  wire [0:0] arrdiv32_fs597_or0;
  wire [0:0] arrdiv32_fs598_xor1;
  wire [0:0] arrdiv32_fs598_or0;
  wire [0:0] arrdiv32_fs599_xor1;
  wire [0:0] arrdiv32_fs599_or0;
  wire [0:0] arrdiv32_fs600_xor1;
  wire [0:0] arrdiv32_fs600_or0;
  wire [0:0] arrdiv32_fs601_xor1;
  wire [0:0] arrdiv32_fs601_or0;
  wire [0:0] arrdiv32_fs602_xor1;
  wire [0:0] arrdiv32_fs602_or0;
  wire [0:0] arrdiv32_fs603_xor1;
  wire [0:0] arrdiv32_fs603_or0;
  wire [0:0] arrdiv32_fs604_xor1;
  wire [0:0] arrdiv32_fs604_or0;
  wire [0:0] arrdiv32_fs605_xor1;
  wire [0:0] arrdiv32_fs605_or0;
  wire [0:0] arrdiv32_fs606_xor1;
  wire [0:0] arrdiv32_fs606_or0;
  wire [0:0] arrdiv32_fs607_xor1;
  wire [0:0] arrdiv32_fs607_or0;
  wire [0:0] arrdiv32_mux2to1558_xor0;
  wire [0:0] arrdiv32_mux2to1559_xor0;
  wire [0:0] arrdiv32_mux2to1560_xor0;
  wire [0:0] arrdiv32_mux2to1561_xor0;
  wire [0:0] arrdiv32_mux2to1562_xor0;
  wire [0:0] arrdiv32_mux2to1563_xor0;
  wire [0:0] arrdiv32_mux2to1564_xor0;
  wire [0:0] arrdiv32_mux2to1565_xor0;
  wire [0:0] arrdiv32_mux2to1566_xor0;
  wire [0:0] arrdiv32_mux2to1567_xor0;
  wire [0:0] arrdiv32_mux2to1568_xor0;
  wire [0:0] arrdiv32_mux2to1569_xor0;
  wire [0:0] arrdiv32_mux2to1570_xor0;
  wire [0:0] arrdiv32_mux2to1571_xor0;
  wire [0:0] arrdiv32_mux2to1572_xor0;
  wire [0:0] arrdiv32_mux2to1573_xor0;
  wire [0:0] arrdiv32_mux2to1574_xor0;
  wire [0:0] arrdiv32_mux2to1575_xor0;
  wire [0:0] arrdiv32_mux2to1576_xor0;
  wire [0:0] arrdiv32_mux2to1577_xor0;
  wire [0:0] arrdiv32_mux2to1578_xor0;
  wire [0:0] arrdiv32_mux2to1579_xor0;
  wire [0:0] arrdiv32_mux2to1580_xor0;
  wire [0:0] arrdiv32_mux2to1581_xor0;
  wire [0:0] arrdiv32_mux2to1582_xor0;
  wire [0:0] arrdiv32_mux2to1583_xor0;
  wire [0:0] arrdiv32_mux2to1584_xor0;
  wire [0:0] arrdiv32_mux2to1585_xor0;
  wire [0:0] arrdiv32_mux2to1586_xor0;
  wire [0:0] arrdiv32_mux2to1587_xor0;
  wire [0:0] arrdiv32_mux2to1588_xor0;
  wire [0:0] arrdiv32_not18;
  wire [0:0] arrdiv32_fs608_xor0;
  wire [0:0] arrdiv32_fs608_and0;
  wire [0:0] arrdiv32_fs609_xor1;
  wire [0:0] arrdiv32_fs609_or0;
  wire [0:0] arrdiv32_fs610_xor1;
  wire [0:0] arrdiv32_fs610_or0;
  wire [0:0] arrdiv32_fs611_xor1;
  wire [0:0] arrdiv32_fs611_or0;
  wire [0:0] arrdiv32_fs612_xor1;
  wire [0:0] arrdiv32_fs612_or0;
  wire [0:0] arrdiv32_fs613_xor1;
  wire [0:0] arrdiv32_fs613_or0;
  wire [0:0] arrdiv32_fs614_xor1;
  wire [0:0] arrdiv32_fs614_or0;
  wire [0:0] arrdiv32_fs615_xor1;
  wire [0:0] arrdiv32_fs615_or0;
  wire [0:0] arrdiv32_fs616_xor1;
  wire [0:0] arrdiv32_fs616_or0;
  wire [0:0] arrdiv32_fs617_xor1;
  wire [0:0] arrdiv32_fs617_or0;
  wire [0:0] arrdiv32_fs618_xor1;
  wire [0:0] arrdiv32_fs618_or0;
  wire [0:0] arrdiv32_fs619_xor1;
  wire [0:0] arrdiv32_fs619_or0;
  wire [0:0] arrdiv32_fs620_xor1;
  wire [0:0] arrdiv32_fs620_or0;
  wire [0:0] arrdiv32_fs621_xor1;
  wire [0:0] arrdiv32_fs621_or0;
  wire [0:0] arrdiv32_fs622_xor1;
  wire [0:0] arrdiv32_fs622_or0;
  wire [0:0] arrdiv32_fs623_xor1;
  wire [0:0] arrdiv32_fs623_or0;
  wire [0:0] arrdiv32_fs624_xor1;
  wire [0:0] arrdiv32_fs624_or0;
  wire [0:0] arrdiv32_fs625_xor1;
  wire [0:0] arrdiv32_fs625_or0;
  wire [0:0] arrdiv32_fs626_xor1;
  wire [0:0] arrdiv32_fs626_or0;
  wire [0:0] arrdiv32_fs627_xor1;
  wire [0:0] arrdiv32_fs627_or0;
  wire [0:0] arrdiv32_fs628_xor1;
  wire [0:0] arrdiv32_fs628_or0;
  wire [0:0] arrdiv32_fs629_xor1;
  wire [0:0] arrdiv32_fs629_or0;
  wire [0:0] arrdiv32_fs630_xor1;
  wire [0:0] arrdiv32_fs630_or0;
  wire [0:0] arrdiv32_fs631_xor1;
  wire [0:0] arrdiv32_fs631_or0;
  wire [0:0] arrdiv32_fs632_xor1;
  wire [0:0] arrdiv32_fs632_or0;
  wire [0:0] arrdiv32_fs633_xor1;
  wire [0:0] arrdiv32_fs633_or0;
  wire [0:0] arrdiv32_fs634_xor1;
  wire [0:0] arrdiv32_fs634_or0;
  wire [0:0] arrdiv32_fs635_xor1;
  wire [0:0] arrdiv32_fs635_or0;
  wire [0:0] arrdiv32_fs636_xor1;
  wire [0:0] arrdiv32_fs636_or0;
  wire [0:0] arrdiv32_fs637_xor1;
  wire [0:0] arrdiv32_fs637_or0;
  wire [0:0] arrdiv32_fs638_xor1;
  wire [0:0] arrdiv32_fs638_or0;
  wire [0:0] arrdiv32_fs639_xor1;
  wire [0:0] arrdiv32_fs639_or0;
  wire [0:0] arrdiv32_mux2to1589_xor0;
  wire [0:0] arrdiv32_mux2to1590_xor0;
  wire [0:0] arrdiv32_mux2to1591_xor0;
  wire [0:0] arrdiv32_mux2to1592_xor0;
  wire [0:0] arrdiv32_mux2to1593_xor0;
  wire [0:0] arrdiv32_mux2to1594_xor0;
  wire [0:0] arrdiv32_mux2to1595_xor0;
  wire [0:0] arrdiv32_mux2to1596_xor0;
  wire [0:0] arrdiv32_mux2to1597_xor0;
  wire [0:0] arrdiv32_mux2to1598_xor0;
  wire [0:0] arrdiv32_mux2to1599_xor0;
  wire [0:0] arrdiv32_mux2to1600_xor0;
  wire [0:0] arrdiv32_mux2to1601_xor0;
  wire [0:0] arrdiv32_mux2to1602_xor0;
  wire [0:0] arrdiv32_mux2to1603_xor0;
  wire [0:0] arrdiv32_mux2to1604_xor0;
  wire [0:0] arrdiv32_mux2to1605_xor0;
  wire [0:0] arrdiv32_mux2to1606_xor0;
  wire [0:0] arrdiv32_mux2to1607_xor0;
  wire [0:0] arrdiv32_mux2to1608_xor0;
  wire [0:0] arrdiv32_mux2to1609_xor0;
  wire [0:0] arrdiv32_mux2to1610_xor0;
  wire [0:0] arrdiv32_mux2to1611_xor0;
  wire [0:0] arrdiv32_mux2to1612_xor0;
  wire [0:0] arrdiv32_mux2to1613_xor0;
  wire [0:0] arrdiv32_mux2to1614_xor0;
  wire [0:0] arrdiv32_mux2to1615_xor0;
  wire [0:0] arrdiv32_mux2to1616_xor0;
  wire [0:0] arrdiv32_mux2to1617_xor0;
  wire [0:0] arrdiv32_mux2to1618_xor0;
  wire [0:0] arrdiv32_mux2to1619_xor0;
  wire [0:0] arrdiv32_not19;
  wire [0:0] arrdiv32_fs640_xor0;
  wire [0:0] arrdiv32_fs640_and0;
  wire [0:0] arrdiv32_fs641_xor1;
  wire [0:0] arrdiv32_fs641_or0;
  wire [0:0] arrdiv32_fs642_xor1;
  wire [0:0] arrdiv32_fs642_or0;
  wire [0:0] arrdiv32_fs643_xor1;
  wire [0:0] arrdiv32_fs643_or0;
  wire [0:0] arrdiv32_fs644_xor1;
  wire [0:0] arrdiv32_fs644_or0;
  wire [0:0] arrdiv32_fs645_xor1;
  wire [0:0] arrdiv32_fs645_or0;
  wire [0:0] arrdiv32_fs646_xor1;
  wire [0:0] arrdiv32_fs646_or0;
  wire [0:0] arrdiv32_fs647_xor1;
  wire [0:0] arrdiv32_fs647_or0;
  wire [0:0] arrdiv32_fs648_xor1;
  wire [0:0] arrdiv32_fs648_or0;
  wire [0:0] arrdiv32_fs649_xor1;
  wire [0:0] arrdiv32_fs649_or0;
  wire [0:0] arrdiv32_fs650_xor1;
  wire [0:0] arrdiv32_fs650_or0;
  wire [0:0] arrdiv32_fs651_xor1;
  wire [0:0] arrdiv32_fs651_or0;
  wire [0:0] arrdiv32_fs652_xor1;
  wire [0:0] arrdiv32_fs652_or0;
  wire [0:0] arrdiv32_fs653_xor1;
  wire [0:0] arrdiv32_fs653_or0;
  wire [0:0] arrdiv32_fs654_xor1;
  wire [0:0] arrdiv32_fs654_or0;
  wire [0:0] arrdiv32_fs655_xor1;
  wire [0:0] arrdiv32_fs655_or0;
  wire [0:0] arrdiv32_fs656_xor1;
  wire [0:0] arrdiv32_fs656_or0;
  wire [0:0] arrdiv32_fs657_xor1;
  wire [0:0] arrdiv32_fs657_or0;
  wire [0:0] arrdiv32_fs658_xor1;
  wire [0:0] arrdiv32_fs658_or0;
  wire [0:0] arrdiv32_fs659_xor1;
  wire [0:0] arrdiv32_fs659_or0;
  wire [0:0] arrdiv32_fs660_xor1;
  wire [0:0] arrdiv32_fs660_or0;
  wire [0:0] arrdiv32_fs661_xor1;
  wire [0:0] arrdiv32_fs661_or0;
  wire [0:0] arrdiv32_fs662_xor1;
  wire [0:0] arrdiv32_fs662_or0;
  wire [0:0] arrdiv32_fs663_xor1;
  wire [0:0] arrdiv32_fs663_or0;
  wire [0:0] arrdiv32_fs664_xor1;
  wire [0:0] arrdiv32_fs664_or0;
  wire [0:0] arrdiv32_fs665_xor1;
  wire [0:0] arrdiv32_fs665_or0;
  wire [0:0] arrdiv32_fs666_xor1;
  wire [0:0] arrdiv32_fs666_or0;
  wire [0:0] arrdiv32_fs667_xor1;
  wire [0:0] arrdiv32_fs667_or0;
  wire [0:0] arrdiv32_fs668_xor1;
  wire [0:0] arrdiv32_fs668_or0;
  wire [0:0] arrdiv32_fs669_xor1;
  wire [0:0] arrdiv32_fs669_or0;
  wire [0:0] arrdiv32_fs670_xor1;
  wire [0:0] arrdiv32_fs670_or0;
  wire [0:0] arrdiv32_fs671_xor1;
  wire [0:0] arrdiv32_fs671_or0;
  wire [0:0] arrdiv32_mux2to1620_xor0;
  wire [0:0] arrdiv32_mux2to1621_xor0;
  wire [0:0] arrdiv32_mux2to1622_xor0;
  wire [0:0] arrdiv32_mux2to1623_xor0;
  wire [0:0] arrdiv32_mux2to1624_xor0;
  wire [0:0] arrdiv32_mux2to1625_xor0;
  wire [0:0] arrdiv32_mux2to1626_xor0;
  wire [0:0] arrdiv32_mux2to1627_xor0;
  wire [0:0] arrdiv32_mux2to1628_xor0;
  wire [0:0] arrdiv32_mux2to1629_xor0;
  wire [0:0] arrdiv32_mux2to1630_xor0;
  wire [0:0] arrdiv32_mux2to1631_xor0;
  wire [0:0] arrdiv32_mux2to1632_xor0;
  wire [0:0] arrdiv32_mux2to1633_xor0;
  wire [0:0] arrdiv32_mux2to1634_xor0;
  wire [0:0] arrdiv32_mux2to1635_xor0;
  wire [0:0] arrdiv32_mux2to1636_xor0;
  wire [0:0] arrdiv32_mux2to1637_xor0;
  wire [0:0] arrdiv32_mux2to1638_xor0;
  wire [0:0] arrdiv32_mux2to1639_xor0;
  wire [0:0] arrdiv32_mux2to1640_xor0;
  wire [0:0] arrdiv32_mux2to1641_xor0;
  wire [0:0] arrdiv32_mux2to1642_xor0;
  wire [0:0] arrdiv32_mux2to1643_xor0;
  wire [0:0] arrdiv32_mux2to1644_xor0;
  wire [0:0] arrdiv32_mux2to1645_xor0;
  wire [0:0] arrdiv32_mux2to1646_xor0;
  wire [0:0] arrdiv32_mux2to1647_xor0;
  wire [0:0] arrdiv32_mux2to1648_xor0;
  wire [0:0] arrdiv32_mux2to1649_xor0;
  wire [0:0] arrdiv32_mux2to1650_xor0;
  wire [0:0] arrdiv32_not20;
  wire [0:0] arrdiv32_fs672_xor0;
  wire [0:0] arrdiv32_fs672_and0;
  wire [0:0] arrdiv32_fs673_xor1;
  wire [0:0] arrdiv32_fs673_or0;
  wire [0:0] arrdiv32_fs674_xor1;
  wire [0:0] arrdiv32_fs674_or0;
  wire [0:0] arrdiv32_fs675_xor1;
  wire [0:0] arrdiv32_fs675_or0;
  wire [0:0] arrdiv32_fs676_xor1;
  wire [0:0] arrdiv32_fs676_or0;
  wire [0:0] arrdiv32_fs677_xor1;
  wire [0:0] arrdiv32_fs677_or0;
  wire [0:0] arrdiv32_fs678_xor1;
  wire [0:0] arrdiv32_fs678_or0;
  wire [0:0] arrdiv32_fs679_xor1;
  wire [0:0] arrdiv32_fs679_or0;
  wire [0:0] arrdiv32_fs680_xor1;
  wire [0:0] arrdiv32_fs680_or0;
  wire [0:0] arrdiv32_fs681_xor1;
  wire [0:0] arrdiv32_fs681_or0;
  wire [0:0] arrdiv32_fs682_xor1;
  wire [0:0] arrdiv32_fs682_or0;
  wire [0:0] arrdiv32_fs683_xor1;
  wire [0:0] arrdiv32_fs683_or0;
  wire [0:0] arrdiv32_fs684_xor1;
  wire [0:0] arrdiv32_fs684_or0;
  wire [0:0] arrdiv32_fs685_xor1;
  wire [0:0] arrdiv32_fs685_or0;
  wire [0:0] arrdiv32_fs686_xor1;
  wire [0:0] arrdiv32_fs686_or0;
  wire [0:0] arrdiv32_fs687_xor1;
  wire [0:0] arrdiv32_fs687_or0;
  wire [0:0] arrdiv32_fs688_xor1;
  wire [0:0] arrdiv32_fs688_or0;
  wire [0:0] arrdiv32_fs689_xor1;
  wire [0:0] arrdiv32_fs689_or0;
  wire [0:0] arrdiv32_fs690_xor1;
  wire [0:0] arrdiv32_fs690_or0;
  wire [0:0] arrdiv32_fs691_xor1;
  wire [0:0] arrdiv32_fs691_or0;
  wire [0:0] arrdiv32_fs692_xor1;
  wire [0:0] arrdiv32_fs692_or0;
  wire [0:0] arrdiv32_fs693_xor1;
  wire [0:0] arrdiv32_fs693_or0;
  wire [0:0] arrdiv32_fs694_xor1;
  wire [0:0] arrdiv32_fs694_or0;
  wire [0:0] arrdiv32_fs695_xor1;
  wire [0:0] arrdiv32_fs695_or0;
  wire [0:0] arrdiv32_fs696_xor1;
  wire [0:0] arrdiv32_fs696_or0;
  wire [0:0] arrdiv32_fs697_xor1;
  wire [0:0] arrdiv32_fs697_or0;
  wire [0:0] arrdiv32_fs698_xor1;
  wire [0:0] arrdiv32_fs698_or0;
  wire [0:0] arrdiv32_fs699_xor1;
  wire [0:0] arrdiv32_fs699_or0;
  wire [0:0] arrdiv32_fs700_xor1;
  wire [0:0] arrdiv32_fs700_or0;
  wire [0:0] arrdiv32_fs701_xor1;
  wire [0:0] arrdiv32_fs701_or0;
  wire [0:0] arrdiv32_fs702_xor1;
  wire [0:0] arrdiv32_fs702_or0;
  wire [0:0] arrdiv32_fs703_xor1;
  wire [0:0] arrdiv32_fs703_or0;
  wire [0:0] arrdiv32_mux2to1651_xor0;
  wire [0:0] arrdiv32_mux2to1652_xor0;
  wire [0:0] arrdiv32_mux2to1653_xor0;
  wire [0:0] arrdiv32_mux2to1654_xor0;
  wire [0:0] arrdiv32_mux2to1655_xor0;
  wire [0:0] arrdiv32_mux2to1656_xor0;
  wire [0:0] arrdiv32_mux2to1657_xor0;
  wire [0:0] arrdiv32_mux2to1658_xor0;
  wire [0:0] arrdiv32_mux2to1659_xor0;
  wire [0:0] arrdiv32_mux2to1660_xor0;
  wire [0:0] arrdiv32_mux2to1661_xor0;
  wire [0:0] arrdiv32_mux2to1662_xor0;
  wire [0:0] arrdiv32_mux2to1663_xor0;
  wire [0:0] arrdiv32_mux2to1664_xor0;
  wire [0:0] arrdiv32_mux2to1665_xor0;
  wire [0:0] arrdiv32_mux2to1666_xor0;
  wire [0:0] arrdiv32_mux2to1667_xor0;
  wire [0:0] arrdiv32_mux2to1668_xor0;
  wire [0:0] arrdiv32_mux2to1669_xor0;
  wire [0:0] arrdiv32_mux2to1670_xor0;
  wire [0:0] arrdiv32_mux2to1671_xor0;
  wire [0:0] arrdiv32_mux2to1672_xor0;
  wire [0:0] arrdiv32_mux2to1673_xor0;
  wire [0:0] arrdiv32_mux2to1674_xor0;
  wire [0:0] arrdiv32_mux2to1675_xor0;
  wire [0:0] arrdiv32_mux2to1676_xor0;
  wire [0:0] arrdiv32_mux2to1677_xor0;
  wire [0:0] arrdiv32_mux2to1678_xor0;
  wire [0:0] arrdiv32_mux2to1679_xor0;
  wire [0:0] arrdiv32_mux2to1680_xor0;
  wire [0:0] arrdiv32_mux2to1681_xor0;
  wire [0:0] arrdiv32_not21;
  wire [0:0] arrdiv32_fs704_xor0;
  wire [0:0] arrdiv32_fs704_and0;
  wire [0:0] arrdiv32_fs705_xor1;
  wire [0:0] arrdiv32_fs705_or0;
  wire [0:0] arrdiv32_fs706_xor1;
  wire [0:0] arrdiv32_fs706_or0;
  wire [0:0] arrdiv32_fs707_xor1;
  wire [0:0] arrdiv32_fs707_or0;
  wire [0:0] arrdiv32_fs708_xor1;
  wire [0:0] arrdiv32_fs708_or0;
  wire [0:0] arrdiv32_fs709_xor1;
  wire [0:0] arrdiv32_fs709_or0;
  wire [0:0] arrdiv32_fs710_xor1;
  wire [0:0] arrdiv32_fs710_or0;
  wire [0:0] arrdiv32_fs711_xor1;
  wire [0:0] arrdiv32_fs711_or0;
  wire [0:0] arrdiv32_fs712_xor1;
  wire [0:0] arrdiv32_fs712_or0;
  wire [0:0] arrdiv32_fs713_xor1;
  wire [0:0] arrdiv32_fs713_or0;
  wire [0:0] arrdiv32_fs714_xor1;
  wire [0:0] arrdiv32_fs714_or0;
  wire [0:0] arrdiv32_fs715_xor1;
  wire [0:0] arrdiv32_fs715_or0;
  wire [0:0] arrdiv32_fs716_xor1;
  wire [0:0] arrdiv32_fs716_or0;
  wire [0:0] arrdiv32_fs717_xor1;
  wire [0:0] arrdiv32_fs717_or0;
  wire [0:0] arrdiv32_fs718_xor1;
  wire [0:0] arrdiv32_fs718_or0;
  wire [0:0] arrdiv32_fs719_xor1;
  wire [0:0] arrdiv32_fs719_or0;
  wire [0:0] arrdiv32_fs720_xor1;
  wire [0:0] arrdiv32_fs720_or0;
  wire [0:0] arrdiv32_fs721_xor1;
  wire [0:0] arrdiv32_fs721_or0;
  wire [0:0] arrdiv32_fs722_xor1;
  wire [0:0] arrdiv32_fs722_or0;
  wire [0:0] arrdiv32_fs723_xor1;
  wire [0:0] arrdiv32_fs723_or0;
  wire [0:0] arrdiv32_fs724_xor1;
  wire [0:0] arrdiv32_fs724_or0;
  wire [0:0] arrdiv32_fs725_xor1;
  wire [0:0] arrdiv32_fs725_or0;
  wire [0:0] arrdiv32_fs726_xor1;
  wire [0:0] arrdiv32_fs726_or0;
  wire [0:0] arrdiv32_fs727_xor1;
  wire [0:0] arrdiv32_fs727_or0;
  wire [0:0] arrdiv32_fs728_xor1;
  wire [0:0] arrdiv32_fs728_or0;
  wire [0:0] arrdiv32_fs729_xor1;
  wire [0:0] arrdiv32_fs729_or0;
  wire [0:0] arrdiv32_fs730_xor1;
  wire [0:0] arrdiv32_fs730_or0;
  wire [0:0] arrdiv32_fs731_xor1;
  wire [0:0] arrdiv32_fs731_or0;
  wire [0:0] arrdiv32_fs732_xor1;
  wire [0:0] arrdiv32_fs732_or0;
  wire [0:0] arrdiv32_fs733_xor1;
  wire [0:0] arrdiv32_fs733_or0;
  wire [0:0] arrdiv32_fs734_xor1;
  wire [0:0] arrdiv32_fs734_or0;
  wire [0:0] arrdiv32_fs735_xor1;
  wire [0:0] arrdiv32_fs735_or0;
  wire [0:0] arrdiv32_mux2to1682_xor0;
  wire [0:0] arrdiv32_mux2to1683_xor0;
  wire [0:0] arrdiv32_mux2to1684_xor0;
  wire [0:0] arrdiv32_mux2to1685_xor0;
  wire [0:0] arrdiv32_mux2to1686_xor0;
  wire [0:0] arrdiv32_mux2to1687_xor0;
  wire [0:0] arrdiv32_mux2to1688_xor0;
  wire [0:0] arrdiv32_mux2to1689_xor0;
  wire [0:0] arrdiv32_mux2to1690_xor0;
  wire [0:0] arrdiv32_mux2to1691_xor0;
  wire [0:0] arrdiv32_mux2to1692_xor0;
  wire [0:0] arrdiv32_mux2to1693_xor0;
  wire [0:0] arrdiv32_mux2to1694_xor0;
  wire [0:0] arrdiv32_mux2to1695_xor0;
  wire [0:0] arrdiv32_mux2to1696_xor0;
  wire [0:0] arrdiv32_mux2to1697_xor0;
  wire [0:0] arrdiv32_mux2to1698_xor0;
  wire [0:0] arrdiv32_mux2to1699_xor0;
  wire [0:0] arrdiv32_mux2to1700_xor0;
  wire [0:0] arrdiv32_mux2to1701_xor0;
  wire [0:0] arrdiv32_mux2to1702_xor0;
  wire [0:0] arrdiv32_mux2to1703_xor0;
  wire [0:0] arrdiv32_mux2to1704_xor0;
  wire [0:0] arrdiv32_mux2to1705_xor0;
  wire [0:0] arrdiv32_mux2to1706_xor0;
  wire [0:0] arrdiv32_mux2to1707_xor0;
  wire [0:0] arrdiv32_mux2to1708_xor0;
  wire [0:0] arrdiv32_mux2to1709_xor0;
  wire [0:0] arrdiv32_mux2to1710_xor0;
  wire [0:0] arrdiv32_mux2to1711_xor0;
  wire [0:0] arrdiv32_mux2to1712_xor0;
  wire [0:0] arrdiv32_not22;
  wire [0:0] arrdiv32_fs736_xor0;
  wire [0:0] arrdiv32_fs736_and0;
  wire [0:0] arrdiv32_fs737_xor1;
  wire [0:0] arrdiv32_fs737_or0;
  wire [0:0] arrdiv32_fs738_xor1;
  wire [0:0] arrdiv32_fs738_or0;
  wire [0:0] arrdiv32_fs739_xor1;
  wire [0:0] arrdiv32_fs739_or0;
  wire [0:0] arrdiv32_fs740_xor1;
  wire [0:0] arrdiv32_fs740_or0;
  wire [0:0] arrdiv32_fs741_xor1;
  wire [0:0] arrdiv32_fs741_or0;
  wire [0:0] arrdiv32_fs742_xor1;
  wire [0:0] arrdiv32_fs742_or0;
  wire [0:0] arrdiv32_fs743_xor1;
  wire [0:0] arrdiv32_fs743_or0;
  wire [0:0] arrdiv32_fs744_xor1;
  wire [0:0] arrdiv32_fs744_or0;
  wire [0:0] arrdiv32_fs745_xor1;
  wire [0:0] arrdiv32_fs745_or0;
  wire [0:0] arrdiv32_fs746_xor1;
  wire [0:0] arrdiv32_fs746_or0;
  wire [0:0] arrdiv32_fs747_xor1;
  wire [0:0] arrdiv32_fs747_or0;
  wire [0:0] arrdiv32_fs748_xor1;
  wire [0:0] arrdiv32_fs748_or0;
  wire [0:0] arrdiv32_fs749_xor1;
  wire [0:0] arrdiv32_fs749_or0;
  wire [0:0] arrdiv32_fs750_xor1;
  wire [0:0] arrdiv32_fs750_or0;
  wire [0:0] arrdiv32_fs751_xor1;
  wire [0:0] arrdiv32_fs751_or0;
  wire [0:0] arrdiv32_fs752_xor1;
  wire [0:0] arrdiv32_fs752_or0;
  wire [0:0] arrdiv32_fs753_xor1;
  wire [0:0] arrdiv32_fs753_or0;
  wire [0:0] arrdiv32_fs754_xor1;
  wire [0:0] arrdiv32_fs754_or0;
  wire [0:0] arrdiv32_fs755_xor1;
  wire [0:0] arrdiv32_fs755_or0;
  wire [0:0] arrdiv32_fs756_xor1;
  wire [0:0] arrdiv32_fs756_or0;
  wire [0:0] arrdiv32_fs757_xor1;
  wire [0:0] arrdiv32_fs757_or0;
  wire [0:0] arrdiv32_fs758_xor1;
  wire [0:0] arrdiv32_fs758_or0;
  wire [0:0] arrdiv32_fs759_xor1;
  wire [0:0] arrdiv32_fs759_or0;
  wire [0:0] arrdiv32_fs760_xor1;
  wire [0:0] arrdiv32_fs760_or0;
  wire [0:0] arrdiv32_fs761_xor1;
  wire [0:0] arrdiv32_fs761_or0;
  wire [0:0] arrdiv32_fs762_xor1;
  wire [0:0] arrdiv32_fs762_or0;
  wire [0:0] arrdiv32_fs763_xor1;
  wire [0:0] arrdiv32_fs763_or0;
  wire [0:0] arrdiv32_fs764_xor1;
  wire [0:0] arrdiv32_fs764_or0;
  wire [0:0] arrdiv32_fs765_xor1;
  wire [0:0] arrdiv32_fs765_or0;
  wire [0:0] arrdiv32_fs766_xor1;
  wire [0:0] arrdiv32_fs766_or0;
  wire [0:0] arrdiv32_fs767_xor1;
  wire [0:0] arrdiv32_fs767_or0;
  wire [0:0] arrdiv32_mux2to1713_xor0;
  wire [0:0] arrdiv32_mux2to1714_xor0;
  wire [0:0] arrdiv32_mux2to1715_xor0;
  wire [0:0] arrdiv32_mux2to1716_xor0;
  wire [0:0] arrdiv32_mux2to1717_xor0;
  wire [0:0] arrdiv32_mux2to1718_xor0;
  wire [0:0] arrdiv32_mux2to1719_xor0;
  wire [0:0] arrdiv32_mux2to1720_xor0;
  wire [0:0] arrdiv32_mux2to1721_xor0;
  wire [0:0] arrdiv32_mux2to1722_xor0;
  wire [0:0] arrdiv32_mux2to1723_xor0;
  wire [0:0] arrdiv32_mux2to1724_xor0;
  wire [0:0] arrdiv32_mux2to1725_xor0;
  wire [0:0] arrdiv32_mux2to1726_xor0;
  wire [0:0] arrdiv32_mux2to1727_xor0;
  wire [0:0] arrdiv32_mux2to1728_xor0;
  wire [0:0] arrdiv32_mux2to1729_xor0;
  wire [0:0] arrdiv32_mux2to1730_xor0;
  wire [0:0] arrdiv32_mux2to1731_xor0;
  wire [0:0] arrdiv32_mux2to1732_xor0;
  wire [0:0] arrdiv32_mux2to1733_xor0;
  wire [0:0] arrdiv32_mux2to1734_xor0;
  wire [0:0] arrdiv32_mux2to1735_xor0;
  wire [0:0] arrdiv32_mux2to1736_xor0;
  wire [0:0] arrdiv32_mux2to1737_xor0;
  wire [0:0] arrdiv32_mux2to1738_xor0;
  wire [0:0] arrdiv32_mux2to1739_xor0;
  wire [0:0] arrdiv32_mux2to1740_xor0;
  wire [0:0] arrdiv32_mux2to1741_xor0;
  wire [0:0] arrdiv32_mux2to1742_xor0;
  wire [0:0] arrdiv32_mux2to1743_xor0;
  wire [0:0] arrdiv32_not23;
  wire [0:0] arrdiv32_fs768_xor0;
  wire [0:0] arrdiv32_fs768_and0;
  wire [0:0] arrdiv32_fs769_xor1;
  wire [0:0] arrdiv32_fs769_or0;
  wire [0:0] arrdiv32_fs770_xor1;
  wire [0:0] arrdiv32_fs770_or0;
  wire [0:0] arrdiv32_fs771_xor1;
  wire [0:0] arrdiv32_fs771_or0;
  wire [0:0] arrdiv32_fs772_xor1;
  wire [0:0] arrdiv32_fs772_or0;
  wire [0:0] arrdiv32_fs773_xor1;
  wire [0:0] arrdiv32_fs773_or0;
  wire [0:0] arrdiv32_fs774_xor1;
  wire [0:0] arrdiv32_fs774_or0;
  wire [0:0] arrdiv32_fs775_xor1;
  wire [0:0] arrdiv32_fs775_or0;
  wire [0:0] arrdiv32_fs776_xor1;
  wire [0:0] arrdiv32_fs776_or0;
  wire [0:0] arrdiv32_fs777_xor1;
  wire [0:0] arrdiv32_fs777_or0;
  wire [0:0] arrdiv32_fs778_xor1;
  wire [0:0] arrdiv32_fs778_or0;
  wire [0:0] arrdiv32_fs779_xor1;
  wire [0:0] arrdiv32_fs779_or0;
  wire [0:0] arrdiv32_fs780_xor1;
  wire [0:0] arrdiv32_fs780_or0;
  wire [0:0] arrdiv32_fs781_xor1;
  wire [0:0] arrdiv32_fs781_or0;
  wire [0:0] arrdiv32_fs782_xor1;
  wire [0:0] arrdiv32_fs782_or0;
  wire [0:0] arrdiv32_fs783_xor1;
  wire [0:0] arrdiv32_fs783_or0;
  wire [0:0] arrdiv32_fs784_xor1;
  wire [0:0] arrdiv32_fs784_or0;
  wire [0:0] arrdiv32_fs785_xor1;
  wire [0:0] arrdiv32_fs785_or0;
  wire [0:0] arrdiv32_fs786_xor1;
  wire [0:0] arrdiv32_fs786_or0;
  wire [0:0] arrdiv32_fs787_xor1;
  wire [0:0] arrdiv32_fs787_or0;
  wire [0:0] arrdiv32_fs788_xor1;
  wire [0:0] arrdiv32_fs788_or0;
  wire [0:0] arrdiv32_fs789_xor1;
  wire [0:0] arrdiv32_fs789_or0;
  wire [0:0] arrdiv32_fs790_xor1;
  wire [0:0] arrdiv32_fs790_or0;
  wire [0:0] arrdiv32_fs791_xor1;
  wire [0:0] arrdiv32_fs791_or0;
  wire [0:0] arrdiv32_fs792_xor1;
  wire [0:0] arrdiv32_fs792_or0;
  wire [0:0] arrdiv32_fs793_xor1;
  wire [0:0] arrdiv32_fs793_or0;
  wire [0:0] arrdiv32_fs794_xor1;
  wire [0:0] arrdiv32_fs794_or0;
  wire [0:0] arrdiv32_fs795_xor1;
  wire [0:0] arrdiv32_fs795_or0;
  wire [0:0] arrdiv32_fs796_xor1;
  wire [0:0] arrdiv32_fs796_or0;
  wire [0:0] arrdiv32_fs797_xor1;
  wire [0:0] arrdiv32_fs797_or0;
  wire [0:0] arrdiv32_fs798_xor1;
  wire [0:0] arrdiv32_fs798_or0;
  wire [0:0] arrdiv32_fs799_xor1;
  wire [0:0] arrdiv32_fs799_or0;
  wire [0:0] arrdiv32_mux2to1744_xor0;
  wire [0:0] arrdiv32_mux2to1745_xor0;
  wire [0:0] arrdiv32_mux2to1746_xor0;
  wire [0:0] arrdiv32_mux2to1747_xor0;
  wire [0:0] arrdiv32_mux2to1748_xor0;
  wire [0:0] arrdiv32_mux2to1749_xor0;
  wire [0:0] arrdiv32_mux2to1750_xor0;
  wire [0:0] arrdiv32_mux2to1751_xor0;
  wire [0:0] arrdiv32_mux2to1752_xor0;
  wire [0:0] arrdiv32_mux2to1753_xor0;
  wire [0:0] arrdiv32_mux2to1754_xor0;
  wire [0:0] arrdiv32_mux2to1755_xor0;
  wire [0:0] arrdiv32_mux2to1756_xor0;
  wire [0:0] arrdiv32_mux2to1757_xor0;
  wire [0:0] arrdiv32_mux2to1758_xor0;
  wire [0:0] arrdiv32_mux2to1759_xor0;
  wire [0:0] arrdiv32_mux2to1760_xor0;
  wire [0:0] arrdiv32_mux2to1761_xor0;
  wire [0:0] arrdiv32_mux2to1762_xor0;
  wire [0:0] arrdiv32_mux2to1763_xor0;
  wire [0:0] arrdiv32_mux2to1764_xor0;
  wire [0:0] arrdiv32_mux2to1765_xor0;
  wire [0:0] arrdiv32_mux2to1766_xor0;
  wire [0:0] arrdiv32_mux2to1767_xor0;
  wire [0:0] arrdiv32_mux2to1768_xor0;
  wire [0:0] arrdiv32_mux2to1769_xor0;
  wire [0:0] arrdiv32_mux2to1770_xor0;
  wire [0:0] arrdiv32_mux2to1771_xor0;
  wire [0:0] arrdiv32_mux2to1772_xor0;
  wire [0:0] arrdiv32_mux2to1773_xor0;
  wire [0:0] arrdiv32_mux2to1774_xor0;
  wire [0:0] arrdiv32_not24;
  wire [0:0] arrdiv32_fs800_xor0;
  wire [0:0] arrdiv32_fs800_and0;
  wire [0:0] arrdiv32_fs801_xor1;
  wire [0:0] arrdiv32_fs801_or0;
  wire [0:0] arrdiv32_fs802_xor1;
  wire [0:0] arrdiv32_fs802_or0;
  wire [0:0] arrdiv32_fs803_xor1;
  wire [0:0] arrdiv32_fs803_or0;
  wire [0:0] arrdiv32_fs804_xor1;
  wire [0:0] arrdiv32_fs804_or0;
  wire [0:0] arrdiv32_fs805_xor1;
  wire [0:0] arrdiv32_fs805_or0;
  wire [0:0] arrdiv32_fs806_xor1;
  wire [0:0] arrdiv32_fs806_or0;
  wire [0:0] arrdiv32_fs807_xor1;
  wire [0:0] arrdiv32_fs807_or0;
  wire [0:0] arrdiv32_fs808_xor1;
  wire [0:0] arrdiv32_fs808_or0;
  wire [0:0] arrdiv32_fs809_xor1;
  wire [0:0] arrdiv32_fs809_or0;
  wire [0:0] arrdiv32_fs810_xor1;
  wire [0:0] arrdiv32_fs810_or0;
  wire [0:0] arrdiv32_fs811_xor1;
  wire [0:0] arrdiv32_fs811_or0;
  wire [0:0] arrdiv32_fs812_xor1;
  wire [0:0] arrdiv32_fs812_or0;
  wire [0:0] arrdiv32_fs813_xor1;
  wire [0:0] arrdiv32_fs813_or0;
  wire [0:0] arrdiv32_fs814_xor1;
  wire [0:0] arrdiv32_fs814_or0;
  wire [0:0] arrdiv32_fs815_xor1;
  wire [0:0] arrdiv32_fs815_or0;
  wire [0:0] arrdiv32_fs816_xor1;
  wire [0:0] arrdiv32_fs816_or0;
  wire [0:0] arrdiv32_fs817_xor1;
  wire [0:0] arrdiv32_fs817_or0;
  wire [0:0] arrdiv32_fs818_xor1;
  wire [0:0] arrdiv32_fs818_or0;
  wire [0:0] arrdiv32_fs819_xor1;
  wire [0:0] arrdiv32_fs819_or0;
  wire [0:0] arrdiv32_fs820_xor1;
  wire [0:0] arrdiv32_fs820_or0;
  wire [0:0] arrdiv32_fs821_xor1;
  wire [0:0] arrdiv32_fs821_or0;
  wire [0:0] arrdiv32_fs822_xor1;
  wire [0:0] arrdiv32_fs822_or0;
  wire [0:0] arrdiv32_fs823_xor1;
  wire [0:0] arrdiv32_fs823_or0;
  wire [0:0] arrdiv32_fs824_xor1;
  wire [0:0] arrdiv32_fs824_or0;
  wire [0:0] arrdiv32_fs825_xor1;
  wire [0:0] arrdiv32_fs825_or0;
  wire [0:0] arrdiv32_fs826_xor1;
  wire [0:0] arrdiv32_fs826_or0;
  wire [0:0] arrdiv32_fs827_xor1;
  wire [0:0] arrdiv32_fs827_or0;
  wire [0:0] arrdiv32_fs828_xor1;
  wire [0:0] arrdiv32_fs828_or0;
  wire [0:0] arrdiv32_fs829_xor1;
  wire [0:0] arrdiv32_fs829_or0;
  wire [0:0] arrdiv32_fs830_xor1;
  wire [0:0] arrdiv32_fs830_or0;
  wire [0:0] arrdiv32_fs831_xor1;
  wire [0:0] arrdiv32_fs831_or0;
  wire [0:0] arrdiv32_mux2to1775_xor0;
  wire [0:0] arrdiv32_mux2to1776_xor0;
  wire [0:0] arrdiv32_mux2to1777_xor0;
  wire [0:0] arrdiv32_mux2to1778_xor0;
  wire [0:0] arrdiv32_mux2to1779_xor0;
  wire [0:0] arrdiv32_mux2to1780_xor0;
  wire [0:0] arrdiv32_mux2to1781_xor0;
  wire [0:0] arrdiv32_mux2to1782_xor0;
  wire [0:0] arrdiv32_mux2to1783_xor0;
  wire [0:0] arrdiv32_mux2to1784_xor0;
  wire [0:0] arrdiv32_mux2to1785_xor0;
  wire [0:0] arrdiv32_mux2to1786_xor0;
  wire [0:0] arrdiv32_mux2to1787_xor0;
  wire [0:0] arrdiv32_mux2to1788_xor0;
  wire [0:0] arrdiv32_mux2to1789_xor0;
  wire [0:0] arrdiv32_mux2to1790_xor0;
  wire [0:0] arrdiv32_mux2to1791_xor0;
  wire [0:0] arrdiv32_mux2to1792_xor0;
  wire [0:0] arrdiv32_mux2to1793_xor0;
  wire [0:0] arrdiv32_mux2to1794_xor0;
  wire [0:0] arrdiv32_mux2to1795_xor0;
  wire [0:0] arrdiv32_mux2to1796_xor0;
  wire [0:0] arrdiv32_mux2to1797_xor0;
  wire [0:0] arrdiv32_mux2to1798_xor0;
  wire [0:0] arrdiv32_mux2to1799_xor0;
  wire [0:0] arrdiv32_mux2to1800_xor0;
  wire [0:0] arrdiv32_mux2to1801_xor0;
  wire [0:0] arrdiv32_mux2to1802_xor0;
  wire [0:0] arrdiv32_mux2to1803_xor0;
  wire [0:0] arrdiv32_mux2to1804_xor0;
  wire [0:0] arrdiv32_mux2to1805_xor0;
  wire [0:0] arrdiv32_not25;
  wire [0:0] arrdiv32_fs832_xor0;
  wire [0:0] arrdiv32_fs832_and0;
  wire [0:0] arrdiv32_fs833_xor1;
  wire [0:0] arrdiv32_fs833_or0;
  wire [0:0] arrdiv32_fs834_xor1;
  wire [0:0] arrdiv32_fs834_or0;
  wire [0:0] arrdiv32_fs835_xor1;
  wire [0:0] arrdiv32_fs835_or0;
  wire [0:0] arrdiv32_fs836_xor1;
  wire [0:0] arrdiv32_fs836_or0;
  wire [0:0] arrdiv32_fs837_xor1;
  wire [0:0] arrdiv32_fs837_or0;
  wire [0:0] arrdiv32_fs838_xor1;
  wire [0:0] arrdiv32_fs838_or0;
  wire [0:0] arrdiv32_fs839_xor1;
  wire [0:0] arrdiv32_fs839_or0;
  wire [0:0] arrdiv32_fs840_xor1;
  wire [0:0] arrdiv32_fs840_or0;
  wire [0:0] arrdiv32_fs841_xor1;
  wire [0:0] arrdiv32_fs841_or0;
  wire [0:0] arrdiv32_fs842_xor1;
  wire [0:0] arrdiv32_fs842_or0;
  wire [0:0] arrdiv32_fs843_xor1;
  wire [0:0] arrdiv32_fs843_or0;
  wire [0:0] arrdiv32_fs844_xor1;
  wire [0:0] arrdiv32_fs844_or0;
  wire [0:0] arrdiv32_fs845_xor1;
  wire [0:0] arrdiv32_fs845_or0;
  wire [0:0] arrdiv32_fs846_xor1;
  wire [0:0] arrdiv32_fs846_or0;
  wire [0:0] arrdiv32_fs847_xor1;
  wire [0:0] arrdiv32_fs847_or0;
  wire [0:0] arrdiv32_fs848_xor1;
  wire [0:0] arrdiv32_fs848_or0;
  wire [0:0] arrdiv32_fs849_xor1;
  wire [0:0] arrdiv32_fs849_or0;
  wire [0:0] arrdiv32_fs850_xor1;
  wire [0:0] arrdiv32_fs850_or0;
  wire [0:0] arrdiv32_fs851_xor1;
  wire [0:0] arrdiv32_fs851_or0;
  wire [0:0] arrdiv32_fs852_xor1;
  wire [0:0] arrdiv32_fs852_or0;
  wire [0:0] arrdiv32_fs853_xor1;
  wire [0:0] arrdiv32_fs853_or0;
  wire [0:0] arrdiv32_fs854_xor1;
  wire [0:0] arrdiv32_fs854_or0;
  wire [0:0] arrdiv32_fs855_xor1;
  wire [0:0] arrdiv32_fs855_or0;
  wire [0:0] arrdiv32_fs856_xor1;
  wire [0:0] arrdiv32_fs856_or0;
  wire [0:0] arrdiv32_fs857_xor1;
  wire [0:0] arrdiv32_fs857_or0;
  wire [0:0] arrdiv32_fs858_xor1;
  wire [0:0] arrdiv32_fs858_or0;
  wire [0:0] arrdiv32_fs859_xor1;
  wire [0:0] arrdiv32_fs859_or0;
  wire [0:0] arrdiv32_fs860_xor1;
  wire [0:0] arrdiv32_fs860_or0;
  wire [0:0] arrdiv32_fs861_xor1;
  wire [0:0] arrdiv32_fs861_or0;
  wire [0:0] arrdiv32_fs862_xor1;
  wire [0:0] arrdiv32_fs862_or0;
  wire [0:0] arrdiv32_fs863_xor1;
  wire [0:0] arrdiv32_fs863_or0;
  wire [0:0] arrdiv32_mux2to1806_xor0;
  wire [0:0] arrdiv32_mux2to1807_xor0;
  wire [0:0] arrdiv32_mux2to1808_xor0;
  wire [0:0] arrdiv32_mux2to1809_xor0;
  wire [0:0] arrdiv32_mux2to1810_xor0;
  wire [0:0] arrdiv32_mux2to1811_xor0;
  wire [0:0] arrdiv32_mux2to1812_xor0;
  wire [0:0] arrdiv32_mux2to1813_xor0;
  wire [0:0] arrdiv32_mux2to1814_xor0;
  wire [0:0] arrdiv32_mux2to1815_xor0;
  wire [0:0] arrdiv32_mux2to1816_xor0;
  wire [0:0] arrdiv32_mux2to1817_xor0;
  wire [0:0] arrdiv32_mux2to1818_xor0;
  wire [0:0] arrdiv32_mux2to1819_xor0;
  wire [0:0] arrdiv32_mux2to1820_xor0;
  wire [0:0] arrdiv32_mux2to1821_xor0;
  wire [0:0] arrdiv32_mux2to1822_xor0;
  wire [0:0] arrdiv32_mux2to1823_xor0;
  wire [0:0] arrdiv32_mux2to1824_xor0;
  wire [0:0] arrdiv32_mux2to1825_xor0;
  wire [0:0] arrdiv32_mux2to1826_xor0;
  wire [0:0] arrdiv32_mux2to1827_xor0;
  wire [0:0] arrdiv32_mux2to1828_xor0;
  wire [0:0] arrdiv32_mux2to1829_xor0;
  wire [0:0] arrdiv32_mux2to1830_xor0;
  wire [0:0] arrdiv32_mux2to1831_xor0;
  wire [0:0] arrdiv32_mux2to1832_xor0;
  wire [0:0] arrdiv32_mux2to1833_xor0;
  wire [0:0] arrdiv32_mux2to1834_xor0;
  wire [0:0] arrdiv32_mux2to1835_xor0;
  wire [0:0] arrdiv32_mux2to1836_xor0;
  wire [0:0] arrdiv32_not26;
  wire [0:0] arrdiv32_fs864_xor0;
  wire [0:0] arrdiv32_fs864_and0;
  wire [0:0] arrdiv32_fs865_xor1;
  wire [0:0] arrdiv32_fs865_or0;
  wire [0:0] arrdiv32_fs866_xor1;
  wire [0:0] arrdiv32_fs866_or0;
  wire [0:0] arrdiv32_fs867_xor1;
  wire [0:0] arrdiv32_fs867_or0;
  wire [0:0] arrdiv32_fs868_xor1;
  wire [0:0] arrdiv32_fs868_or0;
  wire [0:0] arrdiv32_fs869_xor1;
  wire [0:0] arrdiv32_fs869_or0;
  wire [0:0] arrdiv32_fs870_xor1;
  wire [0:0] arrdiv32_fs870_or0;
  wire [0:0] arrdiv32_fs871_xor1;
  wire [0:0] arrdiv32_fs871_or0;
  wire [0:0] arrdiv32_fs872_xor1;
  wire [0:0] arrdiv32_fs872_or0;
  wire [0:0] arrdiv32_fs873_xor1;
  wire [0:0] arrdiv32_fs873_or0;
  wire [0:0] arrdiv32_fs874_xor1;
  wire [0:0] arrdiv32_fs874_or0;
  wire [0:0] arrdiv32_fs875_xor1;
  wire [0:0] arrdiv32_fs875_or0;
  wire [0:0] arrdiv32_fs876_xor1;
  wire [0:0] arrdiv32_fs876_or0;
  wire [0:0] arrdiv32_fs877_xor1;
  wire [0:0] arrdiv32_fs877_or0;
  wire [0:0] arrdiv32_fs878_xor1;
  wire [0:0] arrdiv32_fs878_or0;
  wire [0:0] arrdiv32_fs879_xor1;
  wire [0:0] arrdiv32_fs879_or0;
  wire [0:0] arrdiv32_fs880_xor1;
  wire [0:0] arrdiv32_fs880_or0;
  wire [0:0] arrdiv32_fs881_xor1;
  wire [0:0] arrdiv32_fs881_or0;
  wire [0:0] arrdiv32_fs882_xor1;
  wire [0:0] arrdiv32_fs882_or0;
  wire [0:0] arrdiv32_fs883_xor1;
  wire [0:0] arrdiv32_fs883_or0;
  wire [0:0] arrdiv32_fs884_xor1;
  wire [0:0] arrdiv32_fs884_or0;
  wire [0:0] arrdiv32_fs885_xor1;
  wire [0:0] arrdiv32_fs885_or0;
  wire [0:0] arrdiv32_fs886_xor1;
  wire [0:0] arrdiv32_fs886_or0;
  wire [0:0] arrdiv32_fs887_xor1;
  wire [0:0] arrdiv32_fs887_or0;
  wire [0:0] arrdiv32_fs888_xor1;
  wire [0:0] arrdiv32_fs888_or0;
  wire [0:0] arrdiv32_fs889_xor1;
  wire [0:0] arrdiv32_fs889_or0;
  wire [0:0] arrdiv32_fs890_xor1;
  wire [0:0] arrdiv32_fs890_or0;
  wire [0:0] arrdiv32_fs891_xor1;
  wire [0:0] arrdiv32_fs891_or0;
  wire [0:0] arrdiv32_fs892_xor1;
  wire [0:0] arrdiv32_fs892_or0;
  wire [0:0] arrdiv32_fs893_xor1;
  wire [0:0] arrdiv32_fs893_or0;
  wire [0:0] arrdiv32_fs894_xor1;
  wire [0:0] arrdiv32_fs894_or0;
  wire [0:0] arrdiv32_fs895_xor1;
  wire [0:0] arrdiv32_fs895_or0;
  wire [0:0] arrdiv32_mux2to1837_xor0;
  wire [0:0] arrdiv32_mux2to1838_xor0;
  wire [0:0] arrdiv32_mux2to1839_xor0;
  wire [0:0] arrdiv32_mux2to1840_xor0;
  wire [0:0] arrdiv32_mux2to1841_xor0;
  wire [0:0] arrdiv32_mux2to1842_xor0;
  wire [0:0] arrdiv32_mux2to1843_xor0;
  wire [0:0] arrdiv32_mux2to1844_xor0;
  wire [0:0] arrdiv32_mux2to1845_xor0;
  wire [0:0] arrdiv32_mux2to1846_xor0;
  wire [0:0] arrdiv32_mux2to1847_xor0;
  wire [0:0] arrdiv32_mux2to1848_xor0;
  wire [0:0] arrdiv32_mux2to1849_xor0;
  wire [0:0] arrdiv32_mux2to1850_xor0;
  wire [0:0] arrdiv32_mux2to1851_xor0;
  wire [0:0] arrdiv32_mux2to1852_xor0;
  wire [0:0] arrdiv32_mux2to1853_xor0;
  wire [0:0] arrdiv32_mux2to1854_xor0;
  wire [0:0] arrdiv32_mux2to1855_xor0;
  wire [0:0] arrdiv32_mux2to1856_xor0;
  wire [0:0] arrdiv32_mux2to1857_xor0;
  wire [0:0] arrdiv32_mux2to1858_xor0;
  wire [0:0] arrdiv32_mux2to1859_xor0;
  wire [0:0] arrdiv32_mux2to1860_xor0;
  wire [0:0] arrdiv32_mux2to1861_xor0;
  wire [0:0] arrdiv32_mux2to1862_xor0;
  wire [0:0] arrdiv32_mux2to1863_xor0;
  wire [0:0] arrdiv32_mux2to1864_xor0;
  wire [0:0] arrdiv32_mux2to1865_xor0;
  wire [0:0] arrdiv32_mux2to1866_xor0;
  wire [0:0] arrdiv32_mux2to1867_xor0;
  wire [0:0] arrdiv32_not27;
  wire [0:0] arrdiv32_fs896_xor0;
  wire [0:0] arrdiv32_fs896_and0;
  wire [0:0] arrdiv32_fs897_xor1;
  wire [0:0] arrdiv32_fs897_or0;
  wire [0:0] arrdiv32_fs898_xor1;
  wire [0:0] arrdiv32_fs898_or0;
  wire [0:0] arrdiv32_fs899_xor1;
  wire [0:0] arrdiv32_fs899_or0;
  wire [0:0] arrdiv32_fs900_xor1;
  wire [0:0] arrdiv32_fs900_or0;
  wire [0:0] arrdiv32_fs901_xor1;
  wire [0:0] arrdiv32_fs901_or0;
  wire [0:0] arrdiv32_fs902_xor1;
  wire [0:0] arrdiv32_fs902_or0;
  wire [0:0] arrdiv32_fs903_xor1;
  wire [0:0] arrdiv32_fs903_or0;
  wire [0:0] arrdiv32_fs904_xor1;
  wire [0:0] arrdiv32_fs904_or0;
  wire [0:0] arrdiv32_fs905_xor1;
  wire [0:0] arrdiv32_fs905_or0;
  wire [0:0] arrdiv32_fs906_xor1;
  wire [0:0] arrdiv32_fs906_or0;
  wire [0:0] arrdiv32_fs907_xor1;
  wire [0:0] arrdiv32_fs907_or0;
  wire [0:0] arrdiv32_fs908_xor1;
  wire [0:0] arrdiv32_fs908_or0;
  wire [0:0] arrdiv32_fs909_xor1;
  wire [0:0] arrdiv32_fs909_or0;
  wire [0:0] arrdiv32_fs910_xor1;
  wire [0:0] arrdiv32_fs910_or0;
  wire [0:0] arrdiv32_fs911_xor1;
  wire [0:0] arrdiv32_fs911_or0;
  wire [0:0] arrdiv32_fs912_xor1;
  wire [0:0] arrdiv32_fs912_or0;
  wire [0:0] arrdiv32_fs913_xor1;
  wire [0:0] arrdiv32_fs913_or0;
  wire [0:0] arrdiv32_fs914_xor1;
  wire [0:0] arrdiv32_fs914_or0;
  wire [0:0] arrdiv32_fs915_xor1;
  wire [0:0] arrdiv32_fs915_or0;
  wire [0:0] arrdiv32_fs916_xor1;
  wire [0:0] arrdiv32_fs916_or0;
  wire [0:0] arrdiv32_fs917_xor1;
  wire [0:0] arrdiv32_fs917_or0;
  wire [0:0] arrdiv32_fs918_xor1;
  wire [0:0] arrdiv32_fs918_or0;
  wire [0:0] arrdiv32_fs919_xor1;
  wire [0:0] arrdiv32_fs919_or0;
  wire [0:0] arrdiv32_fs920_xor1;
  wire [0:0] arrdiv32_fs920_or0;
  wire [0:0] arrdiv32_fs921_xor1;
  wire [0:0] arrdiv32_fs921_or0;
  wire [0:0] arrdiv32_fs922_xor1;
  wire [0:0] arrdiv32_fs922_or0;
  wire [0:0] arrdiv32_fs923_xor1;
  wire [0:0] arrdiv32_fs923_or0;
  wire [0:0] arrdiv32_fs924_xor1;
  wire [0:0] arrdiv32_fs924_or0;
  wire [0:0] arrdiv32_fs925_xor1;
  wire [0:0] arrdiv32_fs925_or0;
  wire [0:0] arrdiv32_fs926_xor1;
  wire [0:0] arrdiv32_fs926_or0;
  wire [0:0] arrdiv32_fs927_xor1;
  wire [0:0] arrdiv32_fs927_or0;
  wire [0:0] arrdiv32_mux2to1868_xor0;
  wire [0:0] arrdiv32_mux2to1869_xor0;
  wire [0:0] arrdiv32_mux2to1870_xor0;
  wire [0:0] arrdiv32_mux2to1871_xor0;
  wire [0:0] arrdiv32_mux2to1872_xor0;
  wire [0:0] arrdiv32_mux2to1873_xor0;
  wire [0:0] arrdiv32_mux2to1874_xor0;
  wire [0:0] arrdiv32_mux2to1875_xor0;
  wire [0:0] arrdiv32_mux2to1876_xor0;
  wire [0:0] arrdiv32_mux2to1877_xor0;
  wire [0:0] arrdiv32_mux2to1878_xor0;
  wire [0:0] arrdiv32_mux2to1879_xor0;
  wire [0:0] arrdiv32_mux2to1880_xor0;
  wire [0:0] arrdiv32_mux2to1881_xor0;
  wire [0:0] arrdiv32_mux2to1882_xor0;
  wire [0:0] arrdiv32_mux2to1883_xor0;
  wire [0:0] arrdiv32_mux2to1884_xor0;
  wire [0:0] arrdiv32_mux2to1885_xor0;
  wire [0:0] arrdiv32_mux2to1886_xor0;
  wire [0:0] arrdiv32_mux2to1887_xor0;
  wire [0:0] arrdiv32_mux2to1888_xor0;
  wire [0:0] arrdiv32_mux2to1889_xor0;
  wire [0:0] arrdiv32_mux2to1890_xor0;
  wire [0:0] arrdiv32_mux2to1891_xor0;
  wire [0:0] arrdiv32_mux2to1892_xor0;
  wire [0:0] arrdiv32_mux2to1893_xor0;
  wire [0:0] arrdiv32_mux2to1894_xor0;
  wire [0:0] arrdiv32_mux2to1895_xor0;
  wire [0:0] arrdiv32_mux2to1896_xor0;
  wire [0:0] arrdiv32_mux2to1897_xor0;
  wire [0:0] arrdiv32_mux2to1898_xor0;
  wire [0:0] arrdiv32_not28;
  wire [0:0] arrdiv32_fs928_xor0;
  wire [0:0] arrdiv32_fs928_and0;
  wire [0:0] arrdiv32_fs929_xor1;
  wire [0:0] arrdiv32_fs929_or0;
  wire [0:0] arrdiv32_fs930_xor1;
  wire [0:0] arrdiv32_fs930_or0;
  wire [0:0] arrdiv32_fs931_xor1;
  wire [0:0] arrdiv32_fs931_or0;
  wire [0:0] arrdiv32_fs932_xor1;
  wire [0:0] arrdiv32_fs932_or0;
  wire [0:0] arrdiv32_fs933_xor1;
  wire [0:0] arrdiv32_fs933_or0;
  wire [0:0] arrdiv32_fs934_xor1;
  wire [0:0] arrdiv32_fs934_or0;
  wire [0:0] arrdiv32_fs935_xor1;
  wire [0:0] arrdiv32_fs935_or0;
  wire [0:0] arrdiv32_fs936_xor1;
  wire [0:0] arrdiv32_fs936_or0;
  wire [0:0] arrdiv32_fs937_xor1;
  wire [0:0] arrdiv32_fs937_or0;
  wire [0:0] arrdiv32_fs938_xor1;
  wire [0:0] arrdiv32_fs938_or0;
  wire [0:0] arrdiv32_fs939_xor1;
  wire [0:0] arrdiv32_fs939_or0;
  wire [0:0] arrdiv32_fs940_xor1;
  wire [0:0] arrdiv32_fs940_or0;
  wire [0:0] arrdiv32_fs941_xor1;
  wire [0:0] arrdiv32_fs941_or0;
  wire [0:0] arrdiv32_fs942_xor1;
  wire [0:0] arrdiv32_fs942_or0;
  wire [0:0] arrdiv32_fs943_xor1;
  wire [0:0] arrdiv32_fs943_or0;
  wire [0:0] arrdiv32_fs944_xor1;
  wire [0:0] arrdiv32_fs944_or0;
  wire [0:0] arrdiv32_fs945_xor1;
  wire [0:0] arrdiv32_fs945_or0;
  wire [0:0] arrdiv32_fs946_xor1;
  wire [0:0] arrdiv32_fs946_or0;
  wire [0:0] arrdiv32_fs947_xor1;
  wire [0:0] arrdiv32_fs947_or0;
  wire [0:0] arrdiv32_fs948_xor1;
  wire [0:0] arrdiv32_fs948_or0;
  wire [0:0] arrdiv32_fs949_xor1;
  wire [0:0] arrdiv32_fs949_or0;
  wire [0:0] arrdiv32_fs950_xor1;
  wire [0:0] arrdiv32_fs950_or0;
  wire [0:0] arrdiv32_fs951_xor1;
  wire [0:0] arrdiv32_fs951_or0;
  wire [0:0] arrdiv32_fs952_xor1;
  wire [0:0] arrdiv32_fs952_or0;
  wire [0:0] arrdiv32_fs953_xor1;
  wire [0:0] arrdiv32_fs953_or0;
  wire [0:0] arrdiv32_fs954_xor1;
  wire [0:0] arrdiv32_fs954_or0;
  wire [0:0] arrdiv32_fs955_xor1;
  wire [0:0] arrdiv32_fs955_or0;
  wire [0:0] arrdiv32_fs956_xor1;
  wire [0:0] arrdiv32_fs956_or0;
  wire [0:0] arrdiv32_fs957_xor1;
  wire [0:0] arrdiv32_fs957_or0;
  wire [0:0] arrdiv32_fs958_xor1;
  wire [0:0] arrdiv32_fs958_or0;
  wire [0:0] arrdiv32_fs959_xor1;
  wire [0:0] arrdiv32_fs959_or0;
  wire [0:0] arrdiv32_mux2to1899_xor0;
  wire [0:0] arrdiv32_mux2to1900_xor0;
  wire [0:0] arrdiv32_mux2to1901_xor0;
  wire [0:0] arrdiv32_mux2to1902_xor0;
  wire [0:0] arrdiv32_mux2to1903_xor0;
  wire [0:0] arrdiv32_mux2to1904_xor0;
  wire [0:0] arrdiv32_mux2to1905_xor0;
  wire [0:0] arrdiv32_mux2to1906_xor0;
  wire [0:0] arrdiv32_mux2to1907_xor0;
  wire [0:0] arrdiv32_mux2to1908_xor0;
  wire [0:0] arrdiv32_mux2to1909_xor0;
  wire [0:0] arrdiv32_mux2to1910_xor0;
  wire [0:0] arrdiv32_mux2to1911_xor0;
  wire [0:0] arrdiv32_mux2to1912_xor0;
  wire [0:0] arrdiv32_mux2to1913_xor0;
  wire [0:0] arrdiv32_mux2to1914_xor0;
  wire [0:0] arrdiv32_mux2to1915_xor0;
  wire [0:0] arrdiv32_mux2to1916_xor0;
  wire [0:0] arrdiv32_mux2to1917_xor0;
  wire [0:0] arrdiv32_mux2to1918_xor0;
  wire [0:0] arrdiv32_mux2to1919_xor0;
  wire [0:0] arrdiv32_mux2to1920_xor0;
  wire [0:0] arrdiv32_mux2to1921_xor0;
  wire [0:0] arrdiv32_mux2to1922_xor0;
  wire [0:0] arrdiv32_mux2to1923_xor0;
  wire [0:0] arrdiv32_mux2to1924_xor0;
  wire [0:0] arrdiv32_mux2to1925_xor0;
  wire [0:0] arrdiv32_mux2to1926_xor0;
  wire [0:0] arrdiv32_mux2to1927_xor0;
  wire [0:0] arrdiv32_mux2to1928_xor0;
  wire [0:0] arrdiv32_mux2to1929_xor0;
  wire [0:0] arrdiv32_not29;
  wire [0:0] arrdiv32_fs960_xor0;
  wire [0:0] arrdiv32_fs960_and0;
  wire [0:0] arrdiv32_fs961_xor1;
  wire [0:0] arrdiv32_fs961_or0;
  wire [0:0] arrdiv32_fs962_xor1;
  wire [0:0] arrdiv32_fs962_or0;
  wire [0:0] arrdiv32_fs963_xor1;
  wire [0:0] arrdiv32_fs963_or0;
  wire [0:0] arrdiv32_fs964_xor1;
  wire [0:0] arrdiv32_fs964_or0;
  wire [0:0] arrdiv32_fs965_xor1;
  wire [0:0] arrdiv32_fs965_or0;
  wire [0:0] arrdiv32_fs966_xor1;
  wire [0:0] arrdiv32_fs966_or0;
  wire [0:0] arrdiv32_fs967_xor1;
  wire [0:0] arrdiv32_fs967_or0;
  wire [0:0] arrdiv32_fs968_xor1;
  wire [0:0] arrdiv32_fs968_or0;
  wire [0:0] arrdiv32_fs969_xor1;
  wire [0:0] arrdiv32_fs969_or0;
  wire [0:0] arrdiv32_fs970_xor1;
  wire [0:0] arrdiv32_fs970_or0;
  wire [0:0] arrdiv32_fs971_xor1;
  wire [0:0] arrdiv32_fs971_or0;
  wire [0:0] arrdiv32_fs972_xor1;
  wire [0:0] arrdiv32_fs972_or0;
  wire [0:0] arrdiv32_fs973_xor1;
  wire [0:0] arrdiv32_fs973_or0;
  wire [0:0] arrdiv32_fs974_xor1;
  wire [0:0] arrdiv32_fs974_or0;
  wire [0:0] arrdiv32_fs975_xor1;
  wire [0:0] arrdiv32_fs975_or0;
  wire [0:0] arrdiv32_fs976_xor1;
  wire [0:0] arrdiv32_fs976_or0;
  wire [0:0] arrdiv32_fs977_xor1;
  wire [0:0] arrdiv32_fs977_or0;
  wire [0:0] arrdiv32_fs978_xor1;
  wire [0:0] arrdiv32_fs978_or0;
  wire [0:0] arrdiv32_fs979_xor1;
  wire [0:0] arrdiv32_fs979_or0;
  wire [0:0] arrdiv32_fs980_xor1;
  wire [0:0] arrdiv32_fs980_or0;
  wire [0:0] arrdiv32_fs981_xor1;
  wire [0:0] arrdiv32_fs981_or0;
  wire [0:0] arrdiv32_fs982_xor1;
  wire [0:0] arrdiv32_fs982_or0;
  wire [0:0] arrdiv32_fs983_xor1;
  wire [0:0] arrdiv32_fs983_or0;
  wire [0:0] arrdiv32_fs984_xor1;
  wire [0:0] arrdiv32_fs984_or0;
  wire [0:0] arrdiv32_fs985_xor1;
  wire [0:0] arrdiv32_fs985_or0;
  wire [0:0] arrdiv32_fs986_xor1;
  wire [0:0] arrdiv32_fs986_or0;
  wire [0:0] arrdiv32_fs987_xor1;
  wire [0:0] arrdiv32_fs987_or0;
  wire [0:0] arrdiv32_fs988_xor1;
  wire [0:0] arrdiv32_fs988_or0;
  wire [0:0] arrdiv32_fs989_xor1;
  wire [0:0] arrdiv32_fs989_or0;
  wire [0:0] arrdiv32_fs990_xor1;
  wire [0:0] arrdiv32_fs990_or0;
  wire [0:0] arrdiv32_fs991_xor1;
  wire [0:0] arrdiv32_fs991_or0;
  wire [0:0] arrdiv32_mux2to1930_xor0;
  wire [0:0] arrdiv32_mux2to1931_xor0;
  wire [0:0] arrdiv32_mux2to1932_xor0;
  wire [0:0] arrdiv32_mux2to1933_xor0;
  wire [0:0] arrdiv32_mux2to1934_xor0;
  wire [0:0] arrdiv32_mux2to1935_xor0;
  wire [0:0] arrdiv32_mux2to1936_xor0;
  wire [0:0] arrdiv32_mux2to1937_xor0;
  wire [0:0] arrdiv32_mux2to1938_xor0;
  wire [0:0] arrdiv32_mux2to1939_xor0;
  wire [0:0] arrdiv32_mux2to1940_xor0;
  wire [0:0] arrdiv32_mux2to1941_xor0;
  wire [0:0] arrdiv32_mux2to1942_xor0;
  wire [0:0] arrdiv32_mux2to1943_xor0;
  wire [0:0] arrdiv32_mux2to1944_xor0;
  wire [0:0] arrdiv32_mux2to1945_xor0;
  wire [0:0] arrdiv32_mux2to1946_xor0;
  wire [0:0] arrdiv32_mux2to1947_xor0;
  wire [0:0] arrdiv32_mux2to1948_xor0;
  wire [0:0] arrdiv32_mux2to1949_xor0;
  wire [0:0] arrdiv32_mux2to1950_xor0;
  wire [0:0] arrdiv32_mux2to1951_xor0;
  wire [0:0] arrdiv32_mux2to1952_xor0;
  wire [0:0] arrdiv32_mux2to1953_xor0;
  wire [0:0] arrdiv32_mux2to1954_xor0;
  wire [0:0] arrdiv32_mux2to1955_xor0;
  wire [0:0] arrdiv32_mux2to1956_xor0;
  wire [0:0] arrdiv32_mux2to1957_xor0;
  wire [0:0] arrdiv32_mux2to1958_xor0;
  wire [0:0] arrdiv32_mux2to1959_xor0;
  wire [0:0] arrdiv32_mux2to1960_xor0;
  wire [0:0] arrdiv32_not30;
  wire [0:0] arrdiv32_fs992_xor0;
  wire [0:0] arrdiv32_fs992_and0;
  wire [0:0] arrdiv32_fs993_xor1;
  wire [0:0] arrdiv32_fs993_or0;
  wire [0:0] arrdiv32_fs994_xor1;
  wire [0:0] arrdiv32_fs994_or0;
  wire [0:0] arrdiv32_fs995_xor1;
  wire [0:0] arrdiv32_fs995_or0;
  wire [0:0] arrdiv32_fs996_xor1;
  wire [0:0] arrdiv32_fs996_or0;
  wire [0:0] arrdiv32_fs997_xor1;
  wire [0:0] arrdiv32_fs997_or0;
  wire [0:0] arrdiv32_fs998_xor1;
  wire [0:0] arrdiv32_fs998_or0;
  wire [0:0] arrdiv32_fs999_xor1;
  wire [0:0] arrdiv32_fs999_or0;
  wire [0:0] arrdiv32_fs1000_xor1;
  wire [0:0] arrdiv32_fs1000_or0;
  wire [0:0] arrdiv32_fs1001_xor1;
  wire [0:0] arrdiv32_fs1001_or0;
  wire [0:0] arrdiv32_fs1002_xor1;
  wire [0:0] arrdiv32_fs1002_or0;
  wire [0:0] arrdiv32_fs1003_xor1;
  wire [0:0] arrdiv32_fs1003_or0;
  wire [0:0] arrdiv32_fs1004_xor1;
  wire [0:0] arrdiv32_fs1004_or0;
  wire [0:0] arrdiv32_fs1005_xor1;
  wire [0:0] arrdiv32_fs1005_or0;
  wire [0:0] arrdiv32_fs1006_xor1;
  wire [0:0] arrdiv32_fs1006_or0;
  wire [0:0] arrdiv32_fs1007_xor1;
  wire [0:0] arrdiv32_fs1007_or0;
  wire [0:0] arrdiv32_fs1008_xor1;
  wire [0:0] arrdiv32_fs1008_or0;
  wire [0:0] arrdiv32_fs1009_xor1;
  wire [0:0] arrdiv32_fs1009_or0;
  wire [0:0] arrdiv32_fs1010_xor1;
  wire [0:0] arrdiv32_fs1010_or0;
  wire [0:0] arrdiv32_fs1011_xor1;
  wire [0:0] arrdiv32_fs1011_or0;
  wire [0:0] arrdiv32_fs1012_xor1;
  wire [0:0] arrdiv32_fs1012_or0;
  wire [0:0] arrdiv32_fs1013_xor1;
  wire [0:0] arrdiv32_fs1013_or0;
  wire [0:0] arrdiv32_fs1014_xor1;
  wire [0:0] arrdiv32_fs1014_or0;
  wire [0:0] arrdiv32_fs1015_xor1;
  wire [0:0] arrdiv32_fs1015_or0;
  wire [0:0] arrdiv32_fs1016_xor1;
  wire [0:0] arrdiv32_fs1016_or0;
  wire [0:0] arrdiv32_fs1017_xor1;
  wire [0:0] arrdiv32_fs1017_or0;
  wire [0:0] arrdiv32_fs1018_xor1;
  wire [0:0] arrdiv32_fs1018_or0;
  wire [0:0] arrdiv32_fs1019_xor1;
  wire [0:0] arrdiv32_fs1019_or0;
  wire [0:0] arrdiv32_fs1020_xor1;
  wire [0:0] arrdiv32_fs1020_or0;
  wire [0:0] arrdiv32_fs1021_xor1;
  wire [0:0] arrdiv32_fs1021_or0;
  wire [0:0] arrdiv32_fs1022_xor1;
  wire [0:0] arrdiv32_fs1022_or0;
  wire [0:0] arrdiv32_fs1023_xor1;
  wire [0:0] arrdiv32_fs1023_or0;
  wire [0:0] arrdiv32_not31;

  fs fs_arrdiv32_fs0_out(.a(a[31]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs0_xor0), .fs_or0(arrdiv32_fs0_and0));
  fs fs_arrdiv32_fs1_out(.a(1'b0), .b(b[1]), .bin(arrdiv32_fs0_and0[0]), .fs_xor1(arrdiv32_fs1_xor1), .fs_or0(arrdiv32_fs1_or0));
  fs fs_arrdiv32_fs2_out(.a(1'b0), .b(b[2]), .bin(arrdiv32_fs1_or0[0]), .fs_xor1(arrdiv32_fs2_xor1), .fs_or0(arrdiv32_fs2_or0));
  fs fs_arrdiv32_fs3_out(.a(1'b0), .b(b[3]), .bin(arrdiv32_fs2_or0[0]), .fs_xor1(arrdiv32_fs3_xor1), .fs_or0(arrdiv32_fs3_or0));
  fs fs_arrdiv32_fs4_out(.a(1'b0), .b(b[4]), .bin(arrdiv32_fs3_or0[0]), .fs_xor1(arrdiv32_fs4_xor1), .fs_or0(arrdiv32_fs4_or0));
  fs fs_arrdiv32_fs5_out(.a(1'b0), .b(b[5]), .bin(arrdiv32_fs4_or0[0]), .fs_xor1(arrdiv32_fs5_xor1), .fs_or0(arrdiv32_fs5_or0));
  fs fs_arrdiv32_fs6_out(.a(1'b0), .b(b[6]), .bin(arrdiv32_fs5_or0[0]), .fs_xor1(arrdiv32_fs6_xor1), .fs_or0(arrdiv32_fs6_or0));
  fs fs_arrdiv32_fs7_out(.a(1'b0), .b(b[7]), .bin(arrdiv32_fs6_or0[0]), .fs_xor1(arrdiv32_fs7_xor1), .fs_or0(arrdiv32_fs7_or0));
  fs fs_arrdiv32_fs8_out(.a(1'b0), .b(b[8]), .bin(arrdiv32_fs7_or0[0]), .fs_xor1(arrdiv32_fs8_xor1), .fs_or0(arrdiv32_fs8_or0));
  fs fs_arrdiv32_fs9_out(.a(1'b0), .b(b[9]), .bin(arrdiv32_fs8_or0[0]), .fs_xor1(arrdiv32_fs9_xor1), .fs_or0(arrdiv32_fs9_or0));
  fs fs_arrdiv32_fs10_out(.a(1'b0), .b(b[10]), .bin(arrdiv32_fs9_or0[0]), .fs_xor1(arrdiv32_fs10_xor1), .fs_or0(arrdiv32_fs10_or0));
  fs fs_arrdiv32_fs11_out(.a(1'b0), .b(b[11]), .bin(arrdiv32_fs10_or0[0]), .fs_xor1(arrdiv32_fs11_xor1), .fs_or0(arrdiv32_fs11_or0));
  fs fs_arrdiv32_fs12_out(.a(1'b0), .b(b[12]), .bin(arrdiv32_fs11_or0[0]), .fs_xor1(arrdiv32_fs12_xor1), .fs_or0(arrdiv32_fs12_or0));
  fs fs_arrdiv32_fs13_out(.a(1'b0), .b(b[13]), .bin(arrdiv32_fs12_or0[0]), .fs_xor1(arrdiv32_fs13_xor1), .fs_or0(arrdiv32_fs13_or0));
  fs fs_arrdiv32_fs14_out(.a(1'b0), .b(b[14]), .bin(arrdiv32_fs13_or0[0]), .fs_xor1(arrdiv32_fs14_xor1), .fs_or0(arrdiv32_fs14_or0));
  fs fs_arrdiv32_fs15_out(.a(1'b0), .b(b[15]), .bin(arrdiv32_fs14_or0[0]), .fs_xor1(arrdiv32_fs15_xor1), .fs_or0(arrdiv32_fs15_or0));
  fs fs_arrdiv32_fs16_out(.a(1'b0), .b(b[16]), .bin(arrdiv32_fs15_or0[0]), .fs_xor1(arrdiv32_fs16_xor1), .fs_or0(arrdiv32_fs16_or0));
  fs fs_arrdiv32_fs17_out(.a(1'b0), .b(b[17]), .bin(arrdiv32_fs16_or0[0]), .fs_xor1(arrdiv32_fs17_xor1), .fs_or0(arrdiv32_fs17_or0));
  fs fs_arrdiv32_fs18_out(.a(1'b0), .b(b[18]), .bin(arrdiv32_fs17_or0[0]), .fs_xor1(arrdiv32_fs18_xor1), .fs_or0(arrdiv32_fs18_or0));
  fs fs_arrdiv32_fs19_out(.a(1'b0), .b(b[19]), .bin(arrdiv32_fs18_or0[0]), .fs_xor1(arrdiv32_fs19_xor1), .fs_or0(arrdiv32_fs19_or0));
  fs fs_arrdiv32_fs20_out(.a(1'b0), .b(b[20]), .bin(arrdiv32_fs19_or0[0]), .fs_xor1(arrdiv32_fs20_xor1), .fs_or0(arrdiv32_fs20_or0));
  fs fs_arrdiv32_fs21_out(.a(1'b0), .b(b[21]), .bin(arrdiv32_fs20_or0[0]), .fs_xor1(arrdiv32_fs21_xor1), .fs_or0(arrdiv32_fs21_or0));
  fs fs_arrdiv32_fs22_out(.a(1'b0), .b(b[22]), .bin(arrdiv32_fs21_or0[0]), .fs_xor1(arrdiv32_fs22_xor1), .fs_or0(arrdiv32_fs22_or0));
  fs fs_arrdiv32_fs23_out(.a(1'b0), .b(b[23]), .bin(arrdiv32_fs22_or0[0]), .fs_xor1(arrdiv32_fs23_xor1), .fs_or0(arrdiv32_fs23_or0));
  fs fs_arrdiv32_fs24_out(.a(1'b0), .b(b[24]), .bin(arrdiv32_fs23_or0[0]), .fs_xor1(arrdiv32_fs24_xor1), .fs_or0(arrdiv32_fs24_or0));
  fs fs_arrdiv32_fs25_out(.a(1'b0), .b(b[25]), .bin(arrdiv32_fs24_or0[0]), .fs_xor1(arrdiv32_fs25_xor1), .fs_or0(arrdiv32_fs25_or0));
  fs fs_arrdiv32_fs26_out(.a(1'b0), .b(b[26]), .bin(arrdiv32_fs25_or0[0]), .fs_xor1(arrdiv32_fs26_xor1), .fs_or0(arrdiv32_fs26_or0));
  fs fs_arrdiv32_fs27_out(.a(1'b0), .b(b[27]), .bin(arrdiv32_fs26_or0[0]), .fs_xor1(arrdiv32_fs27_xor1), .fs_or0(arrdiv32_fs27_or0));
  fs fs_arrdiv32_fs28_out(.a(1'b0), .b(b[28]), .bin(arrdiv32_fs27_or0[0]), .fs_xor1(arrdiv32_fs28_xor1), .fs_or0(arrdiv32_fs28_or0));
  fs fs_arrdiv32_fs29_out(.a(1'b0), .b(b[29]), .bin(arrdiv32_fs28_or0[0]), .fs_xor1(arrdiv32_fs29_xor1), .fs_or0(arrdiv32_fs29_or0));
  fs fs_arrdiv32_fs30_out(.a(1'b0), .b(b[30]), .bin(arrdiv32_fs29_or0[0]), .fs_xor1(arrdiv32_fs30_xor1), .fs_or0(arrdiv32_fs30_or0));
  fs fs_arrdiv32_fs31_out(.a(1'b0), .b(b[31]), .bin(arrdiv32_fs30_or0[0]), .fs_xor1(arrdiv32_fs31_xor1), .fs_or0(arrdiv32_fs31_or0));
  mux2to1 mux2to1_arrdiv32_mux2to10_out(.d0(arrdiv32_fs0_xor0[0]), .d1(a[31]), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to10_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to11_out(.d0(arrdiv32_fs1_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to11_and1));
  mux2to1 mux2to1_arrdiv32_mux2to12_out(.d0(arrdiv32_fs2_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to12_and1));
  mux2to1 mux2to1_arrdiv32_mux2to13_out(.d0(arrdiv32_fs3_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to13_and1));
  mux2to1 mux2to1_arrdiv32_mux2to14_out(.d0(arrdiv32_fs4_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to14_and1));
  mux2to1 mux2to1_arrdiv32_mux2to15_out(.d0(arrdiv32_fs5_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to15_and1));
  mux2to1 mux2to1_arrdiv32_mux2to16_out(.d0(arrdiv32_fs6_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to16_and1));
  mux2to1 mux2to1_arrdiv32_mux2to17_out(.d0(arrdiv32_fs7_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to17_and1));
  mux2to1 mux2to1_arrdiv32_mux2to18_out(.d0(arrdiv32_fs8_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to18_and1));
  mux2to1 mux2to1_arrdiv32_mux2to19_out(.d0(arrdiv32_fs9_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to19_and1));
  mux2to1 mux2to1_arrdiv32_mux2to110_out(.d0(arrdiv32_fs10_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to110_and1));
  mux2to1 mux2to1_arrdiv32_mux2to111_out(.d0(arrdiv32_fs11_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to111_and1));
  mux2to1 mux2to1_arrdiv32_mux2to112_out(.d0(arrdiv32_fs12_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to112_and1));
  mux2to1 mux2to1_arrdiv32_mux2to113_out(.d0(arrdiv32_fs13_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to113_and1));
  mux2to1 mux2to1_arrdiv32_mux2to114_out(.d0(arrdiv32_fs14_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to114_and1));
  mux2to1 mux2to1_arrdiv32_mux2to115_out(.d0(arrdiv32_fs15_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to115_and1));
  mux2to1 mux2to1_arrdiv32_mux2to116_out(.d0(arrdiv32_fs16_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to116_and1));
  mux2to1 mux2to1_arrdiv32_mux2to117_out(.d0(arrdiv32_fs17_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to117_and1));
  mux2to1 mux2to1_arrdiv32_mux2to118_out(.d0(arrdiv32_fs18_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to118_and1));
  mux2to1 mux2to1_arrdiv32_mux2to119_out(.d0(arrdiv32_fs19_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to119_and1));
  mux2to1 mux2to1_arrdiv32_mux2to120_out(.d0(arrdiv32_fs20_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to120_and1));
  mux2to1 mux2to1_arrdiv32_mux2to121_out(.d0(arrdiv32_fs21_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to121_and1));
  mux2to1 mux2to1_arrdiv32_mux2to122_out(.d0(arrdiv32_fs22_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to122_and1));
  mux2to1 mux2to1_arrdiv32_mux2to123_out(.d0(arrdiv32_fs23_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to123_and1));
  mux2to1 mux2to1_arrdiv32_mux2to124_out(.d0(arrdiv32_fs24_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to124_and1));
  mux2to1 mux2to1_arrdiv32_mux2to125_out(.d0(arrdiv32_fs25_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to125_and1));
  mux2to1 mux2to1_arrdiv32_mux2to126_out(.d0(arrdiv32_fs26_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to126_and1));
  mux2to1 mux2to1_arrdiv32_mux2to127_out(.d0(arrdiv32_fs27_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to127_and1));
  mux2to1 mux2to1_arrdiv32_mux2to128_out(.d0(arrdiv32_fs28_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to128_and1));
  mux2to1 mux2to1_arrdiv32_mux2to129_out(.d0(arrdiv32_fs29_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to129_and1));
  mux2to1 mux2to1_arrdiv32_mux2to130_out(.d0(arrdiv32_fs30_xor1[0]), .d1(1'b0), .sel(arrdiv32_fs31_or0[0]), .mux2to1_xor0(arrdiv32_mux2to130_and1));
  not_gate not_gate_arrdiv32_not0(.a(arrdiv32_fs31_or0[0]), .out(arrdiv32_not0));
  fs fs_arrdiv32_fs32_out(.a(a[30]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs32_xor0), .fs_or0(arrdiv32_fs32_and0));
  fs fs_arrdiv32_fs33_out(.a(arrdiv32_mux2to10_xor0[0]), .b(b[1]), .bin(arrdiv32_fs32_and0[0]), .fs_xor1(arrdiv32_fs33_xor1), .fs_or0(arrdiv32_fs33_or0));
  fs fs_arrdiv32_fs34_out(.a(arrdiv32_mux2to11_and1[0]), .b(b[2]), .bin(arrdiv32_fs33_or0[0]), .fs_xor1(arrdiv32_fs34_xor1), .fs_or0(arrdiv32_fs34_or0));
  fs fs_arrdiv32_fs35_out(.a(arrdiv32_mux2to12_and1[0]), .b(b[3]), .bin(arrdiv32_fs34_or0[0]), .fs_xor1(arrdiv32_fs35_xor1), .fs_or0(arrdiv32_fs35_or0));
  fs fs_arrdiv32_fs36_out(.a(arrdiv32_mux2to13_and1[0]), .b(b[4]), .bin(arrdiv32_fs35_or0[0]), .fs_xor1(arrdiv32_fs36_xor1), .fs_or0(arrdiv32_fs36_or0));
  fs fs_arrdiv32_fs37_out(.a(arrdiv32_mux2to14_and1[0]), .b(b[5]), .bin(arrdiv32_fs36_or0[0]), .fs_xor1(arrdiv32_fs37_xor1), .fs_or0(arrdiv32_fs37_or0));
  fs fs_arrdiv32_fs38_out(.a(arrdiv32_mux2to15_and1[0]), .b(b[6]), .bin(arrdiv32_fs37_or0[0]), .fs_xor1(arrdiv32_fs38_xor1), .fs_or0(arrdiv32_fs38_or0));
  fs fs_arrdiv32_fs39_out(.a(arrdiv32_mux2to16_and1[0]), .b(b[7]), .bin(arrdiv32_fs38_or0[0]), .fs_xor1(arrdiv32_fs39_xor1), .fs_or0(arrdiv32_fs39_or0));
  fs fs_arrdiv32_fs40_out(.a(arrdiv32_mux2to17_and1[0]), .b(b[8]), .bin(arrdiv32_fs39_or0[0]), .fs_xor1(arrdiv32_fs40_xor1), .fs_or0(arrdiv32_fs40_or0));
  fs fs_arrdiv32_fs41_out(.a(arrdiv32_mux2to18_and1[0]), .b(b[9]), .bin(arrdiv32_fs40_or0[0]), .fs_xor1(arrdiv32_fs41_xor1), .fs_or0(arrdiv32_fs41_or0));
  fs fs_arrdiv32_fs42_out(.a(arrdiv32_mux2to19_and1[0]), .b(b[10]), .bin(arrdiv32_fs41_or0[0]), .fs_xor1(arrdiv32_fs42_xor1), .fs_or0(arrdiv32_fs42_or0));
  fs fs_arrdiv32_fs43_out(.a(arrdiv32_mux2to110_and1[0]), .b(b[11]), .bin(arrdiv32_fs42_or0[0]), .fs_xor1(arrdiv32_fs43_xor1), .fs_or0(arrdiv32_fs43_or0));
  fs fs_arrdiv32_fs44_out(.a(arrdiv32_mux2to111_and1[0]), .b(b[12]), .bin(arrdiv32_fs43_or0[0]), .fs_xor1(arrdiv32_fs44_xor1), .fs_or0(arrdiv32_fs44_or0));
  fs fs_arrdiv32_fs45_out(.a(arrdiv32_mux2to112_and1[0]), .b(b[13]), .bin(arrdiv32_fs44_or0[0]), .fs_xor1(arrdiv32_fs45_xor1), .fs_or0(arrdiv32_fs45_or0));
  fs fs_arrdiv32_fs46_out(.a(arrdiv32_mux2to113_and1[0]), .b(b[14]), .bin(arrdiv32_fs45_or0[0]), .fs_xor1(arrdiv32_fs46_xor1), .fs_or0(arrdiv32_fs46_or0));
  fs fs_arrdiv32_fs47_out(.a(arrdiv32_mux2to114_and1[0]), .b(b[15]), .bin(arrdiv32_fs46_or0[0]), .fs_xor1(arrdiv32_fs47_xor1), .fs_or0(arrdiv32_fs47_or0));
  fs fs_arrdiv32_fs48_out(.a(arrdiv32_mux2to115_and1[0]), .b(b[16]), .bin(arrdiv32_fs47_or0[0]), .fs_xor1(arrdiv32_fs48_xor1), .fs_or0(arrdiv32_fs48_or0));
  fs fs_arrdiv32_fs49_out(.a(arrdiv32_mux2to116_and1[0]), .b(b[17]), .bin(arrdiv32_fs48_or0[0]), .fs_xor1(arrdiv32_fs49_xor1), .fs_or0(arrdiv32_fs49_or0));
  fs fs_arrdiv32_fs50_out(.a(arrdiv32_mux2to117_and1[0]), .b(b[18]), .bin(arrdiv32_fs49_or0[0]), .fs_xor1(arrdiv32_fs50_xor1), .fs_or0(arrdiv32_fs50_or0));
  fs fs_arrdiv32_fs51_out(.a(arrdiv32_mux2to118_and1[0]), .b(b[19]), .bin(arrdiv32_fs50_or0[0]), .fs_xor1(arrdiv32_fs51_xor1), .fs_or0(arrdiv32_fs51_or0));
  fs fs_arrdiv32_fs52_out(.a(arrdiv32_mux2to119_and1[0]), .b(b[20]), .bin(arrdiv32_fs51_or0[0]), .fs_xor1(arrdiv32_fs52_xor1), .fs_or0(arrdiv32_fs52_or0));
  fs fs_arrdiv32_fs53_out(.a(arrdiv32_mux2to120_and1[0]), .b(b[21]), .bin(arrdiv32_fs52_or0[0]), .fs_xor1(arrdiv32_fs53_xor1), .fs_or0(arrdiv32_fs53_or0));
  fs fs_arrdiv32_fs54_out(.a(arrdiv32_mux2to121_and1[0]), .b(b[22]), .bin(arrdiv32_fs53_or0[0]), .fs_xor1(arrdiv32_fs54_xor1), .fs_or0(arrdiv32_fs54_or0));
  fs fs_arrdiv32_fs55_out(.a(arrdiv32_mux2to122_and1[0]), .b(b[23]), .bin(arrdiv32_fs54_or0[0]), .fs_xor1(arrdiv32_fs55_xor1), .fs_or0(arrdiv32_fs55_or0));
  fs fs_arrdiv32_fs56_out(.a(arrdiv32_mux2to123_and1[0]), .b(b[24]), .bin(arrdiv32_fs55_or0[0]), .fs_xor1(arrdiv32_fs56_xor1), .fs_or0(arrdiv32_fs56_or0));
  fs fs_arrdiv32_fs57_out(.a(arrdiv32_mux2to124_and1[0]), .b(b[25]), .bin(arrdiv32_fs56_or0[0]), .fs_xor1(arrdiv32_fs57_xor1), .fs_or0(arrdiv32_fs57_or0));
  fs fs_arrdiv32_fs58_out(.a(arrdiv32_mux2to125_and1[0]), .b(b[26]), .bin(arrdiv32_fs57_or0[0]), .fs_xor1(arrdiv32_fs58_xor1), .fs_or0(arrdiv32_fs58_or0));
  fs fs_arrdiv32_fs59_out(.a(arrdiv32_mux2to126_and1[0]), .b(b[27]), .bin(arrdiv32_fs58_or0[0]), .fs_xor1(arrdiv32_fs59_xor1), .fs_or0(arrdiv32_fs59_or0));
  fs fs_arrdiv32_fs60_out(.a(arrdiv32_mux2to127_and1[0]), .b(b[28]), .bin(arrdiv32_fs59_or0[0]), .fs_xor1(arrdiv32_fs60_xor1), .fs_or0(arrdiv32_fs60_or0));
  fs fs_arrdiv32_fs61_out(.a(arrdiv32_mux2to128_and1[0]), .b(b[29]), .bin(arrdiv32_fs60_or0[0]), .fs_xor1(arrdiv32_fs61_xor1), .fs_or0(arrdiv32_fs61_or0));
  fs fs_arrdiv32_fs62_out(.a(arrdiv32_mux2to129_and1[0]), .b(b[30]), .bin(arrdiv32_fs61_or0[0]), .fs_xor1(arrdiv32_fs62_xor1), .fs_or0(arrdiv32_fs62_or0));
  fs fs_arrdiv32_fs63_out(.a(arrdiv32_mux2to130_and1[0]), .b(b[31]), .bin(arrdiv32_fs62_or0[0]), .fs_xor1(arrdiv32_fs63_xor1), .fs_or0(arrdiv32_fs63_or0));
  mux2to1 mux2to1_arrdiv32_mux2to131_out(.d0(arrdiv32_fs32_xor0[0]), .d1(a[30]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to131_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to132_out(.d0(arrdiv32_fs33_xor1[0]), .d1(arrdiv32_mux2to10_xor0[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to132_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to133_out(.d0(arrdiv32_fs34_xor1[0]), .d1(arrdiv32_mux2to11_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to133_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to134_out(.d0(arrdiv32_fs35_xor1[0]), .d1(arrdiv32_mux2to12_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to134_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to135_out(.d0(arrdiv32_fs36_xor1[0]), .d1(arrdiv32_mux2to13_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to135_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to136_out(.d0(arrdiv32_fs37_xor1[0]), .d1(arrdiv32_mux2to14_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to136_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to137_out(.d0(arrdiv32_fs38_xor1[0]), .d1(arrdiv32_mux2to15_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to137_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to138_out(.d0(arrdiv32_fs39_xor1[0]), .d1(arrdiv32_mux2to16_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to138_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to139_out(.d0(arrdiv32_fs40_xor1[0]), .d1(arrdiv32_mux2to17_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to139_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to140_out(.d0(arrdiv32_fs41_xor1[0]), .d1(arrdiv32_mux2to18_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to140_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to141_out(.d0(arrdiv32_fs42_xor1[0]), .d1(arrdiv32_mux2to19_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to141_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to142_out(.d0(arrdiv32_fs43_xor1[0]), .d1(arrdiv32_mux2to110_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to142_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to143_out(.d0(arrdiv32_fs44_xor1[0]), .d1(arrdiv32_mux2to111_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to143_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to144_out(.d0(arrdiv32_fs45_xor1[0]), .d1(arrdiv32_mux2to112_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to144_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to145_out(.d0(arrdiv32_fs46_xor1[0]), .d1(arrdiv32_mux2to113_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to145_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to146_out(.d0(arrdiv32_fs47_xor1[0]), .d1(arrdiv32_mux2to114_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to146_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to147_out(.d0(arrdiv32_fs48_xor1[0]), .d1(arrdiv32_mux2to115_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to147_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to148_out(.d0(arrdiv32_fs49_xor1[0]), .d1(arrdiv32_mux2to116_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to148_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to149_out(.d0(arrdiv32_fs50_xor1[0]), .d1(arrdiv32_mux2to117_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to149_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to150_out(.d0(arrdiv32_fs51_xor1[0]), .d1(arrdiv32_mux2to118_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to150_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to151_out(.d0(arrdiv32_fs52_xor1[0]), .d1(arrdiv32_mux2to119_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to151_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to152_out(.d0(arrdiv32_fs53_xor1[0]), .d1(arrdiv32_mux2to120_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to152_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to153_out(.d0(arrdiv32_fs54_xor1[0]), .d1(arrdiv32_mux2to121_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to153_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to154_out(.d0(arrdiv32_fs55_xor1[0]), .d1(arrdiv32_mux2to122_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to154_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to155_out(.d0(arrdiv32_fs56_xor1[0]), .d1(arrdiv32_mux2to123_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to155_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to156_out(.d0(arrdiv32_fs57_xor1[0]), .d1(arrdiv32_mux2to124_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to156_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to157_out(.d0(arrdiv32_fs58_xor1[0]), .d1(arrdiv32_mux2to125_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to157_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to158_out(.d0(arrdiv32_fs59_xor1[0]), .d1(arrdiv32_mux2to126_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to158_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to159_out(.d0(arrdiv32_fs60_xor1[0]), .d1(arrdiv32_mux2to127_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to159_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to160_out(.d0(arrdiv32_fs61_xor1[0]), .d1(arrdiv32_mux2to128_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to160_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to161_out(.d0(arrdiv32_fs62_xor1[0]), .d1(arrdiv32_mux2to129_and1[0]), .sel(arrdiv32_fs63_or0[0]), .mux2to1_xor0(arrdiv32_mux2to161_xor0));
  not_gate not_gate_arrdiv32_not1(.a(arrdiv32_fs63_or0[0]), .out(arrdiv32_not1));
  fs fs_arrdiv32_fs64_out(.a(a[29]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs64_xor0), .fs_or0(arrdiv32_fs64_and0));
  fs fs_arrdiv32_fs65_out(.a(arrdiv32_mux2to131_xor0[0]), .b(b[1]), .bin(arrdiv32_fs64_and0[0]), .fs_xor1(arrdiv32_fs65_xor1), .fs_or0(arrdiv32_fs65_or0));
  fs fs_arrdiv32_fs66_out(.a(arrdiv32_mux2to132_xor0[0]), .b(b[2]), .bin(arrdiv32_fs65_or0[0]), .fs_xor1(arrdiv32_fs66_xor1), .fs_or0(arrdiv32_fs66_or0));
  fs fs_arrdiv32_fs67_out(.a(arrdiv32_mux2to133_xor0[0]), .b(b[3]), .bin(arrdiv32_fs66_or0[0]), .fs_xor1(arrdiv32_fs67_xor1), .fs_or0(arrdiv32_fs67_or0));
  fs fs_arrdiv32_fs68_out(.a(arrdiv32_mux2to134_xor0[0]), .b(b[4]), .bin(arrdiv32_fs67_or0[0]), .fs_xor1(arrdiv32_fs68_xor1), .fs_or0(arrdiv32_fs68_or0));
  fs fs_arrdiv32_fs69_out(.a(arrdiv32_mux2to135_xor0[0]), .b(b[5]), .bin(arrdiv32_fs68_or0[0]), .fs_xor1(arrdiv32_fs69_xor1), .fs_or0(arrdiv32_fs69_or0));
  fs fs_arrdiv32_fs70_out(.a(arrdiv32_mux2to136_xor0[0]), .b(b[6]), .bin(arrdiv32_fs69_or0[0]), .fs_xor1(arrdiv32_fs70_xor1), .fs_or0(arrdiv32_fs70_or0));
  fs fs_arrdiv32_fs71_out(.a(arrdiv32_mux2to137_xor0[0]), .b(b[7]), .bin(arrdiv32_fs70_or0[0]), .fs_xor1(arrdiv32_fs71_xor1), .fs_or0(arrdiv32_fs71_or0));
  fs fs_arrdiv32_fs72_out(.a(arrdiv32_mux2to138_xor0[0]), .b(b[8]), .bin(arrdiv32_fs71_or0[0]), .fs_xor1(arrdiv32_fs72_xor1), .fs_or0(arrdiv32_fs72_or0));
  fs fs_arrdiv32_fs73_out(.a(arrdiv32_mux2to139_xor0[0]), .b(b[9]), .bin(arrdiv32_fs72_or0[0]), .fs_xor1(arrdiv32_fs73_xor1), .fs_or0(arrdiv32_fs73_or0));
  fs fs_arrdiv32_fs74_out(.a(arrdiv32_mux2to140_xor0[0]), .b(b[10]), .bin(arrdiv32_fs73_or0[0]), .fs_xor1(arrdiv32_fs74_xor1), .fs_or0(arrdiv32_fs74_or0));
  fs fs_arrdiv32_fs75_out(.a(arrdiv32_mux2to141_xor0[0]), .b(b[11]), .bin(arrdiv32_fs74_or0[0]), .fs_xor1(arrdiv32_fs75_xor1), .fs_or0(arrdiv32_fs75_or0));
  fs fs_arrdiv32_fs76_out(.a(arrdiv32_mux2to142_xor0[0]), .b(b[12]), .bin(arrdiv32_fs75_or0[0]), .fs_xor1(arrdiv32_fs76_xor1), .fs_or0(arrdiv32_fs76_or0));
  fs fs_arrdiv32_fs77_out(.a(arrdiv32_mux2to143_xor0[0]), .b(b[13]), .bin(arrdiv32_fs76_or0[0]), .fs_xor1(arrdiv32_fs77_xor1), .fs_or0(arrdiv32_fs77_or0));
  fs fs_arrdiv32_fs78_out(.a(arrdiv32_mux2to144_xor0[0]), .b(b[14]), .bin(arrdiv32_fs77_or0[0]), .fs_xor1(arrdiv32_fs78_xor1), .fs_or0(arrdiv32_fs78_or0));
  fs fs_arrdiv32_fs79_out(.a(arrdiv32_mux2to145_xor0[0]), .b(b[15]), .bin(arrdiv32_fs78_or0[0]), .fs_xor1(arrdiv32_fs79_xor1), .fs_or0(arrdiv32_fs79_or0));
  fs fs_arrdiv32_fs80_out(.a(arrdiv32_mux2to146_xor0[0]), .b(b[16]), .bin(arrdiv32_fs79_or0[0]), .fs_xor1(arrdiv32_fs80_xor1), .fs_or0(arrdiv32_fs80_or0));
  fs fs_arrdiv32_fs81_out(.a(arrdiv32_mux2to147_xor0[0]), .b(b[17]), .bin(arrdiv32_fs80_or0[0]), .fs_xor1(arrdiv32_fs81_xor1), .fs_or0(arrdiv32_fs81_or0));
  fs fs_arrdiv32_fs82_out(.a(arrdiv32_mux2to148_xor0[0]), .b(b[18]), .bin(arrdiv32_fs81_or0[0]), .fs_xor1(arrdiv32_fs82_xor1), .fs_or0(arrdiv32_fs82_or0));
  fs fs_arrdiv32_fs83_out(.a(arrdiv32_mux2to149_xor0[0]), .b(b[19]), .bin(arrdiv32_fs82_or0[0]), .fs_xor1(arrdiv32_fs83_xor1), .fs_or0(arrdiv32_fs83_or0));
  fs fs_arrdiv32_fs84_out(.a(arrdiv32_mux2to150_xor0[0]), .b(b[20]), .bin(arrdiv32_fs83_or0[0]), .fs_xor1(arrdiv32_fs84_xor1), .fs_or0(arrdiv32_fs84_or0));
  fs fs_arrdiv32_fs85_out(.a(arrdiv32_mux2to151_xor0[0]), .b(b[21]), .bin(arrdiv32_fs84_or0[0]), .fs_xor1(arrdiv32_fs85_xor1), .fs_or0(arrdiv32_fs85_or0));
  fs fs_arrdiv32_fs86_out(.a(arrdiv32_mux2to152_xor0[0]), .b(b[22]), .bin(arrdiv32_fs85_or0[0]), .fs_xor1(arrdiv32_fs86_xor1), .fs_or0(arrdiv32_fs86_or0));
  fs fs_arrdiv32_fs87_out(.a(arrdiv32_mux2to153_xor0[0]), .b(b[23]), .bin(arrdiv32_fs86_or0[0]), .fs_xor1(arrdiv32_fs87_xor1), .fs_or0(arrdiv32_fs87_or0));
  fs fs_arrdiv32_fs88_out(.a(arrdiv32_mux2to154_xor0[0]), .b(b[24]), .bin(arrdiv32_fs87_or0[0]), .fs_xor1(arrdiv32_fs88_xor1), .fs_or0(arrdiv32_fs88_or0));
  fs fs_arrdiv32_fs89_out(.a(arrdiv32_mux2to155_xor0[0]), .b(b[25]), .bin(arrdiv32_fs88_or0[0]), .fs_xor1(arrdiv32_fs89_xor1), .fs_or0(arrdiv32_fs89_or0));
  fs fs_arrdiv32_fs90_out(.a(arrdiv32_mux2to156_xor0[0]), .b(b[26]), .bin(arrdiv32_fs89_or0[0]), .fs_xor1(arrdiv32_fs90_xor1), .fs_or0(arrdiv32_fs90_or0));
  fs fs_arrdiv32_fs91_out(.a(arrdiv32_mux2to157_xor0[0]), .b(b[27]), .bin(arrdiv32_fs90_or0[0]), .fs_xor1(arrdiv32_fs91_xor1), .fs_or0(arrdiv32_fs91_or0));
  fs fs_arrdiv32_fs92_out(.a(arrdiv32_mux2to158_xor0[0]), .b(b[28]), .bin(arrdiv32_fs91_or0[0]), .fs_xor1(arrdiv32_fs92_xor1), .fs_or0(arrdiv32_fs92_or0));
  fs fs_arrdiv32_fs93_out(.a(arrdiv32_mux2to159_xor0[0]), .b(b[29]), .bin(arrdiv32_fs92_or0[0]), .fs_xor1(arrdiv32_fs93_xor1), .fs_or0(arrdiv32_fs93_or0));
  fs fs_arrdiv32_fs94_out(.a(arrdiv32_mux2to160_xor0[0]), .b(b[30]), .bin(arrdiv32_fs93_or0[0]), .fs_xor1(arrdiv32_fs94_xor1), .fs_or0(arrdiv32_fs94_or0));
  fs fs_arrdiv32_fs95_out(.a(arrdiv32_mux2to161_xor0[0]), .b(b[31]), .bin(arrdiv32_fs94_or0[0]), .fs_xor1(arrdiv32_fs95_xor1), .fs_or0(arrdiv32_fs95_or0));
  mux2to1 mux2to1_arrdiv32_mux2to162_out(.d0(arrdiv32_fs64_xor0[0]), .d1(a[29]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to162_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to163_out(.d0(arrdiv32_fs65_xor1[0]), .d1(arrdiv32_mux2to131_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to163_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to164_out(.d0(arrdiv32_fs66_xor1[0]), .d1(arrdiv32_mux2to132_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to164_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to165_out(.d0(arrdiv32_fs67_xor1[0]), .d1(arrdiv32_mux2to133_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to165_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to166_out(.d0(arrdiv32_fs68_xor1[0]), .d1(arrdiv32_mux2to134_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to166_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to167_out(.d0(arrdiv32_fs69_xor1[0]), .d1(arrdiv32_mux2to135_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to167_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to168_out(.d0(arrdiv32_fs70_xor1[0]), .d1(arrdiv32_mux2to136_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to168_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to169_out(.d0(arrdiv32_fs71_xor1[0]), .d1(arrdiv32_mux2to137_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to169_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to170_out(.d0(arrdiv32_fs72_xor1[0]), .d1(arrdiv32_mux2to138_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to170_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to171_out(.d0(arrdiv32_fs73_xor1[0]), .d1(arrdiv32_mux2to139_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to171_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to172_out(.d0(arrdiv32_fs74_xor1[0]), .d1(arrdiv32_mux2to140_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to172_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to173_out(.d0(arrdiv32_fs75_xor1[0]), .d1(arrdiv32_mux2to141_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to173_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to174_out(.d0(arrdiv32_fs76_xor1[0]), .d1(arrdiv32_mux2to142_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to174_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to175_out(.d0(arrdiv32_fs77_xor1[0]), .d1(arrdiv32_mux2to143_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to175_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to176_out(.d0(arrdiv32_fs78_xor1[0]), .d1(arrdiv32_mux2to144_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to176_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to177_out(.d0(arrdiv32_fs79_xor1[0]), .d1(arrdiv32_mux2to145_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to177_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to178_out(.d0(arrdiv32_fs80_xor1[0]), .d1(arrdiv32_mux2to146_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to178_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to179_out(.d0(arrdiv32_fs81_xor1[0]), .d1(arrdiv32_mux2to147_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to179_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to180_out(.d0(arrdiv32_fs82_xor1[0]), .d1(arrdiv32_mux2to148_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to180_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to181_out(.d0(arrdiv32_fs83_xor1[0]), .d1(arrdiv32_mux2to149_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to181_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to182_out(.d0(arrdiv32_fs84_xor1[0]), .d1(arrdiv32_mux2to150_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to182_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to183_out(.d0(arrdiv32_fs85_xor1[0]), .d1(arrdiv32_mux2to151_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to183_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to184_out(.d0(arrdiv32_fs86_xor1[0]), .d1(arrdiv32_mux2to152_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to184_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to185_out(.d0(arrdiv32_fs87_xor1[0]), .d1(arrdiv32_mux2to153_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to185_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to186_out(.d0(arrdiv32_fs88_xor1[0]), .d1(arrdiv32_mux2to154_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to186_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to187_out(.d0(arrdiv32_fs89_xor1[0]), .d1(arrdiv32_mux2to155_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to187_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to188_out(.d0(arrdiv32_fs90_xor1[0]), .d1(arrdiv32_mux2to156_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to188_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to189_out(.d0(arrdiv32_fs91_xor1[0]), .d1(arrdiv32_mux2to157_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to189_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to190_out(.d0(arrdiv32_fs92_xor1[0]), .d1(arrdiv32_mux2to158_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to190_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to191_out(.d0(arrdiv32_fs93_xor1[0]), .d1(arrdiv32_mux2to159_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to191_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to192_out(.d0(arrdiv32_fs94_xor1[0]), .d1(arrdiv32_mux2to160_xor0[0]), .sel(arrdiv32_fs95_or0[0]), .mux2to1_xor0(arrdiv32_mux2to192_xor0));
  not_gate not_gate_arrdiv32_not2(.a(arrdiv32_fs95_or0[0]), .out(arrdiv32_not2));
  fs fs_arrdiv32_fs96_out(.a(a[28]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs96_xor0), .fs_or0(arrdiv32_fs96_and0));
  fs fs_arrdiv32_fs97_out(.a(arrdiv32_mux2to162_xor0[0]), .b(b[1]), .bin(arrdiv32_fs96_and0[0]), .fs_xor1(arrdiv32_fs97_xor1), .fs_or0(arrdiv32_fs97_or0));
  fs fs_arrdiv32_fs98_out(.a(arrdiv32_mux2to163_xor0[0]), .b(b[2]), .bin(arrdiv32_fs97_or0[0]), .fs_xor1(arrdiv32_fs98_xor1), .fs_or0(arrdiv32_fs98_or0));
  fs fs_arrdiv32_fs99_out(.a(arrdiv32_mux2to164_xor0[0]), .b(b[3]), .bin(arrdiv32_fs98_or0[0]), .fs_xor1(arrdiv32_fs99_xor1), .fs_or0(arrdiv32_fs99_or0));
  fs fs_arrdiv32_fs100_out(.a(arrdiv32_mux2to165_xor0[0]), .b(b[4]), .bin(arrdiv32_fs99_or0[0]), .fs_xor1(arrdiv32_fs100_xor1), .fs_or0(arrdiv32_fs100_or0));
  fs fs_arrdiv32_fs101_out(.a(arrdiv32_mux2to166_xor0[0]), .b(b[5]), .bin(arrdiv32_fs100_or0[0]), .fs_xor1(arrdiv32_fs101_xor1), .fs_or0(arrdiv32_fs101_or0));
  fs fs_arrdiv32_fs102_out(.a(arrdiv32_mux2to167_xor0[0]), .b(b[6]), .bin(arrdiv32_fs101_or0[0]), .fs_xor1(arrdiv32_fs102_xor1), .fs_or0(arrdiv32_fs102_or0));
  fs fs_arrdiv32_fs103_out(.a(arrdiv32_mux2to168_xor0[0]), .b(b[7]), .bin(arrdiv32_fs102_or0[0]), .fs_xor1(arrdiv32_fs103_xor1), .fs_or0(arrdiv32_fs103_or0));
  fs fs_arrdiv32_fs104_out(.a(arrdiv32_mux2to169_xor0[0]), .b(b[8]), .bin(arrdiv32_fs103_or0[0]), .fs_xor1(arrdiv32_fs104_xor1), .fs_or0(arrdiv32_fs104_or0));
  fs fs_arrdiv32_fs105_out(.a(arrdiv32_mux2to170_xor0[0]), .b(b[9]), .bin(arrdiv32_fs104_or0[0]), .fs_xor1(arrdiv32_fs105_xor1), .fs_or0(arrdiv32_fs105_or0));
  fs fs_arrdiv32_fs106_out(.a(arrdiv32_mux2to171_xor0[0]), .b(b[10]), .bin(arrdiv32_fs105_or0[0]), .fs_xor1(arrdiv32_fs106_xor1), .fs_or0(arrdiv32_fs106_or0));
  fs fs_arrdiv32_fs107_out(.a(arrdiv32_mux2to172_xor0[0]), .b(b[11]), .bin(arrdiv32_fs106_or0[0]), .fs_xor1(arrdiv32_fs107_xor1), .fs_or0(arrdiv32_fs107_or0));
  fs fs_arrdiv32_fs108_out(.a(arrdiv32_mux2to173_xor0[0]), .b(b[12]), .bin(arrdiv32_fs107_or0[0]), .fs_xor1(arrdiv32_fs108_xor1), .fs_or0(arrdiv32_fs108_or0));
  fs fs_arrdiv32_fs109_out(.a(arrdiv32_mux2to174_xor0[0]), .b(b[13]), .bin(arrdiv32_fs108_or0[0]), .fs_xor1(arrdiv32_fs109_xor1), .fs_or0(arrdiv32_fs109_or0));
  fs fs_arrdiv32_fs110_out(.a(arrdiv32_mux2to175_xor0[0]), .b(b[14]), .bin(arrdiv32_fs109_or0[0]), .fs_xor1(arrdiv32_fs110_xor1), .fs_or0(arrdiv32_fs110_or0));
  fs fs_arrdiv32_fs111_out(.a(arrdiv32_mux2to176_xor0[0]), .b(b[15]), .bin(arrdiv32_fs110_or0[0]), .fs_xor1(arrdiv32_fs111_xor1), .fs_or0(arrdiv32_fs111_or0));
  fs fs_arrdiv32_fs112_out(.a(arrdiv32_mux2to177_xor0[0]), .b(b[16]), .bin(arrdiv32_fs111_or0[0]), .fs_xor1(arrdiv32_fs112_xor1), .fs_or0(arrdiv32_fs112_or0));
  fs fs_arrdiv32_fs113_out(.a(arrdiv32_mux2to178_xor0[0]), .b(b[17]), .bin(arrdiv32_fs112_or0[0]), .fs_xor1(arrdiv32_fs113_xor1), .fs_or0(arrdiv32_fs113_or0));
  fs fs_arrdiv32_fs114_out(.a(arrdiv32_mux2to179_xor0[0]), .b(b[18]), .bin(arrdiv32_fs113_or0[0]), .fs_xor1(arrdiv32_fs114_xor1), .fs_or0(arrdiv32_fs114_or0));
  fs fs_arrdiv32_fs115_out(.a(arrdiv32_mux2to180_xor0[0]), .b(b[19]), .bin(arrdiv32_fs114_or0[0]), .fs_xor1(arrdiv32_fs115_xor1), .fs_or0(arrdiv32_fs115_or0));
  fs fs_arrdiv32_fs116_out(.a(arrdiv32_mux2to181_xor0[0]), .b(b[20]), .bin(arrdiv32_fs115_or0[0]), .fs_xor1(arrdiv32_fs116_xor1), .fs_or0(arrdiv32_fs116_or0));
  fs fs_arrdiv32_fs117_out(.a(arrdiv32_mux2to182_xor0[0]), .b(b[21]), .bin(arrdiv32_fs116_or0[0]), .fs_xor1(arrdiv32_fs117_xor1), .fs_or0(arrdiv32_fs117_or0));
  fs fs_arrdiv32_fs118_out(.a(arrdiv32_mux2to183_xor0[0]), .b(b[22]), .bin(arrdiv32_fs117_or0[0]), .fs_xor1(arrdiv32_fs118_xor1), .fs_or0(arrdiv32_fs118_or0));
  fs fs_arrdiv32_fs119_out(.a(arrdiv32_mux2to184_xor0[0]), .b(b[23]), .bin(arrdiv32_fs118_or0[0]), .fs_xor1(arrdiv32_fs119_xor1), .fs_or0(arrdiv32_fs119_or0));
  fs fs_arrdiv32_fs120_out(.a(arrdiv32_mux2to185_xor0[0]), .b(b[24]), .bin(arrdiv32_fs119_or0[0]), .fs_xor1(arrdiv32_fs120_xor1), .fs_or0(arrdiv32_fs120_or0));
  fs fs_arrdiv32_fs121_out(.a(arrdiv32_mux2to186_xor0[0]), .b(b[25]), .bin(arrdiv32_fs120_or0[0]), .fs_xor1(arrdiv32_fs121_xor1), .fs_or0(arrdiv32_fs121_or0));
  fs fs_arrdiv32_fs122_out(.a(arrdiv32_mux2to187_xor0[0]), .b(b[26]), .bin(arrdiv32_fs121_or0[0]), .fs_xor1(arrdiv32_fs122_xor1), .fs_or0(arrdiv32_fs122_or0));
  fs fs_arrdiv32_fs123_out(.a(arrdiv32_mux2to188_xor0[0]), .b(b[27]), .bin(arrdiv32_fs122_or0[0]), .fs_xor1(arrdiv32_fs123_xor1), .fs_or0(arrdiv32_fs123_or0));
  fs fs_arrdiv32_fs124_out(.a(arrdiv32_mux2to189_xor0[0]), .b(b[28]), .bin(arrdiv32_fs123_or0[0]), .fs_xor1(arrdiv32_fs124_xor1), .fs_or0(arrdiv32_fs124_or0));
  fs fs_arrdiv32_fs125_out(.a(arrdiv32_mux2to190_xor0[0]), .b(b[29]), .bin(arrdiv32_fs124_or0[0]), .fs_xor1(arrdiv32_fs125_xor1), .fs_or0(arrdiv32_fs125_or0));
  fs fs_arrdiv32_fs126_out(.a(arrdiv32_mux2to191_xor0[0]), .b(b[30]), .bin(arrdiv32_fs125_or0[0]), .fs_xor1(arrdiv32_fs126_xor1), .fs_or0(arrdiv32_fs126_or0));
  fs fs_arrdiv32_fs127_out(.a(arrdiv32_mux2to192_xor0[0]), .b(b[31]), .bin(arrdiv32_fs126_or0[0]), .fs_xor1(arrdiv32_fs127_xor1), .fs_or0(arrdiv32_fs127_or0));
  mux2to1 mux2to1_arrdiv32_mux2to193_out(.d0(arrdiv32_fs96_xor0[0]), .d1(a[28]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to193_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to194_out(.d0(arrdiv32_fs97_xor1[0]), .d1(arrdiv32_mux2to162_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to194_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to195_out(.d0(arrdiv32_fs98_xor1[0]), .d1(arrdiv32_mux2to163_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to195_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to196_out(.d0(arrdiv32_fs99_xor1[0]), .d1(arrdiv32_mux2to164_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to196_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to197_out(.d0(arrdiv32_fs100_xor1[0]), .d1(arrdiv32_mux2to165_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to197_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to198_out(.d0(arrdiv32_fs101_xor1[0]), .d1(arrdiv32_mux2to166_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to198_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to199_out(.d0(arrdiv32_fs102_xor1[0]), .d1(arrdiv32_mux2to167_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to199_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1100_out(.d0(arrdiv32_fs103_xor1[0]), .d1(arrdiv32_mux2to168_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1100_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1101_out(.d0(arrdiv32_fs104_xor1[0]), .d1(arrdiv32_mux2to169_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1101_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1102_out(.d0(arrdiv32_fs105_xor1[0]), .d1(arrdiv32_mux2to170_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1102_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1103_out(.d0(arrdiv32_fs106_xor1[0]), .d1(arrdiv32_mux2to171_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1103_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1104_out(.d0(arrdiv32_fs107_xor1[0]), .d1(arrdiv32_mux2to172_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1104_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1105_out(.d0(arrdiv32_fs108_xor1[0]), .d1(arrdiv32_mux2to173_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1105_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1106_out(.d0(arrdiv32_fs109_xor1[0]), .d1(arrdiv32_mux2to174_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1106_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1107_out(.d0(arrdiv32_fs110_xor1[0]), .d1(arrdiv32_mux2to175_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1107_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1108_out(.d0(arrdiv32_fs111_xor1[0]), .d1(arrdiv32_mux2to176_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1108_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1109_out(.d0(arrdiv32_fs112_xor1[0]), .d1(arrdiv32_mux2to177_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1109_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1110_out(.d0(arrdiv32_fs113_xor1[0]), .d1(arrdiv32_mux2to178_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1110_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1111_out(.d0(arrdiv32_fs114_xor1[0]), .d1(arrdiv32_mux2to179_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1111_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1112_out(.d0(arrdiv32_fs115_xor1[0]), .d1(arrdiv32_mux2to180_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1112_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1113_out(.d0(arrdiv32_fs116_xor1[0]), .d1(arrdiv32_mux2to181_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1113_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1114_out(.d0(arrdiv32_fs117_xor1[0]), .d1(arrdiv32_mux2to182_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1114_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1115_out(.d0(arrdiv32_fs118_xor1[0]), .d1(arrdiv32_mux2to183_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1115_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1116_out(.d0(arrdiv32_fs119_xor1[0]), .d1(arrdiv32_mux2to184_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1116_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1117_out(.d0(arrdiv32_fs120_xor1[0]), .d1(arrdiv32_mux2to185_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1117_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1118_out(.d0(arrdiv32_fs121_xor1[0]), .d1(arrdiv32_mux2to186_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1118_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1119_out(.d0(arrdiv32_fs122_xor1[0]), .d1(arrdiv32_mux2to187_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1119_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1120_out(.d0(arrdiv32_fs123_xor1[0]), .d1(arrdiv32_mux2to188_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1120_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1121_out(.d0(arrdiv32_fs124_xor1[0]), .d1(arrdiv32_mux2to189_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1121_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1122_out(.d0(arrdiv32_fs125_xor1[0]), .d1(arrdiv32_mux2to190_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1122_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1123_out(.d0(arrdiv32_fs126_xor1[0]), .d1(arrdiv32_mux2to191_xor0[0]), .sel(arrdiv32_fs127_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1123_xor0));
  not_gate not_gate_arrdiv32_not3(.a(arrdiv32_fs127_or0[0]), .out(arrdiv32_not3));
  fs fs_arrdiv32_fs128_out(.a(a[27]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs128_xor0), .fs_or0(arrdiv32_fs128_and0));
  fs fs_arrdiv32_fs129_out(.a(arrdiv32_mux2to193_xor0[0]), .b(b[1]), .bin(arrdiv32_fs128_and0[0]), .fs_xor1(arrdiv32_fs129_xor1), .fs_or0(arrdiv32_fs129_or0));
  fs fs_arrdiv32_fs130_out(.a(arrdiv32_mux2to194_xor0[0]), .b(b[2]), .bin(arrdiv32_fs129_or0[0]), .fs_xor1(arrdiv32_fs130_xor1), .fs_or0(arrdiv32_fs130_or0));
  fs fs_arrdiv32_fs131_out(.a(arrdiv32_mux2to195_xor0[0]), .b(b[3]), .bin(arrdiv32_fs130_or0[0]), .fs_xor1(arrdiv32_fs131_xor1), .fs_or0(arrdiv32_fs131_or0));
  fs fs_arrdiv32_fs132_out(.a(arrdiv32_mux2to196_xor0[0]), .b(b[4]), .bin(arrdiv32_fs131_or0[0]), .fs_xor1(arrdiv32_fs132_xor1), .fs_or0(arrdiv32_fs132_or0));
  fs fs_arrdiv32_fs133_out(.a(arrdiv32_mux2to197_xor0[0]), .b(b[5]), .bin(arrdiv32_fs132_or0[0]), .fs_xor1(arrdiv32_fs133_xor1), .fs_or0(arrdiv32_fs133_or0));
  fs fs_arrdiv32_fs134_out(.a(arrdiv32_mux2to198_xor0[0]), .b(b[6]), .bin(arrdiv32_fs133_or0[0]), .fs_xor1(arrdiv32_fs134_xor1), .fs_or0(arrdiv32_fs134_or0));
  fs fs_arrdiv32_fs135_out(.a(arrdiv32_mux2to199_xor0[0]), .b(b[7]), .bin(arrdiv32_fs134_or0[0]), .fs_xor1(arrdiv32_fs135_xor1), .fs_or0(arrdiv32_fs135_or0));
  fs fs_arrdiv32_fs136_out(.a(arrdiv32_mux2to1100_xor0[0]), .b(b[8]), .bin(arrdiv32_fs135_or0[0]), .fs_xor1(arrdiv32_fs136_xor1), .fs_or0(arrdiv32_fs136_or0));
  fs fs_arrdiv32_fs137_out(.a(arrdiv32_mux2to1101_xor0[0]), .b(b[9]), .bin(arrdiv32_fs136_or0[0]), .fs_xor1(arrdiv32_fs137_xor1), .fs_or0(arrdiv32_fs137_or0));
  fs fs_arrdiv32_fs138_out(.a(arrdiv32_mux2to1102_xor0[0]), .b(b[10]), .bin(arrdiv32_fs137_or0[0]), .fs_xor1(arrdiv32_fs138_xor1), .fs_or0(arrdiv32_fs138_or0));
  fs fs_arrdiv32_fs139_out(.a(arrdiv32_mux2to1103_xor0[0]), .b(b[11]), .bin(arrdiv32_fs138_or0[0]), .fs_xor1(arrdiv32_fs139_xor1), .fs_or0(arrdiv32_fs139_or0));
  fs fs_arrdiv32_fs140_out(.a(arrdiv32_mux2to1104_xor0[0]), .b(b[12]), .bin(arrdiv32_fs139_or0[0]), .fs_xor1(arrdiv32_fs140_xor1), .fs_or0(arrdiv32_fs140_or0));
  fs fs_arrdiv32_fs141_out(.a(arrdiv32_mux2to1105_xor0[0]), .b(b[13]), .bin(arrdiv32_fs140_or0[0]), .fs_xor1(arrdiv32_fs141_xor1), .fs_or0(arrdiv32_fs141_or0));
  fs fs_arrdiv32_fs142_out(.a(arrdiv32_mux2to1106_xor0[0]), .b(b[14]), .bin(arrdiv32_fs141_or0[0]), .fs_xor1(arrdiv32_fs142_xor1), .fs_or0(arrdiv32_fs142_or0));
  fs fs_arrdiv32_fs143_out(.a(arrdiv32_mux2to1107_xor0[0]), .b(b[15]), .bin(arrdiv32_fs142_or0[0]), .fs_xor1(arrdiv32_fs143_xor1), .fs_or0(arrdiv32_fs143_or0));
  fs fs_arrdiv32_fs144_out(.a(arrdiv32_mux2to1108_xor0[0]), .b(b[16]), .bin(arrdiv32_fs143_or0[0]), .fs_xor1(arrdiv32_fs144_xor1), .fs_or0(arrdiv32_fs144_or0));
  fs fs_arrdiv32_fs145_out(.a(arrdiv32_mux2to1109_xor0[0]), .b(b[17]), .bin(arrdiv32_fs144_or0[0]), .fs_xor1(arrdiv32_fs145_xor1), .fs_or0(arrdiv32_fs145_or0));
  fs fs_arrdiv32_fs146_out(.a(arrdiv32_mux2to1110_xor0[0]), .b(b[18]), .bin(arrdiv32_fs145_or0[0]), .fs_xor1(arrdiv32_fs146_xor1), .fs_or0(arrdiv32_fs146_or0));
  fs fs_arrdiv32_fs147_out(.a(arrdiv32_mux2to1111_xor0[0]), .b(b[19]), .bin(arrdiv32_fs146_or0[0]), .fs_xor1(arrdiv32_fs147_xor1), .fs_or0(arrdiv32_fs147_or0));
  fs fs_arrdiv32_fs148_out(.a(arrdiv32_mux2to1112_xor0[0]), .b(b[20]), .bin(arrdiv32_fs147_or0[0]), .fs_xor1(arrdiv32_fs148_xor1), .fs_or0(arrdiv32_fs148_or0));
  fs fs_arrdiv32_fs149_out(.a(arrdiv32_mux2to1113_xor0[0]), .b(b[21]), .bin(arrdiv32_fs148_or0[0]), .fs_xor1(arrdiv32_fs149_xor1), .fs_or0(arrdiv32_fs149_or0));
  fs fs_arrdiv32_fs150_out(.a(arrdiv32_mux2to1114_xor0[0]), .b(b[22]), .bin(arrdiv32_fs149_or0[0]), .fs_xor1(arrdiv32_fs150_xor1), .fs_or0(arrdiv32_fs150_or0));
  fs fs_arrdiv32_fs151_out(.a(arrdiv32_mux2to1115_xor0[0]), .b(b[23]), .bin(arrdiv32_fs150_or0[0]), .fs_xor1(arrdiv32_fs151_xor1), .fs_or0(arrdiv32_fs151_or0));
  fs fs_arrdiv32_fs152_out(.a(arrdiv32_mux2to1116_xor0[0]), .b(b[24]), .bin(arrdiv32_fs151_or0[0]), .fs_xor1(arrdiv32_fs152_xor1), .fs_or0(arrdiv32_fs152_or0));
  fs fs_arrdiv32_fs153_out(.a(arrdiv32_mux2to1117_xor0[0]), .b(b[25]), .bin(arrdiv32_fs152_or0[0]), .fs_xor1(arrdiv32_fs153_xor1), .fs_or0(arrdiv32_fs153_or0));
  fs fs_arrdiv32_fs154_out(.a(arrdiv32_mux2to1118_xor0[0]), .b(b[26]), .bin(arrdiv32_fs153_or0[0]), .fs_xor1(arrdiv32_fs154_xor1), .fs_or0(arrdiv32_fs154_or0));
  fs fs_arrdiv32_fs155_out(.a(arrdiv32_mux2to1119_xor0[0]), .b(b[27]), .bin(arrdiv32_fs154_or0[0]), .fs_xor1(arrdiv32_fs155_xor1), .fs_or0(arrdiv32_fs155_or0));
  fs fs_arrdiv32_fs156_out(.a(arrdiv32_mux2to1120_xor0[0]), .b(b[28]), .bin(arrdiv32_fs155_or0[0]), .fs_xor1(arrdiv32_fs156_xor1), .fs_or0(arrdiv32_fs156_or0));
  fs fs_arrdiv32_fs157_out(.a(arrdiv32_mux2to1121_xor0[0]), .b(b[29]), .bin(arrdiv32_fs156_or0[0]), .fs_xor1(arrdiv32_fs157_xor1), .fs_or0(arrdiv32_fs157_or0));
  fs fs_arrdiv32_fs158_out(.a(arrdiv32_mux2to1122_xor0[0]), .b(b[30]), .bin(arrdiv32_fs157_or0[0]), .fs_xor1(arrdiv32_fs158_xor1), .fs_or0(arrdiv32_fs158_or0));
  fs fs_arrdiv32_fs159_out(.a(arrdiv32_mux2to1123_xor0[0]), .b(b[31]), .bin(arrdiv32_fs158_or0[0]), .fs_xor1(arrdiv32_fs159_xor1), .fs_or0(arrdiv32_fs159_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1124_out(.d0(arrdiv32_fs128_xor0[0]), .d1(a[27]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1124_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1125_out(.d0(arrdiv32_fs129_xor1[0]), .d1(arrdiv32_mux2to193_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1125_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1126_out(.d0(arrdiv32_fs130_xor1[0]), .d1(arrdiv32_mux2to194_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1126_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1127_out(.d0(arrdiv32_fs131_xor1[0]), .d1(arrdiv32_mux2to195_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1127_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1128_out(.d0(arrdiv32_fs132_xor1[0]), .d1(arrdiv32_mux2to196_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1128_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1129_out(.d0(arrdiv32_fs133_xor1[0]), .d1(arrdiv32_mux2to197_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1129_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1130_out(.d0(arrdiv32_fs134_xor1[0]), .d1(arrdiv32_mux2to198_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1130_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1131_out(.d0(arrdiv32_fs135_xor1[0]), .d1(arrdiv32_mux2to199_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1131_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1132_out(.d0(arrdiv32_fs136_xor1[0]), .d1(arrdiv32_mux2to1100_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1132_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1133_out(.d0(arrdiv32_fs137_xor1[0]), .d1(arrdiv32_mux2to1101_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1133_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1134_out(.d0(arrdiv32_fs138_xor1[0]), .d1(arrdiv32_mux2to1102_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1134_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1135_out(.d0(arrdiv32_fs139_xor1[0]), .d1(arrdiv32_mux2to1103_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1135_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1136_out(.d0(arrdiv32_fs140_xor1[0]), .d1(arrdiv32_mux2to1104_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1136_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1137_out(.d0(arrdiv32_fs141_xor1[0]), .d1(arrdiv32_mux2to1105_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1137_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1138_out(.d0(arrdiv32_fs142_xor1[0]), .d1(arrdiv32_mux2to1106_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1138_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1139_out(.d0(arrdiv32_fs143_xor1[0]), .d1(arrdiv32_mux2to1107_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1139_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1140_out(.d0(arrdiv32_fs144_xor1[0]), .d1(arrdiv32_mux2to1108_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1140_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1141_out(.d0(arrdiv32_fs145_xor1[0]), .d1(arrdiv32_mux2to1109_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1141_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1142_out(.d0(arrdiv32_fs146_xor1[0]), .d1(arrdiv32_mux2to1110_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1142_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1143_out(.d0(arrdiv32_fs147_xor1[0]), .d1(arrdiv32_mux2to1111_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1143_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1144_out(.d0(arrdiv32_fs148_xor1[0]), .d1(arrdiv32_mux2to1112_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1144_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1145_out(.d0(arrdiv32_fs149_xor1[0]), .d1(arrdiv32_mux2to1113_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1145_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1146_out(.d0(arrdiv32_fs150_xor1[0]), .d1(arrdiv32_mux2to1114_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1146_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1147_out(.d0(arrdiv32_fs151_xor1[0]), .d1(arrdiv32_mux2to1115_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1147_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1148_out(.d0(arrdiv32_fs152_xor1[0]), .d1(arrdiv32_mux2to1116_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1148_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1149_out(.d0(arrdiv32_fs153_xor1[0]), .d1(arrdiv32_mux2to1117_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1149_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1150_out(.d0(arrdiv32_fs154_xor1[0]), .d1(arrdiv32_mux2to1118_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1150_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1151_out(.d0(arrdiv32_fs155_xor1[0]), .d1(arrdiv32_mux2to1119_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1151_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1152_out(.d0(arrdiv32_fs156_xor1[0]), .d1(arrdiv32_mux2to1120_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1152_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1153_out(.d0(arrdiv32_fs157_xor1[0]), .d1(arrdiv32_mux2to1121_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1153_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1154_out(.d0(arrdiv32_fs158_xor1[0]), .d1(arrdiv32_mux2to1122_xor0[0]), .sel(arrdiv32_fs159_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1154_xor0));
  not_gate not_gate_arrdiv32_not4(.a(arrdiv32_fs159_or0[0]), .out(arrdiv32_not4));
  fs fs_arrdiv32_fs160_out(.a(a[26]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs160_xor0), .fs_or0(arrdiv32_fs160_and0));
  fs fs_arrdiv32_fs161_out(.a(arrdiv32_mux2to1124_xor0[0]), .b(b[1]), .bin(arrdiv32_fs160_and0[0]), .fs_xor1(arrdiv32_fs161_xor1), .fs_or0(arrdiv32_fs161_or0));
  fs fs_arrdiv32_fs162_out(.a(arrdiv32_mux2to1125_xor0[0]), .b(b[2]), .bin(arrdiv32_fs161_or0[0]), .fs_xor1(arrdiv32_fs162_xor1), .fs_or0(arrdiv32_fs162_or0));
  fs fs_arrdiv32_fs163_out(.a(arrdiv32_mux2to1126_xor0[0]), .b(b[3]), .bin(arrdiv32_fs162_or0[0]), .fs_xor1(arrdiv32_fs163_xor1), .fs_or0(arrdiv32_fs163_or0));
  fs fs_arrdiv32_fs164_out(.a(arrdiv32_mux2to1127_xor0[0]), .b(b[4]), .bin(arrdiv32_fs163_or0[0]), .fs_xor1(arrdiv32_fs164_xor1), .fs_or0(arrdiv32_fs164_or0));
  fs fs_arrdiv32_fs165_out(.a(arrdiv32_mux2to1128_xor0[0]), .b(b[5]), .bin(arrdiv32_fs164_or0[0]), .fs_xor1(arrdiv32_fs165_xor1), .fs_or0(arrdiv32_fs165_or0));
  fs fs_arrdiv32_fs166_out(.a(arrdiv32_mux2to1129_xor0[0]), .b(b[6]), .bin(arrdiv32_fs165_or0[0]), .fs_xor1(arrdiv32_fs166_xor1), .fs_or0(arrdiv32_fs166_or0));
  fs fs_arrdiv32_fs167_out(.a(arrdiv32_mux2to1130_xor0[0]), .b(b[7]), .bin(arrdiv32_fs166_or0[0]), .fs_xor1(arrdiv32_fs167_xor1), .fs_or0(arrdiv32_fs167_or0));
  fs fs_arrdiv32_fs168_out(.a(arrdiv32_mux2to1131_xor0[0]), .b(b[8]), .bin(arrdiv32_fs167_or0[0]), .fs_xor1(arrdiv32_fs168_xor1), .fs_or0(arrdiv32_fs168_or0));
  fs fs_arrdiv32_fs169_out(.a(arrdiv32_mux2to1132_xor0[0]), .b(b[9]), .bin(arrdiv32_fs168_or0[0]), .fs_xor1(arrdiv32_fs169_xor1), .fs_or0(arrdiv32_fs169_or0));
  fs fs_arrdiv32_fs170_out(.a(arrdiv32_mux2to1133_xor0[0]), .b(b[10]), .bin(arrdiv32_fs169_or0[0]), .fs_xor1(arrdiv32_fs170_xor1), .fs_or0(arrdiv32_fs170_or0));
  fs fs_arrdiv32_fs171_out(.a(arrdiv32_mux2to1134_xor0[0]), .b(b[11]), .bin(arrdiv32_fs170_or0[0]), .fs_xor1(arrdiv32_fs171_xor1), .fs_or0(arrdiv32_fs171_or0));
  fs fs_arrdiv32_fs172_out(.a(arrdiv32_mux2to1135_xor0[0]), .b(b[12]), .bin(arrdiv32_fs171_or0[0]), .fs_xor1(arrdiv32_fs172_xor1), .fs_or0(arrdiv32_fs172_or0));
  fs fs_arrdiv32_fs173_out(.a(arrdiv32_mux2to1136_xor0[0]), .b(b[13]), .bin(arrdiv32_fs172_or0[0]), .fs_xor1(arrdiv32_fs173_xor1), .fs_or0(arrdiv32_fs173_or0));
  fs fs_arrdiv32_fs174_out(.a(arrdiv32_mux2to1137_xor0[0]), .b(b[14]), .bin(arrdiv32_fs173_or0[0]), .fs_xor1(arrdiv32_fs174_xor1), .fs_or0(arrdiv32_fs174_or0));
  fs fs_arrdiv32_fs175_out(.a(arrdiv32_mux2to1138_xor0[0]), .b(b[15]), .bin(arrdiv32_fs174_or0[0]), .fs_xor1(arrdiv32_fs175_xor1), .fs_or0(arrdiv32_fs175_or0));
  fs fs_arrdiv32_fs176_out(.a(arrdiv32_mux2to1139_xor0[0]), .b(b[16]), .bin(arrdiv32_fs175_or0[0]), .fs_xor1(arrdiv32_fs176_xor1), .fs_or0(arrdiv32_fs176_or0));
  fs fs_arrdiv32_fs177_out(.a(arrdiv32_mux2to1140_xor0[0]), .b(b[17]), .bin(arrdiv32_fs176_or0[0]), .fs_xor1(arrdiv32_fs177_xor1), .fs_or0(arrdiv32_fs177_or0));
  fs fs_arrdiv32_fs178_out(.a(arrdiv32_mux2to1141_xor0[0]), .b(b[18]), .bin(arrdiv32_fs177_or0[0]), .fs_xor1(arrdiv32_fs178_xor1), .fs_or0(arrdiv32_fs178_or0));
  fs fs_arrdiv32_fs179_out(.a(arrdiv32_mux2to1142_xor0[0]), .b(b[19]), .bin(arrdiv32_fs178_or0[0]), .fs_xor1(arrdiv32_fs179_xor1), .fs_or0(arrdiv32_fs179_or0));
  fs fs_arrdiv32_fs180_out(.a(arrdiv32_mux2to1143_xor0[0]), .b(b[20]), .bin(arrdiv32_fs179_or0[0]), .fs_xor1(arrdiv32_fs180_xor1), .fs_or0(arrdiv32_fs180_or0));
  fs fs_arrdiv32_fs181_out(.a(arrdiv32_mux2to1144_xor0[0]), .b(b[21]), .bin(arrdiv32_fs180_or0[0]), .fs_xor1(arrdiv32_fs181_xor1), .fs_or0(arrdiv32_fs181_or0));
  fs fs_arrdiv32_fs182_out(.a(arrdiv32_mux2to1145_xor0[0]), .b(b[22]), .bin(arrdiv32_fs181_or0[0]), .fs_xor1(arrdiv32_fs182_xor1), .fs_or0(arrdiv32_fs182_or0));
  fs fs_arrdiv32_fs183_out(.a(arrdiv32_mux2to1146_xor0[0]), .b(b[23]), .bin(arrdiv32_fs182_or0[0]), .fs_xor1(arrdiv32_fs183_xor1), .fs_or0(arrdiv32_fs183_or0));
  fs fs_arrdiv32_fs184_out(.a(arrdiv32_mux2to1147_xor0[0]), .b(b[24]), .bin(arrdiv32_fs183_or0[0]), .fs_xor1(arrdiv32_fs184_xor1), .fs_or0(arrdiv32_fs184_or0));
  fs fs_arrdiv32_fs185_out(.a(arrdiv32_mux2to1148_xor0[0]), .b(b[25]), .bin(arrdiv32_fs184_or0[0]), .fs_xor1(arrdiv32_fs185_xor1), .fs_or0(arrdiv32_fs185_or0));
  fs fs_arrdiv32_fs186_out(.a(arrdiv32_mux2to1149_xor0[0]), .b(b[26]), .bin(arrdiv32_fs185_or0[0]), .fs_xor1(arrdiv32_fs186_xor1), .fs_or0(arrdiv32_fs186_or0));
  fs fs_arrdiv32_fs187_out(.a(arrdiv32_mux2to1150_xor0[0]), .b(b[27]), .bin(arrdiv32_fs186_or0[0]), .fs_xor1(arrdiv32_fs187_xor1), .fs_or0(arrdiv32_fs187_or0));
  fs fs_arrdiv32_fs188_out(.a(arrdiv32_mux2to1151_xor0[0]), .b(b[28]), .bin(arrdiv32_fs187_or0[0]), .fs_xor1(arrdiv32_fs188_xor1), .fs_or0(arrdiv32_fs188_or0));
  fs fs_arrdiv32_fs189_out(.a(arrdiv32_mux2to1152_xor0[0]), .b(b[29]), .bin(arrdiv32_fs188_or0[0]), .fs_xor1(arrdiv32_fs189_xor1), .fs_or0(arrdiv32_fs189_or0));
  fs fs_arrdiv32_fs190_out(.a(arrdiv32_mux2to1153_xor0[0]), .b(b[30]), .bin(arrdiv32_fs189_or0[0]), .fs_xor1(arrdiv32_fs190_xor1), .fs_or0(arrdiv32_fs190_or0));
  fs fs_arrdiv32_fs191_out(.a(arrdiv32_mux2to1154_xor0[0]), .b(b[31]), .bin(arrdiv32_fs190_or0[0]), .fs_xor1(arrdiv32_fs191_xor1), .fs_or0(arrdiv32_fs191_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1155_out(.d0(arrdiv32_fs160_xor0[0]), .d1(a[26]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1155_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1156_out(.d0(arrdiv32_fs161_xor1[0]), .d1(arrdiv32_mux2to1124_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1156_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1157_out(.d0(arrdiv32_fs162_xor1[0]), .d1(arrdiv32_mux2to1125_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1157_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1158_out(.d0(arrdiv32_fs163_xor1[0]), .d1(arrdiv32_mux2to1126_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1158_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1159_out(.d0(arrdiv32_fs164_xor1[0]), .d1(arrdiv32_mux2to1127_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1159_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1160_out(.d0(arrdiv32_fs165_xor1[0]), .d1(arrdiv32_mux2to1128_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1160_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1161_out(.d0(arrdiv32_fs166_xor1[0]), .d1(arrdiv32_mux2to1129_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1161_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1162_out(.d0(arrdiv32_fs167_xor1[0]), .d1(arrdiv32_mux2to1130_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1162_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1163_out(.d0(arrdiv32_fs168_xor1[0]), .d1(arrdiv32_mux2to1131_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1163_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1164_out(.d0(arrdiv32_fs169_xor1[0]), .d1(arrdiv32_mux2to1132_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1164_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1165_out(.d0(arrdiv32_fs170_xor1[0]), .d1(arrdiv32_mux2to1133_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1165_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1166_out(.d0(arrdiv32_fs171_xor1[0]), .d1(arrdiv32_mux2to1134_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1166_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1167_out(.d0(arrdiv32_fs172_xor1[0]), .d1(arrdiv32_mux2to1135_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1167_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1168_out(.d0(arrdiv32_fs173_xor1[0]), .d1(arrdiv32_mux2to1136_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1168_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1169_out(.d0(arrdiv32_fs174_xor1[0]), .d1(arrdiv32_mux2to1137_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1169_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1170_out(.d0(arrdiv32_fs175_xor1[0]), .d1(arrdiv32_mux2to1138_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1170_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1171_out(.d0(arrdiv32_fs176_xor1[0]), .d1(arrdiv32_mux2to1139_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1171_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1172_out(.d0(arrdiv32_fs177_xor1[0]), .d1(arrdiv32_mux2to1140_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1172_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1173_out(.d0(arrdiv32_fs178_xor1[0]), .d1(arrdiv32_mux2to1141_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1173_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1174_out(.d0(arrdiv32_fs179_xor1[0]), .d1(arrdiv32_mux2to1142_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1174_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1175_out(.d0(arrdiv32_fs180_xor1[0]), .d1(arrdiv32_mux2to1143_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1175_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1176_out(.d0(arrdiv32_fs181_xor1[0]), .d1(arrdiv32_mux2to1144_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1176_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1177_out(.d0(arrdiv32_fs182_xor1[0]), .d1(arrdiv32_mux2to1145_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1177_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1178_out(.d0(arrdiv32_fs183_xor1[0]), .d1(arrdiv32_mux2to1146_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1178_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1179_out(.d0(arrdiv32_fs184_xor1[0]), .d1(arrdiv32_mux2to1147_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1179_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1180_out(.d0(arrdiv32_fs185_xor1[0]), .d1(arrdiv32_mux2to1148_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1180_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1181_out(.d0(arrdiv32_fs186_xor1[0]), .d1(arrdiv32_mux2to1149_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1181_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1182_out(.d0(arrdiv32_fs187_xor1[0]), .d1(arrdiv32_mux2to1150_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1182_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1183_out(.d0(arrdiv32_fs188_xor1[0]), .d1(arrdiv32_mux2to1151_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1183_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1184_out(.d0(arrdiv32_fs189_xor1[0]), .d1(arrdiv32_mux2to1152_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1184_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1185_out(.d0(arrdiv32_fs190_xor1[0]), .d1(arrdiv32_mux2to1153_xor0[0]), .sel(arrdiv32_fs191_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1185_xor0));
  not_gate not_gate_arrdiv32_not5(.a(arrdiv32_fs191_or0[0]), .out(arrdiv32_not5));
  fs fs_arrdiv32_fs192_out(.a(a[25]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs192_xor0), .fs_or0(arrdiv32_fs192_and0));
  fs fs_arrdiv32_fs193_out(.a(arrdiv32_mux2to1155_xor0[0]), .b(b[1]), .bin(arrdiv32_fs192_and0[0]), .fs_xor1(arrdiv32_fs193_xor1), .fs_or0(arrdiv32_fs193_or0));
  fs fs_arrdiv32_fs194_out(.a(arrdiv32_mux2to1156_xor0[0]), .b(b[2]), .bin(arrdiv32_fs193_or0[0]), .fs_xor1(arrdiv32_fs194_xor1), .fs_or0(arrdiv32_fs194_or0));
  fs fs_arrdiv32_fs195_out(.a(arrdiv32_mux2to1157_xor0[0]), .b(b[3]), .bin(arrdiv32_fs194_or0[0]), .fs_xor1(arrdiv32_fs195_xor1), .fs_or0(arrdiv32_fs195_or0));
  fs fs_arrdiv32_fs196_out(.a(arrdiv32_mux2to1158_xor0[0]), .b(b[4]), .bin(arrdiv32_fs195_or0[0]), .fs_xor1(arrdiv32_fs196_xor1), .fs_or0(arrdiv32_fs196_or0));
  fs fs_arrdiv32_fs197_out(.a(arrdiv32_mux2to1159_xor0[0]), .b(b[5]), .bin(arrdiv32_fs196_or0[0]), .fs_xor1(arrdiv32_fs197_xor1), .fs_or0(arrdiv32_fs197_or0));
  fs fs_arrdiv32_fs198_out(.a(arrdiv32_mux2to1160_xor0[0]), .b(b[6]), .bin(arrdiv32_fs197_or0[0]), .fs_xor1(arrdiv32_fs198_xor1), .fs_or0(arrdiv32_fs198_or0));
  fs fs_arrdiv32_fs199_out(.a(arrdiv32_mux2to1161_xor0[0]), .b(b[7]), .bin(arrdiv32_fs198_or0[0]), .fs_xor1(arrdiv32_fs199_xor1), .fs_or0(arrdiv32_fs199_or0));
  fs fs_arrdiv32_fs200_out(.a(arrdiv32_mux2to1162_xor0[0]), .b(b[8]), .bin(arrdiv32_fs199_or0[0]), .fs_xor1(arrdiv32_fs200_xor1), .fs_or0(arrdiv32_fs200_or0));
  fs fs_arrdiv32_fs201_out(.a(arrdiv32_mux2to1163_xor0[0]), .b(b[9]), .bin(arrdiv32_fs200_or0[0]), .fs_xor1(arrdiv32_fs201_xor1), .fs_or0(arrdiv32_fs201_or0));
  fs fs_arrdiv32_fs202_out(.a(arrdiv32_mux2to1164_xor0[0]), .b(b[10]), .bin(arrdiv32_fs201_or0[0]), .fs_xor1(arrdiv32_fs202_xor1), .fs_or0(arrdiv32_fs202_or0));
  fs fs_arrdiv32_fs203_out(.a(arrdiv32_mux2to1165_xor0[0]), .b(b[11]), .bin(arrdiv32_fs202_or0[0]), .fs_xor1(arrdiv32_fs203_xor1), .fs_or0(arrdiv32_fs203_or0));
  fs fs_arrdiv32_fs204_out(.a(arrdiv32_mux2to1166_xor0[0]), .b(b[12]), .bin(arrdiv32_fs203_or0[0]), .fs_xor1(arrdiv32_fs204_xor1), .fs_or0(arrdiv32_fs204_or0));
  fs fs_arrdiv32_fs205_out(.a(arrdiv32_mux2to1167_xor0[0]), .b(b[13]), .bin(arrdiv32_fs204_or0[0]), .fs_xor1(arrdiv32_fs205_xor1), .fs_or0(arrdiv32_fs205_or0));
  fs fs_arrdiv32_fs206_out(.a(arrdiv32_mux2to1168_xor0[0]), .b(b[14]), .bin(arrdiv32_fs205_or0[0]), .fs_xor1(arrdiv32_fs206_xor1), .fs_or0(arrdiv32_fs206_or0));
  fs fs_arrdiv32_fs207_out(.a(arrdiv32_mux2to1169_xor0[0]), .b(b[15]), .bin(arrdiv32_fs206_or0[0]), .fs_xor1(arrdiv32_fs207_xor1), .fs_or0(arrdiv32_fs207_or0));
  fs fs_arrdiv32_fs208_out(.a(arrdiv32_mux2to1170_xor0[0]), .b(b[16]), .bin(arrdiv32_fs207_or0[0]), .fs_xor1(arrdiv32_fs208_xor1), .fs_or0(arrdiv32_fs208_or0));
  fs fs_arrdiv32_fs209_out(.a(arrdiv32_mux2to1171_xor0[0]), .b(b[17]), .bin(arrdiv32_fs208_or0[0]), .fs_xor1(arrdiv32_fs209_xor1), .fs_or0(arrdiv32_fs209_or0));
  fs fs_arrdiv32_fs210_out(.a(arrdiv32_mux2to1172_xor0[0]), .b(b[18]), .bin(arrdiv32_fs209_or0[0]), .fs_xor1(arrdiv32_fs210_xor1), .fs_or0(arrdiv32_fs210_or0));
  fs fs_arrdiv32_fs211_out(.a(arrdiv32_mux2to1173_xor0[0]), .b(b[19]), .bin(arrdiv32_fs210_or0[0]), .fs_xor1(arrdiv32_fs211_xor1), .fs_or0(arrdiv32_fs211_or0));
  fs fs_arrdiv32_fs212_out(.a(arrdiv32_mux2to1174_xor0[0]), .b(b[20]), .bin(arrdiv32_fs211_or0[0]), .fs_xor1(arrdiv32_fs212_xor1), .fs_or0(arrdiv32_fs212_or0));
  fs fs_arrdiv32_fs213_out(.a(arrdiv32_mux2to1175_xor0[0]), .b(b[21]), .bin(arrdiv32_fs212_or0[0]), .fs_xor1(arrdiv32_fs213_xor1), .fs_or0(arrdiv32_fs213_or0));
  fs fs_arrdiv32_fs214_out(.a(arrdiv32_mux2to1176_xor0[0]), .b(b[22]), .bin(arrdiv32_fs213_or0[0]), .fs_xor1(arrdiv32_fs214_xor1), .fs_or0(arrdiv32_fs214_or0));
  fs fs_arrdiv32_fs215_out(.a(arrdiv32_mux2to1177_xor0[0]), .b(b[23]), .bin(arrdiv32_fs214_or0[0]), .fs_xor1(arrdiv32_fs215_xor1), .fs_or0(arrdiv32_fs215_or0));
  fs fs_arrdiv32_fs216_out(.a(arrdiv32_mux2to1178_xor0[0]), .b(b[24]), .bin(arrdiv32_fs215_or0[0]), .fs_xor1(arrdiv32_fs216_xor1), .fs_or0(arrdiv32_fs216_or0));
  fs fs_arrdiv32_fs217_out(.a(arrdiv32_mux2to1179_xor0[0]), .b(b[25]), .bin(arrdiv32_fs216_or0[0]), .fs_xor1(arrdiv32_fs217_xor1), .fs_or0(arrdiv32_fs217_or0));
  fs fs_arrdiv32_fs218_out(.a(arrdiv32_mux2to1180_xor0[0]), .b(b[26]), .bin(arrdiv32_fs217_or0[0]), .fs_xor1(arrdiv32_fs218_xor1), .fs_or0(arrdiv32_fs218_or0));
  fs fs_arrdiv32_fs219_out(.a(arrdiv32_mux2to1181_xor0[0]), .b(b[27]), .bin(arrdiv32_fs218_or0[0]), .fs_xor1(arrdiv32_fs219_xor1), .fs_or0(arrdiv32_fs219_or0));
  fs fs_arrdiv32_fs220_out(.a(arrdiv32_mux2to1182_xor0[0]), .b(b[28]), .bin(arrdiv32_fs219_or0[0]), .fs_xor1(arrdiv32_fs220_xor1), .fs_or0(arrdiv32_fs220_or0));
  fs fs_arrdiv32_fs221_out(.a(arrdiv32_mux2to1183_xor0[0]), .b(b[29]), .bin(arrdiv32_fs220_or0[0]), .fs_xor1(arrdiv32_fs221_xor1), .fs_or0(arrdiv32_fs221_or0));
  fs fs_arrdiv32_fs222_out(.a(arrdiv32_mux2to1184_xor0[0]), .b(b[30]), .bin(arrdiv32_fs221_or0[0]), .fs_xor1(arrdiv32_fs222_xor1), .fs_or0(arrdiv32_fs222_or0));
  fs fs_arrdiv32_fs223_out(.a(arrdiv32_mux2to1185_xor0[0]), .b(b[31]), .bin(arrdiv32_fs222_or0[0]), .fs_xor1(arrdiv32_fs223_xor1), .fs_or0(arrdiv32_fs223_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1186_out(.d0(arrdiv32_fs192_xor0[0]), .d1(a[25]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1186_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1187_out(.d0(arrdiv32_fs193_xor1[0]), .d1(arrdiv32_mux2to1155_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1187_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1188_out(.d0(arrdiv32_fs194_xor1[0]), .d1(arrdiv32_mux2to1156_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1188_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1189_out(.d0(arrdiv32_fs195_xor1[0]), .d1(arrdiv32_mux2to1157_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1189_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1190_out(.d0(arrdiv32_fs196_xor1[0]), .d1(arrdiv32_mux2to1158_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1190_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1191_out(.d0(arrdiv32_fs197_xor1[0]), .d1(arrdiv32_mux2to1159_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1191_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1192_out(.d0(arrdiv32_fs198_xor1[0]), .d1(arrdiv32_mux2to1160_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1192_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1193_out(.d0(arrdiv32_fs199_xor1[0]), .d1(arrdiv32_mux2to1161_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1193_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1194_out(.d0(arrdiv32_fs200_xor1[0]), .d1(arrdiv32_mux2to1162_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1194_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1195_out(.d0(arrdiv32_fs201_xor1[0]), .d1(arrdiv32_mux2to1163_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1195_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1196_out(.d0(arrdiv32_fs202_xor1[0]), .d1(arrdiv32_mux2to1164_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1196_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1197_out(.d0(arrdiv32_fs203_xor1[0]), .d1(arrdiv32_mux2to1165_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1197_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1198_out(.d0(arrdiv32_fs204_xor1[0]), .d1(arrdiv32_mux2to1166_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1198_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1199_out(.d0(arrdiv32_fs205_xor1[0]), .d1(arrdiv32_mux2to1167_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1199_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1200_out(.d0(arrdiv32_fs206_xor1[0]), .d1(arrdiv32_mux2to1168_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1200_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1201_out(.d0(arrdiv32_fs207_xor1[0]), .d1(arrdiv32_mux2to1169_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1201_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1202_out(.d0(arrdiv32_fs208_xor1[0]), .d1(arrdiv32_mux2to1170_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1202_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1203_out(.d0(arrdiv32_fs209_xor1[0]), .d1(arrdiv32_mux2to1171_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1203_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1204_out(.d0(arrdiv32_fs210_xor1[0]), .d1(arrdiv32_mux2to1172_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1204_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1205_out(.d0(arrdiv32_fs211_xor1[0]), .d1(arrdiv32_mux2to1173_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1205_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1206_out(.d0(arrdiv32_fs212_xor1[0]), .d1(arrdiv32_mux2to1174_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1206_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1207_out(.d0(arrdiv32_fs213_xor1[0]), .d1(arrdiv32_mux2to1175_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1207_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1208_out(.d0(arrdiv32_fs214_xor1[0]), .d1(arrdiv32_mux2to1176_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1208_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1209_out(.d0(arrdiv32_fs215_xor1[0]), .d1(arrdiv32_mux2to1177_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1209_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1210_out(.d0(arrdiv32_fs216_xor1[0]), .d1(arrdiv32_mux2to1178_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1210_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1211_out(.d0(arrdiv32_fs217_xor1[0]), .d1(arrdiv32_mux2to1179_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1211_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1212_out(.d0(arrdiv32_fs218_xor1[0]), .d1(arrdiv32_mux2to1180_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1212_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1213_out(.d0(arrdiv32_fs219_xor1[0]), .d1(arrdiv32_mux2to1181_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1213_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1214_out(.d0(arrdiv32_fs220_xor1[0]), .d1(arrdiv32_mux2to1182_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1214_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1215_out(.d0(arrdiv32_fs221_xor1[0]), .d1(arrdiv32_mux2to1183_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1215_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1216_out(.d0(arrdiv32_fs222_xor1[0]), .d1(arrdiv32_mux2to1184_xor0[0]), .sel(arrdiv32_fs223_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1216_xor0));
  not_gate not_gate_arrdiv32_not6(.a(arrdiv32_fs223_or0[0]), .out(arrdiv32_not6));
  fs fs_arrdiv32_fs224_out(.a(a[24]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs224_xor0), .fs_or0(arrdiv32_fs224_and0));
  fs fs_arrdiv32_fs225_out(.a(arrdiv32_mux2to1186_xor0[0]), .b(b[1]), .bin(arrdiv32_fs224_and0[0]), .fs_xor1(arrdiv32_fs225_xor1), .fs_or0(arrdiv32_fs225_or0));
  fs fs_arrdiv32_fs226_out(.a(arrdiv32_mux2to1187_xor0[0]), .b(b[2]), .bin(arrdiv32_fs225_or0[0]), .fs_xor1(arrdiv32_fs226_xor1), .fs_or0(arrdiv32_fs226_or0));
  fs fs_arrdiv32_fs227_out(.a(arrdiv32_mux2to1188_xor0[0]), .b(b[3]), .bin(arrdiv32_fs226_or0[0]), .fs_xor1(arrdiv32_fs227_xor1), .fs_or0(arrdiv32_fs227_or0));
  fs fs_arrdiv32_fs228_out(.a(arrdiv32_mux2to1189_xor0[0]), .b(b[4]), .bin(arrdiv32_fs227_or0[0]), .fs_xor1(arrdiv32_fs228_xor1), .fs_or0(arrdiv32_fs228_or0));
  fs fs_arrdiv32_fs229_out(.a(arrdiv32_mux2to1190_xor0[0]), .b(b[5]), .bin(arrdiv32_fs228_or0[0]), .fs_xor1(arrdiv32_fs229_xor1), .fs_or0(arrdiv32_fs229_or0));
  fs fs_arrdiv32_fs230_out(.a(arrdiv32_mux2to1191_xor0[0]), .b(b[6]), .bin(arrdiv32_fs229_or0[0]), .fs_xor1(arrdiv32_fs230_xor1), .fs_or0(arrdiv32_fs230_or0));
  fs fs_arrdiv32_fs231_out(.a(arrdiv32_mux2to1192_xor0[0]), .b(b[7]), .bin(arrdiv32_fs230_or0[0]), .fs_xor1(arrdiv32_fs231_xor1), .fs_or0(arrdiv32_fs231_or0));
  fs fs_arrdiv32_fs232_out(.a(arrdiv32_mux2to1193_xor0[0]), .b(b[8]), .bin(arrdiv32_fs231_or0[0]), .fs_xor1(arrdiv32_fs232_xor1), .fs_or0(arrdiv32_fs232_or0));
  fs fs_arrdiv32_fs233_out(.a(arrdiv32_mux2to1194_xor0[0]), .b(b[9]), .bin(arrdiv32_fs232_or0[0]), .fs_xor1(arrdiv32_fs233_xor1), .fs_or0(arrdiv32_fs233_or0));
  fs fs_arrdiv32_fs234_out(.a(arrdiv32_mux2to1195_xor0[0]), .b(b[10]), .bin(arrdiv32_fs233_or0[0]), .fs_xor1(arrdiv32_fs234_xor1), .fs_or0(arrdiv32_fs234_or0));
  fs fs_arrdiv32_fs235_out(.a(arrdiv32_mux2to1196_xor0[0]), .b(b[11]), .bin(arrdiv32_fs234_or0[0]), .fs_xor1(arrdiv32_fs235_xor1), .fs_or0(arrdiv32_fs235_or0));
  fs fs_arrdiv32_fs236_out(.a(arrdiv32_mux2to1197_xor0[0]), .b(b[12]), .bin(arrdiv32_fs235_or0[0]), .fs_xor1(arrdiv32_fs236_xor1), .fs_or0(arrdiv32_fs236_or0));
  fs fs_arrdiv32_fs237_out(.a(arrdiv32_mux2to1198_xor0[0]), .b(b[13]), .bin(arrdiv32_fs236_or0[0]), .fs_xor1(arrdiv32_fs237_xor1), .fs_or0(arrdiv32_fs237_or0));
  fs fs_arrdiv32_fs238_out(.a(arrdiv32_mux2to1199_xor0[0]), .b(b[14]), .bin(arrdiv32_fs237_or0[0]), .fs_xor1(arrdiv32_fs238_xor1), .fs_or0(arrdiv32_fs238_or0));
  fs fs_arrdiv32_fs239_out(.a(arrdiv32_mux2to1200_xor0[0]), .b(b[15]), .bin(arrdiv32_fs238_or0[0]), .fs_xor1(arrdiv32_fs239_xor1), .fs_or0(arrdiv32_fs239_or0));
  fs fs_arrdiv32_fs240_out(.a(arrdiv32_mux2to1201_xor0[0]), .b(b[16]), .bin(arrdiv32_fs239_or0[0]), .fs_xor1(arrdiv32_fs240_xor1), .fs_or0(arrdiv32_fs240_or0));
  fs fs_arrdiv32_fs241_out(.a(arrdiv32_mux2to1202_xor0[0]), .b(b[17]), .bin(arrdiv32_fs240_or0[0]), .fs_xor1(arrdiv32_fs241_xor1), .fs_or0(arrdiv32_fs241_or0));
  fs fs_arrdiv32_fs242_out(.a(arrdiv32_mux2to1203_xor0[0]), .b(b[18]), .bin(arrdiv32_fs241_or0[0]), .fs_xor1(arrdiv32_fs242_xor1), .fs_or0(arrdiv32_fs242_or0));
  fs fs_arrdiv32_fs243_out(.a(arrdiv32_mux2to1204_xor0[0]), .b(b[19]), .bin(arrdiv32_fs242_or0[0]), .fs_xor1(arrdiv32_fs243_xor1), .fs_or0(arrdiv32_fs243_or0));
  fs fs_arrdiv32_fs244_out(.a(arrdiv32_mux2to1205_xor0[0]), .b(b[20]), .bin(arrdiv32_fs243_or0[0]), .fs_xor1(arrdiv32_fs244_xor1), .fs_or0(arrdiv32_fs244_or0));
  fs fs_arrdiv32_fs245_out(.a(arrdiv32_mux2to1206_xor0[0]), .b(b[21]), .bin(arrdiv32_fs244_or0[0]), .fs_xor1(arrdiv32_fs245_xor1), .fs_or0(arrdiv32_fs245_or0));
  fs fs_arrdiv32_fs246_out(.a(arrdiv32_mux2to1207_xor0[0]), .b(b[22]), .bin(arrdiv32_fs245_or0[0]), .fs_xor1(arrdiv32_fs246_xor1), .fs_or0(arrdiv32_fs246_or0));
  fs fs_arrdiv32_fs247_out(.a(arrdiv32_mux2to1208_xor0[0]), .b(b[23]), .bin(arrdiv32_fs246_or0[0]), .fs_xor1(arrdiv32_fs247_xor1), .fs_or0(arrdiv32_fs247_or0));
  fs fs_arrdiv32_fs248_out(.a(arrdiv32_mux2to1209_xor0[0]), .b(b[24]), .bin(arrdiv32_fs247_or0[0]), .fs_xor1(arrdiv32_fs248_xor1), .fs_or0(arrdiv32_fs248_or0));
  fs fs_arrdiv32_fs249_out(.a(arrdiv32_mux2to1210_xor0[0]), .b(b[25]), .bin(arrdiv32_fs248_or0[0]), .fs_xor1(arrdiv32_fs249_xor1), .fs_or0(arrdiv32_fs249_or0));
  fs fs_arrdiv32_fs250_out(.a(arrdiv32_mux2to1211_xor0[0]), .b(b[26]), .bin(arrdiv32_fs249_or0[0]), .fs_xor1(arrdiv32_fs250_xor1), .fs_or0(arrdiv32_fs250_or0));
  fs fs_arrdiv32_fs251_out(.a(arrdiv32_mux2to1212_xor0[0]), .b(b[27]), .bin(arrdiv32_fs250_or0[0]), .fs_xor1(arrdiv32_fs251_xor1), .fs_or0(arrdiv32_fs251_or0));
  fs fs_arrdiv32_fs252_out(.a(arrdiv32_mux2to1213_xor0[0]), .b(b[28]), .bin(arrdiv32_fs251_or0[0]), .fs_xor1(arrdiv32_fs252_xor1), .fs_or0(arrdiv32_fs252_or0));
  fs fs_arrdiv32_fs253_out(.a(arrdiv32_mux2to1214_xor0[0]), .b(b[29]), .bin(arrdiv32_fs252_or0[0]), .fs_xor1(arrdiv32_fs253_xor1), .fs_or0(arrdiv32_fs253_or0));
  fs fs_arrdiv32_fs254_out(.a(arrdiv32_mux2to1215_xor0[0]), .b(b[30]), .bin(arrdiv32_fs253_or0[0]), .fs_xor1(arrdiv32_fs254_xor1), .fs_or0(arrdiv32_fs254_or0));
  fs fs_arrdiv32_fs255_out(.a(arrdiv32_mux2to1216_xor0[0]), .b(b[31]), .bin(arrdiv32_fs254_or0[0]), .fs_xor1(arrdiv32_fs255_xor1), .fs_or0(arrdiv32_fs255_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1217_out(.d0(arrdiv32_fs224_xor0[0]), .d1(a[24]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1217_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1218_out(.d0(arrdiv32_fs225_xor1[0]), .d1(arrdiv32_mux2to1186_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1218_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1219_out(.d0(arrdiv32_fs226_xor1[0]), .d1(arrdiv32_mux2to1187_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1219_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1220_out(.d0(arrdiv32_fs227_xor1[0]), .d1(arrdiv32_mux2to1188_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1220_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1221_out(.d0(arrdiv32_fs228_xor1[0]), .d1(arrdiv32_mux2to1189_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1221_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1222_out(.d0(arrdiv32_fs229_xor1[0]), .d1(arrdiv32_mux2to1190_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1222_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1223_out(.d0(arrdiv32_fs230_xor1[0]), .d1(arrdiv32_mux2to1191_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1223_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1224_out(.d0(arrdiv32_fs231_xor1[0]), .d1(arrdiv32_mux2to1192_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1224_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1225_out(.d0(arrdiv32_fs232_xor1[0]), .d1(arrdiv32_mux2to1193_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1225_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1226_out(.d0(arrdiv32_fs233_xor1[0]), .d1(arrdiv32_mux2to1194_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1226_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1227_out(.d0(arrdiv32_fs234_xor1[0]), .d1(arrdiv32_mux2to1195_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1227_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1228_out(.d0(arrdiv32_fs235_xor1[0]), .d1(arrdiv32_mux2to1196_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1228_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1229_out(.d0(arrdiv32_fs236_xor1[0]), .d1(arrdiv32_mux2to1197_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1229_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1230_out(.d0(arrdiv32_fs237_xor1[0]), .d1(arrdiv32_mux2to1198_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1230_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1231_out(.d0(arrdiv32_fs238_xor1[0]), .d1(arrdiv32_mux2to1199_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1231_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1232_out(.d0(arrdiv32_fs239_xor1[0]), .d1(arrdiv32_mux2to1200_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1232_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1233_out(.d0(arrdiv32_fs240_xor1[0]), .d1(arrdiv32_mux2to1201_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1233_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1234_out(.d0(arrdiv32_fs241_xor1[0]), .d1(arrdiv32_mux2to1202_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1234_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1235_out(.d0(arrdiv32_fs242_xor1[0]), .d1(arrdiv32_mux2to1203_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1235_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1236_out(.d0(arrdiv32_fs243_xor1[0]), .d1(arrdiv32_mux2to1204_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1236_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1237_out(.d0(arrdiv32_fs244_xor1[0]), .d1(arrdiv32_mux2to1205_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1237_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1238_out(.d0(arrdiv32_fs245_xor1[0]), .d1(arrdiv32_mux2to1206_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1238_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1239_out(.d0(arrdiv32_fs246_xor1[0]), .d1(arrdiv32_mux2to1207_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1239_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1240_out(.d0(arrdiv32_fs247_xor1[0]), .d1(arrdiv32_mux2to1208_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1240_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1241_out(.d0(arrdiv32_fs248_xor1[0]), .d1(arrdiv32_mux2to1209_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1241_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1242_out(.d0(arrdiv32_fs249_xor1[0]), .d1(arrdiv32_mux2to1210_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1242_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1243_out(.d0(arrdiv32_fs250_xor1[0]), .d1(arrdiv32_mux2to1211_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1243_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1244_out(.d0(arrdiv32_fs251_xor1[0]), .d1(arrdiv32_mux2to1212_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1244_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1245_out(.d0(arrdiv32_fs252_xor1[0]), .d1(arrdiv32_mux2to1213_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1245_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1246_out(.d0(arrdiv32_fs253_xor1[0]), .d1(arrdiv32_mux2to1214_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1246_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1247_out(.d0(arrdiv32_fs254_xor1[0]), .d1(arrdiv32_mux2to1215_xor0[0]), .sel(arrdiv32_fs255_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1247_xor0));
  not_gate not_gate_arrdiv32_not7(.a(arrdiv32_fs255_or0[0]), .out(arrdiv32_not7));
  fs fs_arrdiv32_fs256_out(.a(a[23]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs256_xor0), .fs_or0(arrdiv32_fs256_and0));
  fs fs_arrdiv32_fs257_out(.a(arrdiv32_mux2to1217_xor0[0]), .b(b[1]), .bin(arrdiv32_fs256_and0[0]), .fs_xor1(arrdiv32_fs257_xor1), .fs_or0(arrdiv32_fs257_or0));
  fs fs_arrdiv32_fs258_out(.a(arrdiv32_mux2to1218_xor0[0]), .b(b[2]), .bin(arrdiv32_fs257_or0[0]), .fs_xor1(arrdiv32_fs258_xor1), .fs_or0(arrdiv32_fs258_or0));
  fs fs_arrdiv32_fs259_out(.a(arrdiv32_mux2to1219_xor0[0]), .b(b[3]), .bin(arrdiv32_fs258_or0[0]), .fs_xor1(arrdiv32_fs259_xor1), .fs_or0(arrdiv32_fs259_or0));
  fs fs_arrdiv32_fs260_out(.a(arrdiv32_mux2to1220_xor0[0]), .b(b[4]), .bin(arrdiv32_fs259_or0[0]), .fs_xor1(arrdiv32_fs260_xor1), .fs_or0(arrdiv32_fs260_or0));
  fs fs_arrdiv32_fs261_out(.a(arrdiv32_mux2to1221_xor0[0]), .b(b[5]), .bin(arrdiv32_fs260_or0[0]), .fs_xor1(arrdiv32_fs261_xor1), .fs_or0(arrdiv32_fs261_or0));
  fs fs_arrdiv32_fs262_out(.a(arrdiv32_mux2to1222_xor0[0]), .b(b[6]), .bin(arrdiv32_fs261_or0[0]), .fs_xor1(arrdiv32_fs262_xor1), .fs_or0(arrdiv32_fs262_or0));
  fs fs_arrdiv32_fs263_out(.a(arrdiv32_mux2to1223_xor0[0]), .b(b[7]), .bin(arrdiv32_fs262_or0[0]), .fs_xor1(arrdiv32_fs263_xor1), .fs_or0(arrdiv32_fs263_or0));
  fs fs_arrdiv32_fs264_out(.a(arrdiv32_mux2to1224_xor0[0]), .b(b[8]), .bin(arrdiv32_fs263_or0[0]), .fs_xor1(arrdiv32_fs264_xor1), .fs_or0(arrdiv32_fs264_or0));
  fs fs_arrdiv32_fs265_out(.a(arrdiv32_mux2to1225_xor0[0]), .b(b[9]), .bin(arrdiv32_fs264_or0[0]), .fs_xor1(arrdiv32_fs265_xor1), .fs_or0(arrdiv32_fs265_or0));
  fs fs_arrdiv32_fs266_out(.a(arrdiv32_mux2to1226_xor0[0]), .b(b[10]), .bin(arrdiv32_fs265_or0[0]), .fs_xor1(arrdiv32_fs266_xor1), .fs_or0(arrdiv32_fs266_or0));
  fs fs_arrdiv32_fs267_out(.a(arrdiv32_mux2to1227_xor0[0]), .b(b[11]), .bin(arrdiv32_fs266_or0[0]), .fs_xor1(arrdiv32_fs267_xor1), .fs_or0(arrdiv32_fs267_or0));
  fs fs_arrdiv32_fs268_out(.a(arrdiv32_mux2to1228_xor0[0]), .b(b[12]), .bin(arrdiv32_fs267_or0[0]), .fs_xor1(arrdiv32_fs268_xor1), .fs_or0(arrdiv32_fs268_or0));
  fs fs_arrdiv32_fs269_out(.a(arrdiv32_mux2to1229_xor0[0]), .b(b[13]), .bin(arrdiv32_fs268_or0[0]), .fs_xor1(arrdiv32_fs269_xor1), .fs_or0(arrdiv32_fs269_or0));
  fs fs_arrdiv32_fs270_out(.a(arrdiv32_mux2to1230_xor0[0]), .b(b[14]), .bin(arrdiv32_fs269_or0[0]), .fs_xor1(arrdiv32_fs270_xor1), .fs_or0(arrdiv32_fs270_or0));
  fs fs_arrdiv32_fs271_out(.a(arrdiv32_mux2to1231_xor0[0]), .b(b[15]), .bin(arrdiv32_fs270_or0[0]), .fs_xor1(arrdiv32_fs271_xor1), .fs_or0(arrdiv32_fs271_or0));
  fs fs_arrdiv32_fs272_out(.a(arrdiv32_mux2to1232_xor0[0]), .b(b[16]), .bin(arrdiv32_fs271_or0[0]), .fs_xor1(arrdiv32_fs272_xor1), .fs_or0(arrdiv32_fs272_or0));
  fs fs_arrdiv32_fs273_out(.a(arrdiv32_mux2to1233_xor0[0]), .b(b[17]), .bin(arrdiv32_fs272_or0[0]), .fs_xor1(arrdiv32_fs273_xor1), .fs_or0(arrdiv32_fs273_or0));
  fs fs_arrdiv32_fs274_out(.a(arrdiv32_mux2to1234_xor0[0]), .b(b[18]), .bin(arrdiv32_fs273_or0[0]), .fs_xor1(arrdiv32_fs274_xor1), .fs_or0(arrdiv32_fs274_or0));
  fs fs_arrdiv32_fs275_out(.a(arrdiv32_mux2to1235_xor0[0]), .b(b[19]), .bin(arrdiv32_fs274_or0[0]), .fs_xor1(arrdiv32_fs275_xor1), .fs_or0(arrdiv32_fs275_or0));
  fs fs_arrdiv32_fs276_out(.a(arrdiv32_mux2to1236_xor0[0]), .b(b[20]), .bin(arrdiv32_fs275_or0[0]), .fs_xor1(arrdiv32_fs276_xor1), .fs_or0(arrdiv32_fs276_or0));
  fs fs_arrdiv32_fs277_out(.a(arrdiv32_mux2to1237_xor0[0]), .b(b[21]), .bin(arrdiv32_fs276_or0[0]), .fs_xor1(arrdiv32_fs277_xor1), .fs_or0(arrdiv32_fs277_or0));
  fs fs_arrdiv32_fs278_out(.a(arrdiv32_mux2to1238_xor0[0]), .b(b[22]), .bin(arrdiv32_fs277_or0[0]), .fs_xor1(arrdiv32_fs278_xor1), .fs_or0(arrdiv32_fs278_or0));
  fs fs_arrdiv32_fs279_out(.a(arrdiv32_mux2to1239_xor0[0]), .b(b[23]), .bin(arrdiv32_fs278_or0[0]), .fs_xor1(arrdiv32_fs279_xor1), .fs_or0(arrdiv32_fs279_or0));
  fs fs_arrdiv32_fs280_out(.a(arrdiv32_mux2to1240_xor0[0]), .b(b[24]), .bin(arrdiv32_fs279_or0[0]), .fs_xor1(arrdiv32_fs280_xor1), .fs_or0(arrdiv32_fs280_or0));
  fs fs_arrdiv32_fs281_out(.a(arrdiv32_mux2to1241_xor0[0]), .b(b[25]), .bin(arrdiv32_fs280_or0[0]), .fs_xor1(arrdiv32_fs281_xor1), .fs_or0(arrdiv32_fs281_or0));
  fs fs_arrdiv32_fs282_out(.a(arrdiv32_mux2to1242_xor0[0]), .b(b[26]), .bin(arrdiv32_fs281_or0[0]), .fs_xor1(arrdiv32_fs282_xor1), .fs_or0(arrdiv32_fs282_or0));
  fs fs_arrdiv32_fs283_out(.a(arrdiv32_mux2to1243_xor0[0]), .b(b[27]), .bin(arrdiv32_fs282_or0[0]), .fs_xor1(arrdiv32_fs283_xor1), .fs_or0(arrdiv32_fs283_or0));
  fs fs_arrdiv32_fs284_out(.a(arrdiv32_mux2to1244_xor0[0]), .b(b[28]), .bin(arrdiv32_fs283_or0[0]), .fs_xor1(arrdiv32_fs284_xor1), .fs_or0(arrdiv32_fs284_or0));
  fs fs_arrdiv32_fs285_out(.a(arrdiv32_mux2to1245_xor0[0]), .b(b[29]), .bin(arrdiv32_fs284_or0[0]), .fs_xor1(arrdiv32_fs285_xor1), .fs_or0(arrdiv32_fs285_or0));
  fs fs_arrdiv32_fs286_out(.a(arrdiv32_mux2to1246_xor0[0]), .b(b[30]), .bin(arrdiv32_fs285_or0[0]), .fs_xor1(arrdiv32_fs286_xor1), .fs_or0(arrdiv32_fs286_or0));
  fs fs_arrdiv32_fs287_out(.a(arrdiv32_mux2to1247_xor0[0]), .b(b[31]), .bin(arrdiv32_fs286_or0[0]), .fs_xor1(arrdiv32_fs287_xor1), .fs_or0(arrdiv32_fs287_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1248_out(.d0(arrdiv32_fs256_xor0[0]), .d1(a[23]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1248_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1249_out(.d0(arrdiv32_fs257_xor1[0]), .d1(arrdiv32_mux2to1217_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1249_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1250_out(.d0(arrdiv32_fs258_xor1[0]), .d1(arrdiv32_mux2to1218_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1250_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1251_out(.d0(arrdiv32_fs259_xor1[0]), .d1(arrdiv32_mux2to1219_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1251_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1252_out(.d0(arrdiv32_fs260_xor1[0]), .d1(arrdiv32_mux2to1220_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1252_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1253_out(.d0(arrdiv32_fs261_xor1[0]), .d1(arrdiv32_mux2to1221_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1253_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1254_out(.d0(arrdiv32_fs262_xor1[0]), .d1(arrdiv32_mux2to1222_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1254_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1255_out(.d0(arrdiv32_fs263_xor1[0]), .d1(arrdiv32_mux2to1223_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1255_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1256_out(.d0(arrdiv32_fs264_xor1[0]), .d1(arrdiv32_mux2to1224_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1256_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1257_out(.d0(arrdiv32_fs265_xor1[0]), .d1(arrdiv32_mux2to1225_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1257_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1258_out(.d0(arrdiv32_fs266_xor1[0]), .d1(arrdiv32_mux2to1226_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1258_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1259_out(.d0(arrdiv32_fs267_xor1[0]), .d1(arrdiv32_mux2to1227_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1259_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1260_out(.d0(arrdiv32_fs268_xor1[0]), .d1(arrdiv32_mux2to1228_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1260_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1261_out(.d0(arrdiv32_fs269_xor1[0]), .d1(arrdiv32_mux2to1229_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1261_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1262_out(.d0(arrdiv32_fs270_xor1[0]), .d1(arrdiv32_mux2to1230_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1262_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1263_out(.d0(arrdiv32_fs271_xor1[0]), .d1(arrdiv32_mux2to1231_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1263_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1264_out(.d0(arrdiv32_fs272_xor1[0]), .d1(arrdiv32_mux2to1232_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1264_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1265_out(.d0(arrdiv32_fs273_xor1[0]), .d1(arrdiv32_mux2to1233_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1265_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1266_out(.d0(arrdiv32_fs274_xor1[0]), .d1(arrdiv32_mux2to1234_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1266_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1267_out(.d0(arrdiv32_fs275_xor1[0]), .d1(arrdiv32_mux2to1235_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1267_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1268_out(.d0(arrdiv32_fs276_xor1[0]), .d1(arrdiv32_mux2to1236_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1268_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1269_out(.d0(arrdiv32_fs277_xor1[0]), .d1(arrdiv32_mux2to1237_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1269_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1270_out(.d0(arrdiv32_fs278_xor1[0]), .d1(arrdiv32_mux2to1238_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1270_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1271_out(.d0(arrdiv32_fs279_xor1[0]), .d1(arrdiv32_mux2to1239_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1271_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1272_out(.d0(arrdiv32_fs280_xor1[0]), .d1(arrdiv32_mux2to1240_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1272_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1273_out(.d0(arrdiv32_fs281_xor1[0]), .d1(arrdiv32_mux2to1241_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1273_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1274_out(.d0(arrdiv32_fs282_xor1[0]), .d1(arrdiv32_mux2to1242_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1274_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1275_out(.d0(arrdiv32_fs283_xor1[0]), .d1(arrdiv32_mux2to1243_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1275_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1276_out(.d0(arrdiv32_fs284_xor1[0]), .d1(arrdiv32_mux2to1244_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1276_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1277_out(.d0(arrdiv32_fs285_xor1[0]), .d1(arrdiv32_mux2to1245_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1277_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1278_out(.d0(arrdiv32_fs286_xor1[0]), .d1(arrdiv32_mux2to1246_xor0[0]), .sel(arrdiv32_fs287_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1278_xor0));
  not_gate not_gate_arrdiv32_not8(.a(arrdiv32_fs287_or0[0]), .out(arrdiv32_not8));
  fs fs_arrdiv32_fs288_out(.a(a[22]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs288_xor0), .fs_or0(arrdiv32_fs288_and0));
  fs fs_arrdiv32_fs289_out(.a(arrdiv32_mux2to1248_xor0[0]), .b(b[1]), .bin(arrdiv32_fs288_and0[0]), .fs_xor1(arrdiv32_fs289_xor1), .fs_or0(arrdiv32_fs289_or0));
  fs fs_arrdiv32_fs290_out(.a(arrdiv32_mux2to1249_xor0[0]), .b(b[2]), .bin(arrdiv32_fs289_or0[0]), .fs_xor1(arrdiv32_fs290_xor1), .fs_or0(arrdiv32_fs290_or0));
  fs fs_arrdiv32_fs291_out(.a(arrdiv32_mux2to1250_xor0[0]), .b(b[3]), .bin(arrdiv32_fs290_or0[0]), .fs_xor1(arrdiv32_fs291_xor1), .fs_or0(arrdiv32_fs291_or0));
  fs fs_arrdiv32_fs292_out(.a(arrdiv32_mux2to1251_xor0[0]), .b(b[4]), .bin(arrdiv32_fs291_or0[0]), .fs_xor1(arrdiv32_fs292_xor1), .fs_or0(arrdiv32_fs292_or0));
  fs fs_arrdiv32_fs293_out(.a(arrdiv32_mux2to1252_xor0[0]), .b(b[5]), .bin(arrdiv32_fs292_or0[0]), .fs_xor1(arrdiv32_fs293_xor1), .fs_or0(arrdiv32_fs293_or0));
  fs fs_arrdiv32_fs294_out(.a(arrdiv32_mux2to1253_xor0[0]), .b(b[6]), .bin(arrdiv32_fs293_or0[0]), .fs_xor1(arrdiv32_fs294_xor1), .fs_or0(arrdiv32_fs294_or0));
  fs fs_arrdiv32_fs295_out(.a(arrdiv32_mux2to1254_xor0[0]), .b(b[7]), .bin(arrdiv32_fs294_or0[0]), .fs_xor1(arrdiv32_fs295_xor1), .fs_or0(arrdiv32_fs295_or0));
  fs fs_arrdiv32_fs296_out(.a(arrdiv32_mux2to1255_xor0[0]), .b(b[8]), .bin(arrdiv32_fs295_or0[0]), .fs_xor1(arrdiv32_fs296_xor1), .fs_or0(arrdiv32_fs296_or0));
  fs fs_arrdiv32_fs297_out(.a(arrdiv32_mux2to1256_xor0[0]), .b(b[9]), .bin(arrdiv32_fs296_or0[0]), .fs_xor1(arrdiv32_fs297_xor1), .fs_or0(arrdiv32_fs297_or0));
  fs fs_arrdiv32_fs298_out(.a(arrdiv32_mux2to1257_xor0[0]), .b(b[10]), .bin(arrdiv32_fs297_or0[0]), .fs_xor1(arrdiv32_fs298_xor1), .fs_or0(arrdiv32_fs298_or0));
  fs fs_arrdiv32_fs299_out(.a(arrdiv32_mux2to1258_xor0[0]), .b(b[11]), .bin(arrdiv32_fs298_or0[0]), .fs_xor1(arrdiv32_fs299_xor1), .fs_or0(arrdiv32_fs299_or0));
  fs fs_arrdiv32_fs300_out(.a(arrdiv32_mux2to1259_xor0[0]), .b(b[12]), .bin(arrdiv32_fs299_or0[0]), .fs_xor1(arrdiv32_fs300_xor1), .fs_or0(arrdiv32_fs300_or0));
  fs fs_arrdiv32_fs301_out(.a(arrdiv32_mux2to1260_xor0[0]), .b(b[13]), .bin(arrdiv32_fs300_or0[0]), .fs_xor1(arrdiv32_fs301_xor1), .fs_or0(arrdiv32_fs301_or0));
  fs fs_arrdiv32_fs302_out(.a(arrdiv32_mux2to1261_xor0[0]), .b(b[14]), .bin(arrdiv32_fs301_or0[0]), .fs_xor1(arrdiv32_fs302_xor1), .fs_or0(arrdiv32_fs302_or0));
  fs fs_arrdiv32_fs303_out(.a(arrdiv32_mux2to1262_xor0[0]), .b(b[15]), .bin(arrdiv32_fs302_or0[0]), .fs_xor1(arrdiv32_fs303_xor1), .fs_or0(arrdiv32_fs303_or0));
  fs fs_arrdiv32_fs304_out(.a(arrdiv32_mux2to1263_xor0[0]), .b(b[16]), .bin(arrdiv32_fs303_or0[0]), .fs_xor1(arrdiv32_fs304_xor1), .fs_or0(arrdiv32_fs304_or0));
  fs fs_arrdiv32_fs305_out(.a(arrdiv32_mux2to1264_xor0[0]), .b(b[17]), .bin(arrdiv32_fs304_or0[0]), .fs_xor1(arrdiv32_fs305_xor1), .fs_or0(arrdiv32_fs305_or0));
  fs fs_arrdiv32_fs306_out(.a(arrdiv32_mux2to1265_xor0[0]), .b(b[18]), .bin(arrdiv32_fs305_or0[0]), .fs_xor1(arrdiv32_fs306_xor1), .fs_or0(arrdiv32_fs306_or0));
  fs fs_arrdiv32_fs307_out(.a(arrdiv32_mux2to1266_xor0[0]), .b(b[19]), .bin(arrdiv32_fs306_or0[0]), .fs_xor1(arrdiv32_fs307_xor1), .fs_or0(arrdiv32_fs307_or0));
  fs fs_arrdiv32_fs308_out(.a(arrdiv32_mux2to1267_xor0[0]), .b(b[20]), .bin(arrdiv32_fs307_or0[0]), .fs_xor1(arrdiv32_fs308_xor1), .fs_or0(arrdiv32_fs308_or0));
  fs fs_arrdiv32_fs309_out(.a(arrdiv32_mux2to1268_xor0[0]), .b(b[21]), .bin(arrdiv32_fs308_or0[0]), .fs_xor1(arrdiv32_fs309_xor1), .fs_or0(arrdiv32_fs309_or0));
  fs fs_arrdiv32_fs310_out(.a(arrdiv32_mux2to1269_xor0[0]), .b(b[22]), .bin(arrdiv32_fs309_or0[0]), .fs_xor1(arrdiv32_fs310_xor1), .fs_or0(arrdiv32_fs310_or0));
  fs fs_arrdiv32_fs311_out(.a(arrdiv32_mux2to1270_xor0[0]), .b(b[23]), .bin(arrdiv32_fs310_or0[0]), .fs_xor1(arrdiv32_fs311_xor1), .fs_or0(arrdiv32_fs311_or0));
  fs fs_arrdiv32_fs312_out(.a(arrdiv32_mux2to1271_xor0[0]), .b(b[24]), .bin(arrdiv32_fs311_or0[0]), .fs_xor1(arrdiv32_fs312_xor1), .fs_or0(arrdiv32_fs312_or0));
  fs fs_arrdiv32_fs313_out(.a(arrdiv32_mux2to1272_xor0[0]), .b(b[25]), .bin(arrdiv32_fs312_or0[0]), .fs_xor1(arrdiv32_fs313_xor1), .fs_or0(arrdiv32_fs313_or0));
  fs fs_arrdiv32_fs314_out(.a(arrdiv32_mux2to1273_xor0[0]), .b(b[26]), .bin(arrdiv32_fs313_or0[0]), .fs_xor1(arrdiv32_fs314_xor1), .fs_or0(arrdiv32_fs314_or0));
  fs fs_arrdiv32_fs315_out(.a(arrdiv32_mux2to1274_xor0[0]), .b(b[27]), .bin(arrdiv32_fs314_or0[0]), .fs_xor1(arrdiv32_fs315_xor1), .fs_or0(arrdiv32_fs315_or0));
  fs fs_arrdiv32_fs316_out(.a(arrdiv32_mux2to1275_xor0[0]), .b(b[28]), .bin(arrdiv32_fs315_or0[0]), .fs_xor1(arrdiv32_fs316_xor1), .fs_or0(arrdiv32_fs316_or0));
  fs fs_arrdiv32_fs317_out(.a(arrdiv32_mux2to1276_xor0[0]), .b(b[29]), .bin(arrdiv32_fs316_or0[0]), .fs_xor1(arrdiv32_fs317_xor1), .fs_or0(arrdiv32_fs317_or0));
  fs fs_arrdiv32_fs318_out(.a(arrdiv32_mux2to1277_xor0[0]), .b(b[30]), .bin(arrdiv32_fs317_or0[0]), .fs_xor1(arrdiv32_fs318_xor1), .fs_or0(arrdiv32_fs318_or0));
  fs fs_arrdiv32_fs319_out(.a(arrdiv32_mux2to1278_xor0[0]), .b(b[31]), .bin(arrdiv32_fs318_or0[0]), .fs_xor1(arrdiv32_fs319_xor1), .fs_or0(arrdiv32_fs319_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1279_out(.d0(arrdiv32_fs288_xor0[0]), .d1(a[22]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1279_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1280_out(.d0(arrdiv32_fs289_xor1[0]), .d1(arrdiv32_mux2to1248_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1280_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1281_out(.d0(arrdiv32_fs290_xor1[0]), .d1(arrdiv32_mux2to1249_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1281_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1282_out(.d0(arrdiv32_fs291_xor1[0]), .d1(arrdiv32_mux2to1250_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1282_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1283_out(.d0(arrdiv32_fs292_xor1[0]), .d1(arrdiv32_mux2to1251_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1283_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1284_out(.d0(arrdiv32_fs293_xor1[0]), .d1(arrdiv32_mux2to1252_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1284_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1285_out(.d0(arrdiv32_fs294_xor1[0]), .d1(arrdiv32_mux2to1253_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1285_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1286_out(.d0(arrdiv32_fs295_xor1[0]), .d1(arrdiv32_mux2to1254_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1286_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1287_out(.d0(arrdiv32_fs296_xor1[0]), .d1(arrdiv32_mux2to1255_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1287_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1288_out(.d0(arrdiv32_fs297_xor1[0]), .d1(arrdiv32_mux2to1256_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1288_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1289_out(.d0(arrdiv32_fs298_xor1[0]), .d1(arrdiv32_mux2to1257_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1289_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1290_out(.d0(arrdiv32_fs299_xor1[0]), .d1(arrdiv32_mux2to1258_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1290_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1291_out(.d0(arrdiv32_fs300_xor1[0]), .d1(arrdiv32_mux2to1259_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1291_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1292_out(.d0(arrdiv32_fs301_xor1[0]), .d1(arrdiv32_mux2to1260_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1292_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1293_out(.d0(arrdiv32_fs302_xor1[0]), .d1(arrdiv32_mux2to1261_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1293_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1294_out(.d0(arrdiv32_fs303_xor1[0]), .d1(arrdiv32_mux2to1262_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1294_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1295_out(.d0(arrdiv32_fs304_xor1[0]), .d1(arrdiv32_mux2to1263_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1295_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1296_out(.d0(arrdiv32_fs305_xor1[0]), .d1(arrdiv32_mux2to1264_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1296_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1297_out(.d0(arrdiv32_fs306_xor1[0]), .d1(arrdiv32_mux2to1265_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1297_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1298_out(.d0(arrdiv32_fs307_xor1[0]), .d1(arrdiv32_mux2to1266_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1298_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1299_out(.d0(arrdiv32_fs308_xor1[0]), .d1(arrdiv32_mux2to1267_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1299_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1300_out(.d0(arrdiv32_fs309_xor1[0]), .d1(arrdiv32_mux2to1268_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1300_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1301_out(.d0(arrdiv32_fs310_xor1[0]), .d1(arrdiv32_mux2to1269_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1301_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1302_out(.d0(arrdiv32_fs311_xor1[0]), .d1(arrdiv32_mux2to1270_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1302_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1303_out(.d0(arrdiv32_fs312_xor1[0]), .d1(arrdiv32_mux2to1271_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1303_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1304_out(.d0(arrdiv32_fs313_xor1[0]), .d1(arrdiv32_mux2to1272_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1304_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1305_out(.d0(arrdiv32_fs314_xor1[0]), .d1(arrdiv32_mux2to1273_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1305_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1306_out(.d0(arrdiv32_fs315_xor1[0]), .d1(arrdiv32_mux2to1274_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1306_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1307_out(.d0(arrdiv32_fs316_xor1[0]), .d1(arrdiv32_mux2to1275_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1307_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1308_out(.d0(arrdiv32_fs317_xor1[0]), .d1(arrdiv32_mux2to1276_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1308_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1309_out(.d0(arrdiv32_fs318_xor1[0]), .d1(arrdiv32_mux2to1277_xor0[0]), .sel(arrdiv32_fs319_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1309_xor0));
  not_gate not_gate_arrdiv32_not9(.a(arrdiv32_fs319_or0[0]), .out(arrdiv32_not9));
  fs fs_arrdiv32_fs320_out(.a(a[21]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs320_xor0), .fs_or0(arrdiv32_fs320_and0));
  fs fs_arrdiv32_fs321_out(.a(arrdiv32_mux2to1279_xor0[0]), .b(b[1]), .bin(arrdiv32_fs320_and0[0]), .fs_xor1(arrdiv32_fs321_xor1), .fs_or0(arrdiv32_fs321_or0));
  fs fs_arrdiv32_fs322_out(.a(arrdiv32_mux2to1280_xor0[0]), .b(b[2]), .bin(arrdiv32_fs321_or0[0]), .fs_xor1(arrdiv32_fs322_xor1), .fs_or0(arrdiv32_fs322_or0));
  fs fs_arrdiv32_fs323_out(.a(arrdiv32_mux2to1281_xor0[0]), .b(b[3]), .bin(arrdiv32_fs322_or0[0]), .fs_xor1(arrdiv32_fs323_xor1), .fs_or0(arrdiv32_fs323_or0));
  fs fs_arrdiv32_fs324_out(.a(arrdiv32_mux2to1282_xor0[0]), .b(b[4]), .bin(arrdiv32_fs323_or0[0]), .fs_xor1(arrdiv32_fs324_xor1), .fs_or0(arrdiv32_fs324_or0));
  fs fs_arrdiv32_fs325_out(.a(arrdiv32_mux2to1283_xor0[0]), .b(b[5]), .bin(arrdiv32_fs324_or0[0]), .fs_xor1(arrdiv32_fs325_xor1), .fs_or0(arrdiv32_fs325_or0));
  fs fs_arrdiv32_fs326_out(.a(arrdiv32_mux2to1284_xor0[0]), .b(b[6]), .bin(arrdiv32_fs325_or0[0]), .fs_xor1(arrdiv32_fs326_xor1), .fs_or0(arrdiv32_fs326_or0));
  fs fs_arrdiv32_fs327_out(.a(arrdiv32_mux2to1285_xor0[0]), .b(b[7]), .bin(arrdiv32_fs326_or0[0]), .fs_xor1(arrdiv32_fs327_xor1), .fs_or0(arrdiv32_fs327_or0));
  fs fs_arrdiv32_fs328_out(.a(arrdiv32_mux2to1286_xor0[0]), .b(b[8]), .bin(arrdiv32_fs327_or0[0]), .fs_xor1(arrdiv32_fs328_xor1), .fs_or0(arrdiv32_fs328_or0));
  fs fs_arrdiv32_fs329_out(.a(arrdiv32_mux2to1287_xor0[0]), .b(b[9]), .bin(arrdiv32_fs328_or0[0]), .fs_xor1(arrdiv32_fs329_xor1), .fs_or0(arrdiv32_fs329_or0));
  fs fs_arrdiv32_fs330_out(.a(arrdiv32_mux2to1288_xor0[0]), .b(b[10]), .bin(arrdiv32_fs329_or0[0]), .fs_xor1(arrdiv32_fs330_xor1), .fs_or0(arrdiv32_fs330_or0));
  fs fs_arrdiv32_fs331_out(.a(arrdiv32_mux2to1289_xor0[0]), .b(b[11]), .bin(arrdiv32_fs330_or0[0]), .fs_xor1(arrdiv32_fs331_xor1), .fs_or0(arrdiv32_fs331_or0));
  fs fs_arrdiv32_fs332_out(.a(arrdiv32_mux2to1290_xor0[0]), .b(b[12]), .bin(arrdiv32_fs331_or0[0]), .fs_xor1(arrdiv32_fs332_xor1), .fs_or0(arrdiv32_fs332_or0));
  fs fs_arrdiv32_fs333_out(.a(arrdiv32_mux2to1291_xor0[0]), .b(b[13]), .bin(arrdiv32_fs332_or0[0]), .fs_xor1(arrdiv32_fs333_xor1), .fs_or0(arrdiv32_fs333_or0));
  fs fs_arrdiv32_fs334_out(.a(arrdiv32_mux2to1292_xor0[0]), .b(b[14]), .bin(arrdiv32_fs333_or0[0]), .fs_xor1(arrdiv32_fs334_xor1), .fs_or0(arrdiv32_fs334_or0));
  fs fs_arrdiv32_fs335_out(.a(arrdiv32_mux2to1293_xor0[0]), .b(b[15]), .bin(arrdiv32_fs334_or0[0]), .fs_xor1(arrdiv32_fs335_xor1), .fs_or0(arrdiv32_fs335_or0));
  fs fs_arrdiv32_fs336_out(.a(arrdiv32_mux2to1294_xor0[0]), .b(b[16]), .bin(arrdiv32_fs335_or0[0]), .fs_xor1(arrdiv32_fs336_xor1), .fs_or0(arrdiv32_fs336_or0));
  fs fs_arrdiv32_fs337_out(.a(arrdiv32_mux2to1295_xor0[0]), .b(b[17]), .bin(arrdiv32_fs336_or0[0]), .fs_xor1(arrdiv32_fs337_xor1), .fs_or0(arrdiv32_fs337_or0));
  fs fs_arrdiv32_fs338_out(.a(arrdiv32_mux2to1296_xor0[0]), .b(b[18]), .bin(arrdiv32_fs337_or0[0]), .fs_xor1(arrdiv32_fs338_xor1), .fs_or0(arrdiv32_fs338_or0));
  fs fs_arrdiv32_fs339_out(.a(arrdiv32_mux2to1297_xor0[0]), .b(b[19]), .bin(arrdiv32_fs338_or0[0]), .fs_xor1(arrdiv32_fs339_xor1), .fs_or0(arrdiv32_fs339_or0));
  fs fs_arrdiv32_fs340_out(.a(arrdiv32_mux2to1298_xor0[0]), .b(b[20]), .bin(arrdiv32_fs339_or0[0]), .fs_xor1(arrdiv32_fs340_xor1), .fs_or0(arrdiv32_fs340_or0));
  fs fs_arrdiv32_fs341_out(.a(arrdiv32_mux2to1299_xor0[0]), .b(b[21]), .bin(arrdiv32_fs340_or0[0]), .fs_xor1(arrdiv32_fs341_xor1), .fs_or0(arrdiv32_fs341_or0));
  fs fs_arrdiv32_fs342_out(.a(arrdiv32_mux2to1300_xor0[0]), .b(b[22]), .bin(arrdiv32_fs341_or0[0]), .fs_xor1(arrdiv32_fs342_xor1), .fs_or0(arrdiv32_fs342_or0));
  fs fs_arrdiv32_fs343_out(.a(arrdiv32_mux2to1301_xor0[0]), .b(b[23]), .bin(arrdiv32_fs342_or0[0]), .fs_xor1(arrdiv32_fs343_xor1), .fs_or0(arrdiv32_fs343_or0));
  fs fs_arrdiv32_fs344_out(.a(arrdiv32_mux2to1302_xor0[0]), .b(b[24]), .bin(arrdiv32_fs343_or0[0]), .fs_xor1(arrdiv32_fs344_xor1), .fs_or0(arrdiv32_fs344_or0));
  fs fs_arrdiv32_fs345_out(.a(arrdiv32_mux2to1303_xor0[0]), .b(b[25]), .bin(arrdiv32_fs344_or0[0]), .fs_xor1(arrdiv32_fs345_xor1), .fs_or0(arrdiv32_fs345_or0));
  fs fs_arrdiv32_fs346_out(.a(arrdiv32_mux2to1304_xor0[0]), .b(b[26]), .bin(arrdiv32_fs345_or0[0]), .fs_xor1(arrdiv32_fs346_xor1), .fs_or0(arrdiv32_fs346_or0));
  fs fs_arrdiv32_fs347_out(.a(arrdiv32_mux2to1305_xor0[0]), .b(b[27]), .bin(arrdiv32_fs346_or0[0]), .fs_xor1(arrdiv32_fs347_xor1), .fs_or0(arrdiv32_fs347_or0));
  fs fs_arrdiv32_fs348_out(.a(arrdiv32_mux2to1306_xor0[0]), .b(b[28]), .bin(arrdiv32_fs347_or0[0]), .fs_xor1(arrdiv32_fs348_xor1), .fs_or0(arrdiv32_fs348_or0));
  fs fs_arrdiv32_fs349_out(.a(arrdiv32_mux2to1307_xor0[0]), .b(b[29]), .bin(arrdiv32_fs348_or0[0]), .fs_xor1(arrdiv32_fs349_xor1), .fs_or0(arrdiv32_fs349_or0));
  fs fs_arrdiv32_fs350_out(.a(arrdiv32_mux2to1308_xor0[0]), .b(b[30]), .bin(arrdiv32_fs349_or0[0]), .fs_xor1(arrdiv32_fs350_xor1), .fs_or0(arrdiv32_fs350_or0));
  fs fs_arrdiv32_fs351_out(.a(arrdiv32_mux2to1309_xor0[0]), .b(b[31]), .bin(arrdiv32_fs350_or0[0]), .fs_xor1(arrdiv32_fs351_xor1), .fs_or0(arrdiv32_fs351_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1310_out(.d0(arrdiv32_fs320_xor0[0]), .d1(a[21]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1310_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1311_out(.d0(arrdiv32_fs321_xor1[0]), .d1(arrdiv32_mux2to1279_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1311_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1312_out(.d0(arrdiv32_fs322_xor1[0]), .d1(arrdiv32_mux2to1280_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1312_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1313_out(.d0(arrdiv32_fs323_xor1[0]), .d1(arrdiv32_mux2to1281_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1313_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1314_out(.d0(arrdiv32_fs324_xor1[0]), .d1(arrdiv32_mux2to1282_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1314_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1315_out(.d0(arrdiv32_fs325_xor1[0]), .d1(arrdiv32_mux2to1283_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1315_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1316_out(.d0(arrdiv32_fs326_xor1[0]), .d1(arrdiv32_mux2to1284_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1316_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1317_out(.d0(arrdiv32_fs327_xor1[0]), .d1(arrdiv32_mux2to1285_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1317_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1318_out(.d0(arrdiv32_fs328_xor1[0]), .d1(arrdiv32_mux2to1286_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1318_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1319_out(.d0(arrdiv32_fs329_xor1[0]), .d1(arrdiv32_mux2to1287_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1319_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1320_out(.d0(arrdiv32_fs330_xor1[0]), .d1(arrdiv32_mux2to1288_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1320_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1321_out(.d0(arrdiv32_fs331_xor1[0]), .d1(arrdiv32_mux2to1289_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1321_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1322_out(.d0(arrdiv32_fs332_xor1[0]), .d1(arrdiv32_mux2to1290_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1322_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1323_out(.d0(arrdiv32_fs333_xor1[0]), .d1(arrdiv32_mux2to1291_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1323_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1324_out(.d0(arrdiv32_fs334_xor1[0]), .d1(arrdiv32_mux2to1292_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1324_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1325_out(.d0(arrdiv32_fs335_xor1[0]), .d1(arrdiv32_mux2to1293_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1325_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1326_out(.d0(arrdiv32_fs336_xor1[0]), .d1(arrdiv32_mux2to1294_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1326_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1327_out(.d0(arrdiv32_fs337_xor1[0]), .d1(arrdiv32_mux2to1295_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1327_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1328_out(.d0(arrdiv32_fs338_xor1[0]), .d1(arrdiv32_mux2to1296_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1328_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1329_out(.d0(arrdiv32_fs339_xor1[0]), .d1(arrdiv32_mux2to1297_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1329_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1330_out(.d0(arrdiv32_fs340_xor1[0]), .d1(arrdiv32_mux2to1298_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1330_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1331_out(.d0(arrdiv32_fs341_xor1[0]), .d1(arrdiv32_mux2to1299_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1331_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1332_out(.d0(arrdiv32_fs342_xor1[0]), .d1(arrdiv32_mux2to1300_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1332_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1333_out(.d0(arrdiv32_fs343_xor1[0]), .d1(arrdiv32_mux2to1301_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1333_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1334_out(.d0(arrdiv32_fs344_xor1[0]), .d1(arrdiv32_mux2to1302_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1334_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1335_out(.d0(arrdiv32_fs345_xor1[0]), .d1(arrdiv32_mux2to1303_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1335_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1336_out(.d0(arrdiv32_fs346_xor1[0]), .d1(arrdiv32_mux2to1304_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1336_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1337_out(.d0(arrdiv32_fs347_xor1[0]), .d1(arrdiv32_mux2to1305_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1337_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1338_out(.d0(arrdiv32_fs348_xor1[0]), .d1(arrdiv32_mux2to1306_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1338_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1339_out(.d0(arrdiv32_fs349_xor1[0]), .d1(arrdiv32_mux2to1307_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1339_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1340_out(.d0(arrdiv32_fs350_xor1[0]), .d1(arrdiv32_mux2to1308_xor0[0]), .sel(arrdiv32_fs351_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1340_xor0));
  not_gate not_gate_arrdiv32_not10(.a(arrdiv32_fs351_or0[0]), .out(arrdiv32_not10));
  fs fs_arrdiv32_fs352_out(.a(a[20]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs352_xor0), .fs_or0(arrdiv32_fs352_and0));
  fs fs_arrdiv32_fs353_out(.a(arrdiv32_mux2to1310_xor0[0]), .b(b[1]), .bin(arrdiv32_fs352_and0[0]), .fs_xor1(arrdiv32_fs353_xor1), .fs_or0(arrdiv32_fs353_or0));
  fs fs_arrdiv32_fs354_out(.a(arrdiv32_mux2to1311_xor0[0]), .b(b[2]), .bin(arrdiv32_fs353_or0[0]), .fs_xor1(arrdiv32_fs354_xor1), .fs_or0(arrdiv32_fs354_or0));
  fs fs_arrdiv32_fs355_out(.a(arrdiv32_mux2to1312_xor0[0]), .b(b[3]), .bin(arrdiv32_fs354_or0[0]), .fs_xor1(arrdiv32_fs355_xor1), .fs_or0(arrdiv32_fs355_or0));
  fs fs_arrdiv32_fs356_out(.a(arrdiv32_mux2to1313_xor0[0]), .b(b[4]), .bin(arrdiv32_fs355_or0[0]), .fs_xor1(arrdiv32_fs356_xor1), .fs_or0(arrdiv32_fs356_or0));
  fs fs_arrdiv32_fs357_out(.a(arrdiv32_mux2to1314_xor0[0]), .b(b[5]), .bin(arrdiv32_fs356_or0[0]), .fs_xor1(arrdiv32_fs357_xor1), .fs_or0(arrdiv32_fs357_or0));
  fs fs_arrdiv32_fs358_out(.a(arrdiv32_mux2to1315_xor0[0]), .b(b[6]), .bin(arrdiv32_fs357_or0[0]), .fs_xor1(arrdiv32_fs358_xor1), .fs_or0(arrdiv32_fs358_or0));
  fs fs_arrdiv32_fs359_out(.a(arrdiv32_mux2to1316_xor0[0]), .b(b[7]), .bin(arrdiv32_fs358_or0[0]), .fs_xor1(arrdiv32_fs359_xor1), .fs_or0(arrdiv32_fs359_or0));
  fs fs_arrdiv32_fs360_out(.a(arrdiv32_mux2to1317_xor0[0]), .b(b[8]), .bin(arrdiv32_fs359_or0[0]), .fs_xor1(arrdiv32_fs360_xor1), .fs_or0(arrdiv32_fs360_or0));
  fs fs_arrdiv32_fs361_out(.a(arrdiv32_mux2to1318_xor0[0]), .b(b[9]), .bin(arrdiv32_fs360_or0[0]), .fs_xor1(arrdiv32_fs361_xor1), .fs_or0(arrdiv32_fs361_or0));
  fs fs_arrdiv32_fs362_out(.a(arrdiv32_mux2to1319_xor0[0]), .b(b[10]), .bin(arrdiv32_fs361_or0[0]), .fs_xor1(arrdiv32_fs362_xor1), .fs_or0(arrdiv32_fs362_or0));
  fs fs_arrdiv32_fs363_out(.a(arrdiv32_mux2to1320_xor0[0]), .b(b[11]), .bin(arrdiv32_fs362_or0[0]), .fs_xor1(arrdiv32_fs363_xor1), .fs_or0(arrdiv32_fs363_or0));
  fs fs_arrdiv32_fs364_out(.a(arrdiv32_mux2to1321_xor0[0]), .b(b[12]), .bin(arrdiv32_fs363_or0[0]), .fs_xor1(arrdiv32_fs364_xor1), .fs_or0(arrdiv32_fs364_or0));
  fs fs_arrdiv32_fs365_out(.a(arrdiv32_mux2to1322_xor0[0]), .b(b[13]), .bin(arrdiv32_fs364_or0[0]), .fs_xor1(arrdiv32_fs365_xor1), .fs_or0(arrdiv32_fs365_or0));
  fs fs_arrdiv32_fs366_out(.a(arrdiv32_mux2to1323_xor0[0]), .b(b[14]), .bin(arrdiv32_fs365_or0[0]), .fs_xor1(arrdiv32_fs366_xor1), .fs_or0(arrdiv32_fs366_or0));
  fs fs_arrdiv32_fs367_out(.a(arrdiv32_mux2to1324_xor0[0]), .b(b[15]), .bin(arrdiv32_fs366_or0[0]), .fs_xor1(arrdiv32_fs367_xor1), .fs_or0(arrdiv32_fs367_or0));
  fs fs_arrdiv32_fs368_out(.a(arrdiv32_mux2to1325_xor0[0]), .b(b[16]), .bin(arrdiv32_fs367_or0[0]), .fs_xor1(arrdiv32_fs368_xor1), .fs_or0(arrdiv32_fs368_or0));
  fs fs_arrdiv32_fs369_out(.a(arrdiv32_mux2to1326_xor0[0]), .b(b[17]), .bin(arrdiv32_fs368_or0[0]), .fs_xor1(arrdiv32_fs369_xor1), .fs_or0(arrdiv32_fs369_or0));
  fs fs_arrdiv32_fs370_out(.a(arrdiv32_mux2to1327_xor0[0]), .b(b[18]), .bin(arrdiv32_fs369_or0[0]), .fs_xor1(arrdiv32_fs370_xor1), .fs_or0(arrdiv32_fs370_or0));
  fs fs_arrdiv32_fs371_out(.a(arrdiv32_mux2to1328_xor0[0]), .b(b[19]), .bin(arrdiv32_fs370_or0[0]), .fs_xor1(arrdiv32_fs371_xor1), .fs_or0(arrdiv32_fs371_or0));
  fs fs_arrdiv32_fs372_out(.a(arrdiv32_mux2to1329_xor0[0]), .b(b[20]), .bin(arrdiv32_fs371_or0[0]), .fs_xor1(arrdiv32_fs372_xor1), .fs_or0(arrdiv32_fs372_or0));
  fs fs_arrdiv32_fs373_out(.a(arrdiv32_mux2to1330_xor0[0]), .b(b[21]), .bin(arrdiv32_fs372_or0[0]), .fs_xor1(arrdiv32_fs373_xor1), .fs_or0(arrdiv32_fs373_or0));
  fs fs_arrdiv32_fs374_out(.a(arrdiv32_mux2to1331_xor0[0]), .b(b[22]), .bin(arrdiv32_fs373_or0[0]), .fs_xor1(arrdiv32_fs374_xor1), .fs_or0(arrdiv32_fs374_or0));
  fs fs_arrdiv32_fs375_out(.a(arrdiv32_mux2to1332_xor0[0]), .b(b[23]), .bin(arrdiv32_fs374_or0[0]), .fs_xor1(arrdiv32_fs375_xor1), .fs_or0(arrdiv32_fs375_or0));
  fs fs_arrdiv32_fs376_out(.a(arrdiv32_mux2to1333_xor0[0]), .b(b[24]), .bin(arrdiv32_fs375_or0[0]), .fs_xor1(arrdiv32_fs376_xor1), .fs_or0(arrdiv32_fs376_or0));
  fs fs_arrdiv32_fs377_out(.a(arrdiv32_mux2to1334_xor0[0]), .b(b[25]), .bin(arrdiv32_fs376_or0[0]), .fs_xor1(arrdiv32_fs377_xor1), .fs_or0(arrdiv32_fs377_or0));
  fs fs_arrdiv32_fs378_out(.a(arrdiv32_mux2to1335_xor0[0]), .b(b[26]), .bin(arrdiv32_fs377_or0[0]), .fs_xor1(arrdiv32_fs378_xor1), .fs_or0(arrdiv32_fs378_or0));
  fs fs_arrdiv32_fs379_out(.a(arrdiv32_mux2to1336_xor0[0]), .b(b[27]), .bin(arrdiv32_fs378_or0[0]), .fs_xor1(arrdiv32_fs379_xor1), .fs_or0(arrdiv32_fs379_or0));
  fs fs_arrdiv32_fs380_out(.a(arrdiv32_mux2to1337_xor0[0]), .b(b[28]), .bin(arrdiv32_fs379_or0[0]), .fs_xor1(arrdiv32_fs380_xor1), .fs_or0(arrdiv32_fs380_or0));
  fs fs_arrdiv32_fs381_out(.a(arrdiv32_mux2to1338_xor0[0]), .b(b[29]), .bin(arrdiv32_fs380_or0[0]), .fs_xor1(arrdiv32_fs381_xor1), .fs_or0(arrdiv32_fs381_or0));
  fs fs_arrdiv32_fs382_out(.a(arrdiv32_mux2to1339_xor0[0]), .b(b[30]), .bin(arrdiv32_fs381_or0[0]), .fs_xor1(arrdiv32_fs382_xor1), .fs_or0(arrdiv32_fs382_or0));
  fs fs_arrdiv32_fs383_out(.a(arrdiv32_mux2to1340_xor0[0]), .b(b[31]), .bin(arrdiv32_fs382_or0[0]), .fs_xor1(arrdiv32_fs383_xor1), .fs_or0(arrdiv32_fs383_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1341_out(.d0(arrdiv32_fs352_xor0[0]), .d1(a[20]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1341_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1342_out(.d0(arrdiv32_fs353_xor1[0]), .d1(arrdiv32_mux2to1310_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1342_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1343_out(.d0(arrdiv32_fs354_xor1[0]), .d1(arrdiv32_mux2to1311_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1343_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1344_out(.d0(arrdiv32_fs355_xor1[0]), .d1(arrdiv32_mux2to1312_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1344_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1345_out(.d0(arrdiv32_fs356_xor1[0]), .d1(arrdiv32_mux2to1313_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1345_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1346_out(.d0(arrdiv32_fs357_xor1[0]), .d1(arrdiv32_mux2to1314_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1346_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1347_out(.d0(arrdiv32_fs358_xor1[0]), .d1(arrdiv32_mux2to1315_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1347_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1348_out(.d0(arrdiv32_fs359_xor1[0]), .d1(arrdiv32_mux2to1316_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1348_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1349_out(.d0(arrdiv32_fs360_xor1[0]), .d1(arrdiv32_mux2to1317_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1349_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1350_out(.d0(arrdiv32_fs361_xor1[0]), .d1(arrdiv32_mux2to1318_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1350_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1351_out(.d0(arrdiv32_fs362_xor1[0]), .d1(arrdiv32_mux2to1319_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1351_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1352_out(.d0(arrdiv32_fs363_xor1[0]), .d1(arrdiv32_mux2to1320_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1352_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1353_out(.d0(arrdiv32_fs364_xor1[0]), .d1(arrdiv32_mux2to1321_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1353_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1354_out(.d0(arrdiv32_fs365_xor1[0]), .d1(arrdiv32_mux2to1322_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1354_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1355_out(.d0(arrdiv32_fs366_xor1[0]), .d1(arrdiv32_mux2to1323_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1355_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1356_out(.d0(arrdiv32_fs367_xor1[0]), .d1(arrdiv32_mux2to1324_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1356_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1357_out(.d0(arrdiv32_fs368_xor1[0]), .d1(arrdiv32_mux2to1325_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1357_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1358_out(.d0(arrdiv32_fs369_xor1[0]), .d1(arrdiv32_mux2to1326_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1358_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1359_out(.d0(arrdiv32_fs370_xor1[0]), .d1(arrdiv32_mux2to1327_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1359_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1360_out(.d0(arrdiv32_fs371_xor1[0]), .d1(arrdiv32_mux2to1328_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1360_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1361_out(.d0(arrdiv32_fs372_xor1[0]), .d1(arrdiv32_mux2to1329_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1361_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1362_out(.d0(arrdiv32_fs373_xor1[0]), .d1(arrdiv32_mux2to1330_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1362_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1363_out(.d0(arrdiv32_fs374_xor1[0]), .d1(arrdiv32_mux2to1331_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1363_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1364_out(.d0(arrdiv32_fs375_xor1[0]), .d1(arrdiv32_mux2to1332_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1364_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1365_out(.d0(arrdiv32_fs376_xor1[0]), .d1(arrdiv32_mux2to1333_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1365_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1366_out(.d0(arrdiv32_fs377_xor1[0]), .d1(arrdiv32_mux2to1334_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1366_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1367_out(.d0(arrdiv32_fs378_xor1[0]), .d1(arrdiv32_mux2to1335_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1367_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1368_out(.d0(arrdiv32_fs379_xor1[0]), .d1(arrdiv32_mux2to1336_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1368_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1369_out(.d0(arrdiv32_fs380_xor1[0]), .d1(arrdiv32_mux2to1337_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1369_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1370_out(.d0(arrdiv32_fs381_xor1[0]), .d1(arrdiv32_mux2to1338_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1370_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1371_out(.d0(arrdiv32_fs382_xor1[0]), .d1(arrdiv32_mux2to1339_xor0[0]), .sel(arrdiv32_fs383_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1371_xor0));
  not_gate not_gate_arrdiv32_not11(.a(arrdiv32_fs383_or0[0]), .out(arrdiv32_not11));
  fs fs_arrdiv32_fs384_out(.a(a[19]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs384_xor0), .fs_or0(arrdiv32_fs384_and0));
  fs fs_arrdiv32_fs385_out(.a(arrdiv32_mux2to1341_xor0[0]), .b(b[1]), .bin(arrdiv32_fs384_and0[0]), .fs_xor1(arrdiv32_fs385_xor1), .fs_or0(arrdiv32_fs385_or0));
  fs fs_arrdiv32_fs386_out(.a(arrdiv32_mux2to1342_xor0[0]), .b(b[2]), .bin(arrdiv32_fs385_or0[0]), .fs_xor1(arrdiv32_fs386_xor1), .fs_or0(arrdiv32_fs386_or0));
  fs fs_arrdiv32_fs387_out(.a(arrdiv32_mux2to1343_xor0[0]), .b(b[3]), .bin(arrdiv32_fs386_or0[0]), .fs_xor1(arrdiv32_fs387_xor1), .fs_or0(arrdiv32_fs387_or0));
  fs fs_arrdiv32_fs388_out(.a(arrdiv32_mux2to1344_xor0[0]), .b(b[4]), .bin(arrdiv32_fs387_or0[0]), .fs_xor1(arrdiv32_fs388_xor1), .fs_or0(arrdiv32_fs388_or0));
  fs fs_arrdiv32_fs389_out(.a(arrdiv32_mux2to1345_xor0[0]), .b(b[5]), .bin(arrdiv32_fs388_or0[0]), .fs_xor1(arrdiv32_fs389_xor1), .fs_or0(arrdiv32_fs389_or0));
  fs fs_arrdiv32_fs390_out(.a(arrdiv32_mux2to1346_xor0[0]), .b(b[6]), .bin(arrdiv32_fs389_or0[0]), .fs_xor1(arrdiv32_fs390_xor1), .fs_or0(arrdiv32_fs390_or0));
  fs fs_arrdiv32_fs391_out(.a(arrdiv32_mux2to1347_xor0[0]), .b(b[7]), .bin(arrdiv32_fs390_or0[0]), .fs_xor1(arrdiv32_fs391_xor1), .fs_or0(arrdiv32_fs391_or0));
  fs fs_arrdiv32_fs392_out(.a(arrdiv32_mux2to1348_xor0[0]), .b(b[8]), .bin(arrdiv32_fs391_or0[0]), .fs_xor1(arrdiv32_fs392_xor1), .fs_or0(arrdiv32_fs392_or0));
  fs fs_arrdiv32_fs393_out(.a(arrdiv32_mux2to1349_xor0[0]), .b(b[9]), .bin(arrdiv32_fs392_or0[0]), .fs_xor1(arrdiv32_fs393_xor1), .fs_or0(arrdiv32_fs393_or0));
  fs fs_arrdiv32_fs394_out(.a(arrdiv32_mux2to1350_xor0[0]), .b(b[10]), .bin(arrdiv32_fs393_or0[0]), .fs_xor1(arrdiv32_fs394_xor1), .fs_or0(arrdiv32_fs394_or0));
  fs fs_arrdiv32_fs395_out(.a(arrdiv32_mux2to1351_xor0[0]), .b(b[11]), .bin(arrdiv32_fs394_or0[0]), .fs_xor1(arrdiv32_fs395_xor1), .fs_or0(arrdiv32_fs395_or0));
  fs fs_arrdiv32_fs396_out(.a(arrdiv32_mux2to1352_xor0[0]), .b(b[12]), .bin(arrdiv32_fs395_or0[0]), .fs_xor1(arrdiv32_fs396_xor1), .fs_or0(arrdiv32_fs396_or0));
  fs fs_arrdiv32_fs397_out(.a(arrdiv32_mux2to1353_xor0[0]), .b(b[13]), .bin(arrdiv32_fs396_or0[0]), .fs_xor1(arrdiv32_fs397_xor1), .fs_or0(arrdiv32_fs397_or0));
  fs fs_arrdiv32_fs398_out(.a(arrdiv32_mux2to1354_xor0[0]), .b(b[14]), .bin(arrdiv32_fs397_or0[0]), .fs_xor1(arrdiv32_fs398_xor1), .fs_or0(arrdiv32_fs398_or0));
  fs fs_arrdiv32_fs399_out(.a(arrdiv32_mux2to1355_xor0[0]), .b(b[15]), .bin(arrdiv32_fs398_or0[0]), .fs_xor1(arrdiv32_fs399_xor1), .fs_or0(arrdiv32_fs399_or0));
  fs fs_arrdiv32_fs400_out(.a(arrdiv32_mux2to1356_xor0[0]), .b(b[16]), .bin(arrdiv32_fs399_or0[0]), .fs_xor1(arrdiv32_fs400_xor1), .fs_or0(arrdiv32_fs400_or0));
  fs fs_arrdiv32_fs401_out(.a(arrdiv32_mux2to1357_xor0[0]), .b(b[17]), .bin(arrdiv32_fs400_or0[0]), .fs_xor1(arrdiv32_fs401_xor1), .fs_or0(arrdiv32_fs401_or0));
  fs fs_arrdiv32_fs402_out(.a(arrdiv32_mux2to1358_xor0[0]), .b(b[18]), .bin(arrdiv32_fs401_or0[0]), .fs_xor1(arrdiv32_fs402_xor1), .fs_or0(arrdiv32_fs402_or0));
  fs fs_arrdiv32_fs403_out(.a(arrdiv32_mux2to1359_xor0[0]), .b(b[19]), .bin(arrdiv32_fs402_or0[0]), .fs_xor1(arrdiv32_fs403_xor1), .fs_or0(arrdiv32_fs403_or0));
  fs fs_arrdiv32_fs404_out(.a(arrdiv32_mux2to1360_xor0[0]), .b(b[20]), .bin(arrdiv32_fs403_or0[0]), .fs_xor1(arrdiv32_fs404_xor1), .fs_or0(arrdiv32_fs404_or0));
  fs fs_arrdiv32_fs405_out(.a(arrdiv32_mux2to1361_xor0[0]), .b(b[21]), .bin(arrdiv32_fs404_or0[0]), .fs_xor1(arrdiv32_fs405_xor1), .fs_or0(arrdiv32_fs405_or0));
  fs fs_arrdiv32_fs406_out(.a(arrdiv32_mux2to1362_xor0[0]), .b(b[22]), .bin(arrdiv32_fs405_or0[0]), .fs_xor1(arrdiv32_fs406_xor1), .fs_or0(arrdiv32_fs406_or0));
  fs fs_arrdiv32_fs407_out(.a(arrdiv32_mux2to1363_xor0[0]), .b(b[23]), .bin(arrdiv32_fs406_or0[0]), .fs_xor1(arrdiv32_fs407_xor1), .fs_or0(arrdiv32_fs407_or0));
  fs fs_arrdiv32_fs408_out(.a(arrdiv32_mux2to1364_xor0[0]), .b(b[24]), .bin(arrdiv32_fs407_or0[0]), .fs_xor1(arrdiv32_fs408_xor1), .fs_or0(arrdiv32_fs408_or0));
  fs fs_arrdiv32_fs409_out(.a(arrdiv32_mux2to1365_xor0[0]), .b(b[25]), .bin(arrdiv32_fs408_or0[0]), .fs_xor1(arrdiv32_fs409_xor1), .fs_or0(arrdiv32_fs409_or0));
  fs fs_arrdiv32_fs410_out(.a(arrdiv32_mux2to1366_xor0[0]), .b(b[26]), .bin(arrdiv32_fs409_or0[0]), .fs_xor1(arrdiv32_fs410_xor1), .fs_or0(arrdiv32_fs410_or0));
  fs fs_arrdiv32_fs411_out(.a(arrdiv32_mux2to1367_xor0[0]), .b(b[27]), .bin(arrdiv32_fs410_or0[0]), .fs_xor1(arrdiv32_fs411_xor1), .fs_or0(arrdiv32_fs411_or0));
  fs fs_arrdiv32_fs412_out(.a(arrdiv32_mux2to1368_xor0[0]), .b(b[28]), .bin(arrdiv32_fs411_or0[0]), .fs_xor1(arrdiv32_fs412_xor1), .fs_or0(arrdiv32_fs412_or0));
  fs fs_arrdiv32_fs413_out(.a(arrdiv32_mux2to1369_xor0[0]), .b(b[29]), .bin(arrdiv32_fs412_or0[0]), .fs_xor1(arrdiv32_fs413_xor1), .fs_or0(arrdiv32_fs413_or0));
  fs fs_arrdiv32_fs414_out(.a(arrdiv32_mux2to1370_xor0[0]), .b(b[30]), .bin(arrdiv32_fs413_or0[0]), .fs_xor1(arrdiv32_fs414_xor1), .fs_or0(arrdiv32_fs414_or0));
  fs fs_arrdiv32_fs415_out(.a(arrdiv32_mux2to1371_xor0[0]), .b(b[31]), .bin(arrdiv32_fs414_or0[0]), .fs_xor1(arrdiv32_fs415_xor1), .fs_or0(arrdiv32_fs415_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1372_out(.d0(arrdiv32_fs384_xor0[0]), .d1(a[19]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1372_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1373_out(.d0(arrdiv32_fs385_xor1[0]), .d1(arrdiv32_mux2to1341_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1373_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1374_out(.d0(arrdiv32_fs386_xor1[0]), .d1(arrdiv32_mux2to1342_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1374_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1375_out(.d0(arrdiv32_fs387_xor1[0]), .d1(arrdiv32_mux2to1343_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1375_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1376_out(.d0(arrdiv32_fs388_xor1[0]), .d1(arrdiv32_mux2to1344_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1376_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1377_out(.d0(arrdiv32_fs389_xor1[0]), .d1(arrdiv32_mux2to1345_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1377_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1378_out(.d0(arrdiv32_fs390_xor1[0]), .d1(arrdiv32_mux2to1346_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1378_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1379_out(.d0(arrdiv32_fs391_xor1[0]), .d1(arrdiv32_mux2to1347_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1379_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1380_out(.d0(arrdiv32_fs392_xor1[0]), .d1(arrdiv32_mux2to1348_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1380_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1381_out(.d0(arrdiv32_fs393_xor1[0]), .d1(arrdiv32_mux2to1349_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1381_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1382_out(.d0(arrdiv32_fs394_xor1[0]), .d1(arrdiv32_mux2to1350_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1382_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1383_out(.d0(arrdiv32_fs395_xor1[0]), .d1(arrdiv32_mux2to1351_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1383_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1384_out(.d0(arrdiv32_fs396_xor1[0]), .d1(arrdiv32_mux2to1352_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1384_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1385_out(.d0(arrdiv32_fs397_xor1[0]), .d1(arrdiv32_mux2to1353_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1385_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1386_out(.d0(arrdiv32_fs398_xor1[0]), .d1(arrdiv32_mux2to1354_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1386_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1387_out(.d0(arrdiv32_fs399_xor1[0]), .d1(arrdiv32_mux2to1355_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1387_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1388_out(.d0(arrdiv32_fs400_xor1[0]), .d1(arrdiv32_mux2to1356_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1388_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1389_out(.d0(arrdiv32_fs401_xor1[0]), .d1(arrdiv32_mux2to1357_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1389_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1390_out(.d0(arrdiv32_fs402_xor1[0]), .d1(arrdiv32_mux2to1358_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1390_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1391_out(.d0(arrdiv32_fs403_xor1[0]), .d1(arrdiv32_mux2to1359_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1391_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1392_out(.d0(arrdiv32_fs404_xor1[0]), .d1(arrdiv32_mux2to1360_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1392_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1393_out(.d0(arrdiv32_fs405_xor1[0]), .d1(arrdiv32_mux2to1361_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1393_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1394_out(.d0(arrdiv32_fs406_xor1[0]), .d1(arrdiv32_mux2to1362_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1394_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1395_out(.d0(arrdiv32_fs407_xor1[0]), .d1(arrdiv32_mux2to1363_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1395_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1396_out(.d0(arrdiv32_fs408_xor1[0]), .d1(arrdiv32_mux2to1364_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1396_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1397_out(.d0(arrdiv32_fs409_xor1[0]), .d1(arrdiv32_mux2to1365_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1397_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1398_out(.d0(arrdiv32_fs410_xor1[0]), .d1(arrdiv32_mux2to1366_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1398_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1399_out(.d0(arrdiv32_fs411_xor1[0]), .d1(arrdiv32_mux2to1367_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1399_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1400_out(.d0(arrdiv32_fs412_xor1[0]), .d1(arrdiv32_mux2to1368_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1400_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1401_out(.d0(arrdiv32_fs413_xor1[0]), .d1(arrdiv32_mux2to1369_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1401_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1402_out(.d0(arrdiv32_fs414_xor1[0]), .d1(arrdiv32_mux2to1370_xor0[0]), .sel(arrdiv32_fs415_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1402_xor0));
  not_gate not_gate_arrdiv32_not12(.a(arrdiv32_fs415_or0[0]), .out(arrdiv32_not12));
  fs fs_arrdiv32_fs416_out(.a(a[18]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs416_xor0), .fs_or0(arrdiv32_fs416_and0));
  fs fs_arrdiv32_fs417_out(.a(arrdiv32_mux2to1372_xor0[0]), .b(b[1]), .bin(arrdiv32_fs416_and0[0]), .fs_xor1(arrdiv32_fs417_xor1), .fs_or0(arrdiv32_fs417_or0));
  fs fs_arrdiv32_fs418_out(.a(arrdiv32_mux2to1373_xor0[0]), .b(b[2]), .bin(arrdiv32_fs417_or0[0]), .fs_xor1(arrdiv32_fs418_xor1), .fs_or0(arrdiv32_fs418_or0));
  fs fs_arrdiv32_fs419_out(.a(arrdiv32_mux2to1374_xor0[0]), .b(b[3]), .bin(arrdiv32_fs418_or0[0]), .fs_xor1(arrdiv32_fs419_xor1), .fs_or0(arrdiv32_fs419_or0));
  fs fs_arrdiv32_fs420_out(.a(arrdiv32_mux2to1375_xor0[0]), .b(b[4]), .bin(arrdiv32_fs419_or0[0]), .fs_xor1(arrdiv32_fs420_xor1), .fs_or0(arrdiv32_fs420_or0));
  fs fs_arrdiv32_fs421_out(.a(arrdiv32_mux2to1376_xor0[0]), .b(b[5]), .bin(arrdiv32_fs420_or0[0]), .fs_xor1(arrdiv32_fs421_xor1), .fs_or0(arrdiv32_fs421_or0));
  fs fs_arrdiv32_fs422_out(.a(arrdiv32_mux2to1377_xor0[0]), .b(b[6]), .bin(arrdiv32_fs421_or0[0]), .fs_xor1(arrdiv32_fs422_xor1), .fs_or0(arrdiv32_fs422_or0));
  fs fs_arrdiv32_fs423_out(.a(arrdiv32_mux2to1378_xor0[0]), .b(b[7]), .bin(arrdiv32_fs422_or0[0]), .fs_xor1(arrdiv32_fs423_xor1), .fs_or0(arrdiv32_fs423_or0));
  fs fs_arrdiv32_fs424_out(.a(arrdiv32_mux2to1379_xor0[0]), .b(b[8]), .bin(arrdiv32_fs423_or0[0]), .fs_xor1(arrdiv32_fs424_xor1), .fs_or0(arrdiv32_fs424_or0));
  fs fs_arrdiv32_fs425_out(.a(arrdiv32_mux2to1380_xor0[0]), .b(b[9]), .bin(arrdiv32_fs424_or0[0]), .fs_xor1(arrdiv32_fs425_xor1), .fs_or0(arrdiv32_fs425_or0));
  fs fs_arrdiv32_fs426_out(.a(arrdiv32_mux2to1381_xor0[0]), .b(b[10]), .bin(arrdiv32_fs425_or0[0]), .fs_xor1(arrdiv32_fs426_xor1), .fs_or0(arrdiv32_fs426_or0));
  fs fs_arrdiv32_fs427_out(.a(arrdiv32_mux2to1382_xor0[0]), .b(b[11]), .bin(arrdiv32_fs426_or0[0]), .fs_xor1(arrdiv32_fs427_xor1), .fs_or0(arrdiv32_fs427_or0));
  fs fs_arrdiv32_fs428_out(.a(arrdiv32_mux2to1383_xor0[0]), .b(b[12]), .bin(arrdiv32_fs427_or0[0]), .fs_xor1(arrdiv32_fs428_xor1), .fs_or0(arrdiv32_fs428_or0));
  fs fs_arrdiv32_fs429_out(.a(arrdiv32_mux2to1384_xor0[0]), .b(b[13]), .bin(arrdiv32_fs428_or0[0]), .fs_xor1(arrdiv32_fs429_xor1), .fs_or0(arrdiv32_fs429_or0));
  fs fs_arrdiv32_fs430_out(.a(arrdiv32_mux2to1385_xor0[0]), .b(b[14]), .bin(arrdiv32_fs429_or0[0]), .fs_xor1(arrdiv32_fs430_xor1), .fs_or0(arrdiv32_fs430_or0));
  fs fs_arrdiv32_fs431_out(.a(arrdiv32_mux2to1386_xor0[0]), .b(b[15]), .bin(arrdiv32_fs430_or0[0]), .fs_xor1(arrdiv32_fs431_xor1), .fs_or0(arrdiv32_fs431_or0));
  fs fs_arrdiv32_fs432_out(.a(arrdiv32_mux2to1387_xor0[0]), .b(b[16]), .bin(arrdiv32_fs431_or0[0]), .fs_xor1(arrdiv32_fs432_xor1), .fs_or0(arrdiv32_fs432_or0));
  fs fs_arrdiv32_fs433_out(.a(arrdiv32_mux2to1388_xor0[0]), .b(b[17]), .bin(arrdiv32_fs432_or0[0]), .fs_xor1(arrdiv32_fs433_xor1), .fs_or0(arrdiv32_fs433_or0));
  fs fs_arrdiv32_fs434_out(.a(arrdiv32_mux2to1389_xor0[0]), .b(b[18]), .bin(arrdiv32_fs433_or0[0]), .fs_xor1(arrdiv32_fs434_xor1), .fs_or0(arrdiv32_fs434_or0));
  fs fs_arrdiv32_fs435_out(.a(arrdiv32_mux2to1390_xor0[0]), .b(b[19]), .bin(arrdiv32_fs434_or0[0]), .fs_xor1(arrdiv32_fs435_xor1), .fs_or0(arrdiv32_fs435_or0));
  fs fs_arrdiv32_fs436_out(.a(arrdiv32_mux2to1391_xor0[0]), .b(b[20]), .bin(arrdiv32_fs435_or0[0]), .fs_xor1(arrdiv32_fs436_xor1), .fs_or0(arrdiv32_fs436_or0));
  fs fs_arrdiv32_fs437_out(.a(arrdiv32_mux2to1392_xor0[0]), .b(b[21]), .bin(arrdiv32_fs436_or0[0]), .fs_xor1(arrdiv32_fs437_xor1), .fs_or0(arrdiv32_fs437_or0));
  fs fs_arrdiv32_fs438_out(.a(arrdiv32_mux2to1393_xor0[0]), .b(b[22]), .bin(arrdiv32_fs437_or0[0]), .fs_xor1(arrdiv32_fs438_xor1), .fs_or0(arrdiv32_fs438_or0));
  fs fs_arrdiv32_fs439_out(.a(arrdiv32_mux2to1394_xor0[0]), .b(b[23]), .bin(arrdiv32_fs438_or0[0]), .fs_xor1(arrdiv32_fs439_xor1), .fs_or0(arrdiv32_fs439_or0));
  fs fs_arrdiv32_fs440_out(.a(arrdiv32_mux2to1395_xor0[0]), .b(b[24]), .bin(arrdiv32_fs439_or0[0]), .fs_xor1(arrdiv32_fs440_xor1), .fs_or0(arrdiv32_fs440_or0));
  fs fs_arrdiv32_fs441_out(.a(arrdiv32_mux2to1396_xor0[0]), .b(b[25]), .bin(arrdiv32_fs440_or0[0]), .fs_xor1(arrdiv32_fs441_xor1), .fs_or0(arrdiv32_fs441_or0));
  fs fs_arrdiv32_fs442_out(.a(arrdiv32_mux2to1397_xor0[0]), .b(b[26]), .bin(arrdiv32_fs441_or0[0]), .fs_xor1(arrdiv32_fs442_xor1), .fs_or0(arrdiv32_fs442_or0));
  fs fs_arrdiv32_fs443_out(.a(arrdiv32_mux2to1398_xor0[0]), .b(b[27]), .bin(arrdiv32_fs442_or0[0]), .fs_xor1(arrdiv32_fs443_xor1), .fs_or0(arrdiv32_fs443_or0));
  fs fs_arrdiv32_fs444_out(.a(arrdiv32_mux2to1399_xor0[0]), .b(b[28]), .bin(arrdiv32_fs443_or0[0]), .fs_xor1(arrdiv32_fs444_xor1), .fs_or0(arrdiv32_fs444_or0));
  fs fs_arrdiv32_fs445_out(.a(arrdiv32_mux2to1400_xor0[0]), .b(b[29]), .bin(arrdiv32_fs444_or0[0]), .fs_xor1(arrdiv32_fs445_xor1), .fs_or0(arrdiv32_fs445_or0));
  fs fs_arrdiv32_fs446_out(.a(arrdiv32_mux2to1401_xor0[0]), .b(b[30]), .bin(arrdiv32_fs445_or0[0]), .fs_xor1(arrdiv32_fs446_xor1), .fs_or0(arrdiv32_fs446_or0));
  fs fs_arrdiv32_fs447_out(.a(arrdiv32_mux2to1402_xor0[0]), .b(b[31]), .bin(arrdiv32_fs446_or0[0]), .fs_xor1(arrdiv32_fs447_xor1), .fs_or0(arrdiv32_fs447_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1403_out(.d0(arrdiv32_fs416_xor0[0]), .d1(a[18]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1403_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1404_out(.d0(arrdiv32_fs417_xor1[0]), .d1(arrdiv32_mux2to1372_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1404_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1405_out(.d0(arrdiv32_fs418_xor1[0]), .d1(arrdiv32_mux2to1373_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1405_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1406_out(.d0(arrdiv32_fs419_xor1[0]), .d1(arrdiv32_mux2to1374_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1406_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1407_out(.d0(arrdiv32_fs420_xor1[0]), .d1(arrdiv32_mux2to1375_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1407_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1408_out(.d0(arrdiv32_fs421_xor1[0]), .d1(arrdiv32_mux2to1376_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1408_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1409_out(.d0(arrdiv32_fs422_xor1[0]), .d1(arrdiv32_mux2to1377_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1409_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1410_out(.d0(arrdiv32_fs423_xor1[0]), .d1(arrdiv32_mux2to1378_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1410_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1411_out(.d0(arrdiv32_fs424_xor1[0]), .d1(arrdiv32_mux2to1379_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1411_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1412_out(.d0(arrdiv32_fs425_xor1[0]), .d1(arrdiv32_mux2to1380_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1412_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1413_out(.d0(arrdiv32_fs426_xor1[0]), .d1(arrdiv32_mux2to1381_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1413_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1414_out(.d0(arrdiv32_fs427_xor1[0]), .d1(arrdiv32_mux2to1382_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1414_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1415_out(.d0(arrdiv32_fs428_xor1[0]), .d1(arrdiv32_mux2to1383_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1415_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1416_out(.d0(arrdiv32_fs429_xor1[0]), .d1(arrdiv32_mux2to1384_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1416_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1417_out(.d0(arrdiv32_fs430_xor1[0]), .d1(arrdiv32_mux2to1385_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1417_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1418_out(.d0(arrdiv32_fs431_xor1[0]), .d1(arrdiv32_mux2to1386_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1418_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1419_out(.d0(arrdiv32_fs432_xor1[0]), .d1(arrdiv32_mux2to1387_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1419_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1420_out(.d0(arrdiv32_fs433_xor1[0]), .d1(arrdiv32_mux2to1388_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1420_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1421_out(.d0(arrdiv32_fs434_xor1[0]), .d1(arrdiv32_mux2to1389_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1421_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1422_out(.d0(arrdiv32_fs435_xor1[0]), .d1(arrdiv32_mux2to1390_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1422_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1423_out(.d0(arrdiv32_fs436_xor1[0]), .d1(arrdiv32_mux2to1391_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1423_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1424_out(.d0(arrdiv32_fs437_xor1[0]), .d1(arrdiv32_mux2to1392_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1424_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1425_out(.d0(arrdiv32_fs438_xor1[0]), .d1(arrdiv32_mux2to1393_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1425_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1426_out(.d0(arrdiv32_fs439_xor1[0]), .d1(arrdiv32_mux2to1394_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1426_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1427_out(.d0(arrdiv32_fs440_xor1[0]), .d1(arrdiv32_mux2to1395_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1427_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1428_out(.d0(arrdiv32_fs441_xor1[0]), .d1(arrdiv32_mux2to1396_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1428_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1429_out(.d0(arrdiv32_fs442_xor1[0]), .d1(arrdiv32_mux2to1397_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1429_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1430_out(.d0(arrdiv32_fs443_xor1[0]), .d1(arrdiv32_mux2to1398_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1430_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1431_out(.d0(arrdiv32_fs444_xor1[0]), .d1(arrdiv32_mux2to1399_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1431_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1432_out(.d0(arrdiv32_fs445_xor1[0]), .d1(arrdiv32_mux2to1400_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1432_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1433_out(.d0(arrdiv32_fs446_xor1[0]), .d1(arrdiv32_mux2to1401_xor0[0]), .sel(arrdiv32_fs447_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1433_xor0));
  not_gate not_gate_arrdiv32_not13(.a(arrdiv32_fs447_or0[0]), .out(arrdiv32_not13));
  fs fs_arrdiv32_fs448_out(.a(a[17]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs448_xor0), .fs_or0(arrdiv32_fs448_and0));
  fs fs_arrdiv32_fs449_out(.a(arrdiv32_mux2to1403_xor0[0]), .b(b[1]), .bin(arrdiv32_fs448_and0[0]), .fs_xor1(arrdiv32_fs449_xor1), .fs_or0(arrdiv32_fs449_or0));
  fs fs_arrdiv32_fs450_out(.a(arrdiv32_mux2to1404_xor0[0]), .b(b[2]), .bin(arrdiv32_fs449_or0[0]), .fs_xor1(arrdiv32_fs450_xor1), .fs_or0(arrdiv32_fs450_or0));
  fs fs_arrdiv32_fs451_out(.a(arrdiv32_mux2to1405_xor0[0]), .b(b[3]), .bin(arrdiv32_fs450_or0[0]), .fs_xor1(arrdiv32_fs451_xor1), .fs_or0(arrdiv32_fs451_or0));
  fs fs_arrdiv32_fs452_out(.a(arrdiv32_mux2to1406_xor0[0]), .b(b[4]), .bin(arrdiv32_fs451_or0[0]), .fs_xor1(arrdiv32_fs452_xor1), .fs_or0(arrdiv32_fs452_or0));
  fs fs_arrdiv32_fs453_out(.a(arrdiv32_mux2to1407_xor0[0]), .b(b[5]), .bin(arrdiv32_fs452_or0[0]), .fs_xor1(arrdiv32_fs453_xor1), .fs_or0(arrdiv32_fs453_or0));
  fs fs_arrdiv32_fs454_out(.a(arrdiv32_mux2to1408_xor0[0]), .b(b[6]), .bin(arrdiv32_fs453_or0[0]), .fs_xor1(arrdiv32_fs454_xor1), .fs_or0(arrdiv32_fs454_or0));
  fs fs_arrdiv32_fs455_out(.a(arrdiv32_mux2to1409_xor0[0]), .b(b[7]), .bin(arrdiv32_fs454_or0[0]), .fs_xor1(arrdiv32_fs455_xor1), .fs_or0(arrdiv32_fs455_or0));
  fs fs_arrdiv32_fs456_out(.a(arrdiv32_mux2to1410_xor0[0]), .b(b[8]), .bin(arrdiv32_fs455_or0[0]), .fs_xor1(arrdiv32_fs456_xor1), .fs_or0(arrdiv32_fs456_or0));
  fs fs_arrdiv32_fs457_out(.a(arrdiv32_mux2to1411_xor0[0]), .b(b[9]), .bin(arrdiv32_fs456_or0[0]), .fs_xor1(arrdiv32_fs457_xor1), .fs_or0(arrdiv32_fs457_or0));
  fs fs_arrdiv32_fs458_out(.a(arrdiv32_mux2to1412_xor0[0]), .b(b[10]), .bin(arrdiv32_fs457_or0[0]), .fs_xor1(arrdiv32_fs458_xor1), .fs_or0(arrdiv32_fs458_or0));
  fs fs_arrdiv32_fs459_out(.a(arrdiv32_mux2to1413_xor0[0]), .b(b[11]), .bin(arrdiv32_fs458_or0[0]), .fs_xor1(arrdiv32_fs459_xor1), .fs_or0(arrdiv32_fs459_or0));
  fs fs_arrdiv32_fs460_out(.a(arrdiv32_mux2to1414_xor0[0]), .b(b[12]), .bin(arrdiv32_fs459_or0[0]), .fs_xor1(arrdiv32_fs460_xor1), .fs_or0(arrdiv32_fs460_or0));
  fs fs_arrdiv32_fs461_out(.a(arrdiv32_mux2to1415_xor0[0]), .b(b[13]), .bin(arrdiv32_fs460_or0[0]), .fs_xor1(arrdiv32_fs461_xor1), .fs_or0(arrdiv32_fs461_or0));
  fs fs_arrdiv32_fs462_out(.a(arrdiv32_mux2to1416_xor0[0]), .b(b[14]), .bin(arrdiv32_fs461_or0[0]), .fs_xor1(arrdiv32_fs462_xor1), .fs_or0(arrdiv32_fs462_or0));
  fs fs_arrdiv32_fs463_out(.a(arrdiv32_mux2to1417_xor0[0]), .b(b[15]), .bin(arrdiv32_fs462_or0[0]), .fs_xor1(arrdiv32_fs463_xor1), .fs_or0(arrdiv32_fs463_or0));
  fs fs_arrdiv32_fs464_out(.a(arrdiv32_mux2to1418_xor0[0]), .b(b[16]), .bin(arrdiv32_fs463_or0[0]), .fs_xor1(arrdiv32_fs464_xor1), .fs_or0(arrdiv32_fs464_or0));
  fs fs_arrdiv32_fs465_out(.a(arrdiv32_mux2to1419_xor0[0]), .b(b[17]), .bin(arrdiv32_fs464_or0[0]), .fs_xor1(arrdiv32_fs465_xor1), .fs_or0(arrdiv32_fs465_or0));
  fs fs_arrdiv32_fs466_out(.a(arrdiv32_mux2to1420_xor0[0]), .b(b[18]), .bin(arrdiv32_fs465_or0[0]), .fs_xor1(arrdiv32_fs466_xor1), .fs_or0(arrdiv32_fs466_or0));
  fs fs_arrdiv32_fs467_out(.a(arrdiv32_mux2to1421_xor0[0]), .b(b[19]), .bin(arrdiv32_fs466_or0[0]), .fs_xor1(arrdiv32_fs467_xor1), .fs_or0(arrdiv32_fs467_or0));
  fs fs_arrdiv32_fs468_out(.a(arrdiv32_mux2to1422_xor0[0]), .b(b[20]), .bin(arrdiv32_fs467_or0[0]), .fs_xor1(arrdiv32_fs468_xor1), .fs_or0(arrdiv32_fs468_or0));
  fs fs_arrdiv32_fs469_out(.a(arrdiv32_mux2to1423_xor0[0]), .b(b[21]), .bin(arrdiv32_fs468_or0[0]), .fs_xor1(arrdiv32_fs469_xor1), .fs_or0(arrdiv32_fs469_or0));
  fs fs_arrdiv32_fs470_out(.a(arrdiv32_mux2to1424_xor0[0]), .b(b[22]), .bin(arrdiv32_fs469_or0[0]), .fs_xor1(arrdiv32_fs470_xor1), .fs_or0(arrdiv32_fs470_or0));
  fs fs_arrdiv32_fs471_out(.a(arrdiv32_mux2to1425_xor0[0]), .b(b[23]), .bin(arrdiv32_fs470_or0[0]), .fs_xor1(arrdiv32_fs471_xor1), .fs_or0(arrdiv32_fs471_or0));
  fs fs_arrdiv32_fs472_out(.a(arrdiv32_mux2to1426_xor0[0]), .b(b[24]), .bin(arrdiv32_fs471_or0[0]), .fs_xor1(arrdiv32_fs472_xor1), .fs_or0(arrdiv32_fs472_or0));
  fs fs_arrdiv32_fs473_out(.a(arrdiv32_mux2to1427_xor0[0]), .b(b[25]), .bin(arrdiv32_fs472_or0[0]), .fs_xor1(arrdiv32_fs473_xor1), .fs_or0(arrdiv32_fs473_or0));
  fs fs_arrdiv32_fs474_out(.a(arrdiv32_mux2to1428_xor0[0]), .b(b[26]), .bin(arrdiv32_fs473_or0[0]), .fs_xor1(arrdiv32_fs474_xor1), .fs_or0(arrdiv32_fs474_or0));
  fs fs_arrdiv32_fs475_out(.a(arrdiv32_mux2to1429_xor0[0]), .b(b[27]), .bin(arrdiv32_fs474_or0[0]), .fs_xor1(arrdiv32_fs475_xor1), .fs_or0(arrdiv32_fs475_or0));
  fs fs_arrdiv32_fs476_out(.a(arrdiv32_mux2to1430_xor0[0]), .b(b[28]), .bin(arrdiv32_fs475_or0[0]), .fs_xor1(arrdiv32_fs476_xor1), .fs_or0(arrdiv32_fs476_or0));
  fs fs_arrdiv32_fs477_out(.a(arrdiv32_mux2to1431_xor0[0]), .b(b[29]), .bin(arrdiv32_fs476_or0[0]), .fs_xor1(arrdiv32_fs477_xor1), .fs_or0(arrdiv32_fs477_or0));
  fs fs_arrdiv32_fs478_out(.a(arrdiv32_mux2to1432_xor0[0]), .b(b[30]), .bin(arrdiv32_fs477_or0[0]), .fs_xor1(arrdiv32_fs478_xor1), .fs_or0(arrdiv32_fs478_or0));
  fs fs_arrdiv32_fs479_out(.a(arrdiv32_mux2to1433_xor0[0]), .b(b[31]), .bin(arrdiv32_fs478_or0[0]), .fs_xor1(arrdiv32_fs479_xor1), .fs_or0(arrdiv32_fs479_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1434_out(.d0(arrdiv32_fs448_xor0[0]), .d1(a[17]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1434_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1435_out(.d0(arrdiv32_fs449_xor1[0]), .d1(arrdiv32_mux2to1403_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1435_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1436_out(.d0(arrdiv32_fs450_xor1[0]), .d1(arrdiv32_mux2to1404_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1436_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1437_out(.d0(arrdiv32_fs451_xor1[0]), .d1(arrdiv32_mux2to1405_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1437_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1438_out(.d0(arrdiv32_fs452_xor1[0]), .d1(arrdiv32_mux2to1406_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1438_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1439_out(.d0(arrdiv32_fs453_xor1[0]), .d1(arrdiv32_mux2to1407_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1439_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1440_out(.d0(arrdiv32_fs454_xor1[0]), .d1(arrdiv32_mux2to1408_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1440_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1441_out(.d0(arrdiv32_fs455_xor1[0]), .d1(arrdiv32_mux2to1409_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1441_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1442_out(.d0(arrdiv32_fs456_xor1[0]), .d1(arrdiv32_mux2to1410_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1442_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1443_out(.d0(arrdiv32_fs457_xor1[0]), .d1(arrdiv32_mux2to1411_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1443_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1444_out(.d0(arrdiv32_fs458_xor1[0]), .d1(arrdiv32_mux2to1412_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1444_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1445_out(.d0(arrdiv32_fs459_xor1[0]), .d1(arrdiv32_mux2to1413_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1445_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1446_out(.d0(arrdiv32_fs460_xor1[0]), .d1(arrdiv32_mux2to1414_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1446_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1447_out(.d0(arrdiv32_fs461_xor1[0]), .d1(arrdiv32_mux2to1415_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1447_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1448_out(.d0(arrdiv32_fs462_xor1[0]), .d1(arrdiv32_mux2to1416_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1448_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1449_out(.d0(arrdiv32_fs463_xor1[0]), .d1(arrdiv32_mux2to1417_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1449_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1450_out(.d0(arrdiv32_fs464_xor1[0]), .d1(arrdiv32_mux2to1418_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1450_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1451_out(.d0(arrdiv32_fs465_xor1[0]), .d1(arrdiv32_mux2to1419_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1451_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1452_out(.d0(arrdiv32_fs466_xor1[0]), .d1(arrdiv32_mux2to1420_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1452_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1453_out(.d0(arrdiv32_fs467_xor1[0]), .d1(arrdiv32_mux2to1421_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1453_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1454_out(.d0(arrdiv32_fs468_xor1[0]), .d1(arrdiv32_mux2to1422_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1454_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1455_out(.d0(arrdiv32_fs469_xor1[0]), .d1(arrdiv32_mux2to1423_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1455_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1456_out(.d0(arrdiv32_fs470_xor1[0]), .d1(arrdiv32_mux2to1424_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1456_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1457_out(.d0(arrdiv32_fs471_xor1[0]), .d1(arrdiv32_mux2to1425_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1457_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1458_out(.d0(arrdiv32_fs472_xor1[0]), .d1(arrdiv32_mux2to1426_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1458_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1459_out(.d0(arrdiv32_fs473_xor1[0]), .d1(arrdiv32_mux2to1427_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1459_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1460_out(.d0(arrdiv32_fs474_xor1[0]), .d1(arrdiv32_mux2to1428_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1460_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1461_out(.d0(arrdiv32_fs475_xor1[0]), .d1(arrdiv32_mux2to1429_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1461_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1462_out(.d0(arrdiv32_fs476_xor1[0]), .d1(arrdiv32_mux2to1430_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1462_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1463_out(.d0(arrdiv32_fs477_xor1[0]), .d1(arrdiv32_mux2to1431_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1463_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1464_out(.d0(arrdiv32_fs478_xor1[0]), .d1(arrdiv32_mux2to1432_xor0[0]), .sel(arrdiv32_fs479_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1464_xor0));
  not_gate not_gate_arrdiv32_not14(.a(arrdiv32_fs479_or0[0]), .out(arrdiv32_not14));
  fs fs_arrdiv32_fs480_out(.a(a[16]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs480_xor0), .fs_or0(arrdiv32_fs480_and0));
  fs fs_arrdiv32_fs481_out(.a(arrdiv32_mux2to1434_xor0[0]), .b(b[1]), .bin(arrdiv32_fs480_and0[0]), .fs_xor1(arrdiv32_fs481_xor1), .fs_or0(arrdiv32_fs481_or0));
  fs fs_arrdiv32_fs482_out(.a(arrdiv32_mux2to1435_xor0[0]), .b(b[2]), .bin(arrdiv32_fs481_or0[0]), .fs_xor1(arrdiv32_fs482_xor1), .fs_or0(arrdiv32_fs482_or0));
  fs fs_arrdiv32_fs483_out(.a(arrdiv32_mux2to1436_xor0[0]), .b(b[3]), .bin(arrdiv32_fs482_or0[0]), .fs_xor1(arrdiv32_fs483_xor1), .fs_or0(arrdiv32_fs483_or0));
  fs fs_arrdiv32_fs484_out(.a(arrdiv32_mux2to1437_xor0[0]), .b(b[4]), .bin(arrdiv32_fs483_or0[0]), .fs_xor1(arrdiv32_fs484_xor1), .fs_or0(arrdiv32_fs484_or0));
  fs fs_arrdiv32_fs485_out(.a(arrdiv32_mux2to1438_xor0[0]), .b(b[5]), .bin(arrdiv32_fs484_or0[0]), .fs_xor1(arrdiv32_fs485_xor1), .fs_or0(arrdiv32_fs485_or0));
  fs fs_arrdiv32_fs486_out(.a(arrdiv32_mux2to1439_xor0[0]), .b(b[6]), .bin(arrdiv32_fs485_or0[0]), .fs_xor1(arrdiv32_fs486_xor1), .fs_or0(arrdiv32_fs486_or0));
  fs fs_arrdiv32_fs487_out(.a(arrdiv32_mux2to1440_xor0[0]), .b(b[7]), .bin(arrdiv32_fs486_or0[0]), .fs_xor1(arrdiv32_fs487_xor1), .fs_or0(arrdiv32_fs487_or0));
  fs fs_arrdiv32_fs488_out(.a(arrdiv32_mux2to1441_xor0[0]), .b(b[8]), .bin(arrdiv32_fs487_or0[0]), .fs_xor1(arrdiv32_fs488_xor1), .fs_or0(arrdiv32_fs488_or0));
  fs fs_arrdiv32_fs489_out(.a(arrdiv32_mux2to1442_xor0[0]), .b(b[9]), .bin(arrdiv32_fs488_or0[0]), .fs_xor1(arrdiv32_fs489_xor1), .fs_or0(arrdiv32_fs489_or0));
  fs fs_arrdiv32_fs490_out(.a(arrdiv32_mux2to1443_xor0[0]), .b(b[10]), .bin(arrdiv32_fs489_or0[0]), .fs_xor1(arrdiv32_fs490_xor1), .fs_or0(arrdiv32_fs490_or0));
  fs fs_arrdiv32_fs491_out(.a(arrdiv32_mux2to1444_xor0[0]), .b(b[11]), .bin(arrdiv32_fs490_or0[0]), .fs_xor1(arrdiv32_fs491_xor1), .fs_or0(arrdiv32_fs491_or0));
  fs fs_arrdiv32_fs492_out(.a(arrdiv32_mux2to1445_xor0[0]), .b(b[12]), .bin(arrdiv32_fs491_or0[0]), .fs_xor1(arrdiv32_fs492_xor1), .fs_or0(arrdiv32_fs492_or0));
  fs fs_arrdiv32_fs493_out(.a(arrdiv32_mux2to1446_xor0[0]), .b(b[13]), .bin(arrdiv32_fs492_or0[0]), .fs_xor1(arrdiv32_fs493_xor1), .fs_or0(arrdiv32_fs493_or0));
  fs fs_arrdiv32_fs494_out(.a(arrdiv32_mux2to1447_xor0[0]), .b(b[14]), .bin(arrdiv32_fs493_or0[0]), .fs_xor1(arrdiv32_fs494_xor1), .fs_or0(arrdiv32_fs494_or0));
  fs fs_arrdiv32_fs495_out(.a(arrdiv32_mux2to1448_xor0[0]), .b(b[15]), .bin(arrdiv32_fs494_or0[0]), .fs_xor1(arrdiv32_fs495_xor1), .fs_or0(arrdiv32_fs495_or0));
  fs fs_arrdiv32_fs496_out(.a(arrdiv32_mux2to1449_xor0[0]), .b(b[16]), .bin(arrdiv32_fs495_or0[0]), .fs_xor1(arrdiv32_fs496_xor1), .fs_or0(arrdiv32_fs496_or0));
  fs fs_arrdiv32_fs497_out(.a(arrdiv32_mux2to1450_xor0[0]), .b(b[17]), .bin(arrdiv32_fs496_or0[0]), .fs_xor1(arrdiv32_fs497_xor1), .fs_or0(arrdiv32_fs497_or0));
  fs fs_arrdiv32_fs498_out(.a(arrdiv32_mux2to1451_xor0[0]), .b(b[18]), .bin(arrdiv32_fs497_or0[0]), .fs_xor1(arrdiv32_fs498_xor1), .fs_or0(arrdiv32_fs498_or0));
  fs fs_arrdiv32_fs499_out(.a(arrdiv32_mux2to1452_xor0[0]), .b(b[19]), .bin(arrdiv32_fs498_or0[0]), .fs_xor1(arrdiv32_fs499_xor1), .fs_or0(arrdiv32_fs499_or0));
  fs fs_arrdiv32_fs500_out(.a(arrdiv32_mux2to1453_xor0[0]), .b(b[20]), .bin(arrdiv32_fs499_or0[0]), .fs_xor1(arrdiv32_fs500_xor1), .fs_or0(arrdiv32_fs500_or0));
  fs fs_arrdiv32_fs501_out(.a(arrdiv32_mux2to1454_xor0[0]), .b(b[21]), .bin(arrdiv32_fs500_or0[0]), .fs_xor1(arrdiv32_fs501_xor1), .fs_or0(arrdiv32_fs501_or0));
  fs fs_arrdiv32_fs502_out(.a(arrdiv32_mux2to1455_xor0[0]), .b(b[22]), .bin(arrdiv32_fs501_or0[0]), .fs_xor1(arrdiv32_fs502_xor1), .fs_or0(arrdiv32_fs502_or0));
  fs fs_arrdiv32_fs503_out(.a(arrdiv32_mux2to1456_xor0[0]), .b(b[23]), .bin(arrdiv32_fs502_or0[0]), .fs_xor1(arrdiv32_fs503_xor1), .fs_or0(arrdiv32_fs503_or0));
  fs fs_arrdiv32_fs504_out(.a(arrdiv32_mux2to1457_xor0[0]), .b(b[24]), .bin(arrdiv32_fs503_or0[0]), .fs_xor1(arrdiv32_fs504_xor1), .fs_or0(arrdiv32_fs504_or0));
  fs fs_arrdiv32_fs505_out(.a(arrdiv32_mux2to1458_xor0[0]), .b(b[25]), .bin(arrdiv32_fs504_or0[0]), .fs_xor1(arrdiv32_fs505_xor1), .fs_or0(arrdiv32_fs505_or0));
  fs fs_arrdiv32_fs506_out(.a(arrdiv32_mux2to1459_xor0[0]), .b(b[26]), .bin(arrdiv32_fs505_or0[0]), .fs_xor1(arrdiv32_fs506_xor1), .fs_or0(arrdiv32_fs506_or0));
  fs fs_arrdiv32_fs507_out(.a(arrdiv32_mux2to1460_xor0[0]), .b(b[27]), .bin(arrdiv32_fs506_or0[0]), .fs_xor1(arrdiv32_fs507_xor1), .fs_or0(arrdiv32_fs507_or0));
  fs fs_arrdiv32_fs508_out(.a(arrdiv32_mux2to1461_xor0[0]), .b(b[28]), .bin(arrdiv32_fs507_or0[0]), .fs_xor1(arrdiv32_fs508_xor1), .fs_or0(arrdiv32_fs508_or0));
  fs fs_arrdiv32_fs509_out(.a(arrdiv32_mux2to1462_xor0[0]), .b(b[29]), .bin(arrdiv32_fs508_or0[0]), .fs_xor1(arrdiv32_fs509_xor1), .fs_or0(arrdiv32_fs509_or0));
  fs fs_arrdiv32_fs510_out(.a(arrdiv32_mux2to1463_xor0[0]), .b(b[30]), .bin(arrdiv32_fs509_or0[0]), .fs_xor1(arrdiv32_fs510_xor1), .fs_or0(arrdiv32_fs510_or0));
  fs fs_arrdiv32_fs511_out(.a(arrdiv32_mux2to1464_xor0[0]), .b(b[31]), .bin(arrdiv32_fs510_or0[0]), .fs_xor1(arrdiv32_fs511_xor1), .fs_or0(arrdiv32_fs511_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1465_out(.d0(arrdiv32_fs480_xor0[0]), .d1(a[16]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1465_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1466_out(.d0(arrdiv32_fs481_xor1[0]), .d1(arrdiv32_mux2to1434_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1466_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1467_out(.d0(arrdiv32_fs482_xor1[0]), .d1(arrdiv32_mux2to1435_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1467_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1468_out(.d0(arrdiv32_fs483_xor1[0]), .d1(arrdiv32_mux2to1436_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1468_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1469_out(.d0(arrdiv32_fs484_xor1[0]), .d1(arrdiv32_mux2to1437_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1469_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1470_out(.d0(arrdiv32_fs485_xor1[0]), .d1(arrdiv32_mux2to1438_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1470_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1471_out(.d0(arrdiv32_fs486_xor1[0]), .d1(arrdiv32_mux2to1439_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1471_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1472_out(.d0(arrdiv32_fs487_xor1[0]), .d1(arrdiv32_mux2to1440_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1472_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1473_out(.d0(arrdiv32_fs488_xor1[0]), .d1(arrdiv32_mux2to1441_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1473_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1474_out(.d0(arrdiv32_fs489_xor1[0]), .d1(arrdiv32_mux2to1442_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1474_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1475_out(.d0(arrdiv32_fs490_xor1[0]), .d1(arrdiv32_mux2to1443_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1475_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1476_out(.d0(arrdiv32_fs491_xor1[0]), .d1(arrdiv32_mux2to1444_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1476_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1477_out(.d0(arrdiv32_fs492_xor1[0]), .d1(arrdiv32_mux2to1445_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1477_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1478_out(.d0(arrdiv32_fs493_xor1[0]), .d1(arrdiv32_mux2to1446_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1478_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1479_out(.d0(arrdiv32_fs494_xor1[0]), .d1(arrdiv32_mux2to1447_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1479_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1480_out(.d0(arrdiv32_fs495_xor1[0]), .d1(arrdiv32_mux2to1448_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1480_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1481_out(.d0(arrdiv32_fs496_xor1[0]), .d1(arrdiv32_mux2to1449_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1481_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1482_out(.d0(arrdiv32_fs497_xor1[0]), .d1(arrdiv32_mux2to1450_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1482_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1483_out(.d0(arrdiv32_fs498_xor1[0]), .d1(arrdiv32_mux2to1451_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1483_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1484_out(.d0(arrdiv32_fs499_xor1[0]), .d1(arrdiv32_mux2to1452_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1484_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1485_out(.d0(arrdiv32_fs500_xor1[0]), .d1(arrdiv32_mux2to1453_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1485_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1486_out(.d0(arrdiv32_fs501_xor1[0]), .d1(arrdiv32_mux2to1454_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1486_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1487_out(.d0(arrdiv32_fs502_xor1[0]), .d1(arrdiv32_mux2to1455_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1487_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1488_out(.d0(arrdiv32_fs503_xor1[0]), .d1(arrdiv32_mux2to1456_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1488_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1489_out(.d0(arrdiv32_fs504_xor1[0]), .d1(arrdiv32_mux2to1457_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1489_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1490_out(.d0(arrdiv32_fs505_xor1[0]), .d1(arrdiv32_mux2to1458_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1490_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1491_out(.d0(arrdiv32_fs506_xor1[0]), .d1(arrdiv32_mux2to1459_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1491_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1492_out(.d0(arrdiv32_fs507_xor1[0]), .d1(arrdiv32_mux2to1460_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1492_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1493_out(.d0(arrdiv32_fs508_xor1[0]), .d1(arrdiv32_mux2to1461_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1493_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1494_out(.d0(arrdiv32_fs509_xor1[0]), .d1(arrdiv32_mux2to1462_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1494_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1495_out(.d0(arrdiv32_fs510_xor1[0]), .d1(arrdiv32_mux2to1463_xor0[0]), .sel(arrdiv32_fs511_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1495_xor0));
  not_gate not_gate_arrdiv32_not15(.a(arrdiv32_fs511_or0[0]), .out(arrdiv32_not15));
  fs fs_arrdiv32_fs512_out(.a(a[15]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs512_xor0), .fs_or0(arrdiv32_fs512_and0));
  fs fs_arrdiv32_fs513_out(.a(arrdiv32_mux2to1465_xor0[0]), .b(b[1]), .bin(arrdiv32_fs512_and0[0]), .fs_xor1(arrdiv32_fs513_xor1), .fs_or0(arrdiv32_fs513_or0));
  fs fs_arrdiv32_fs514_out(.a(arrdiv32_mux2to1466_xor0[0]), .b(b[2]), .bin(arrdiv32_fs513_or0[0]), .fs_xor1(arrdiv32_fs514_xor1), .fs_or0(arrdiv32_fs514_or0));
  fs fs_arrdiv32_fs515_out(.a(arrdiv32_mux2to1467_xor0[0]), .b(b[3]), .bin(arrdiv32_fs514_or0[0]), .fs_xor1(arrdiv32_fs515_xor1), .fs_or0(arrdiv32_fs515_or0));
  fs fs_arrdiv32_fs516_out(.a(arrdiv32_mux2to1468_xor0[0]), .b(b[4]), .bin(arrdiv32_fs515_or0[0]), .fs_xor1(arrdiv32_fs516_xor1), .fs_or0(arrdiv32_fs516_or0));
  fs fs_arrdiv32_fs517_out(.a(arrdiv32_mux2to1469_xor0[0]), .b(b[5]), .bin(arrdiv32_fs516_or0[0]), .fs_xor1(arrdiv32_fs517_xor1), .fs_or0(arrdiv32_fs517_or0));
  fs fs_arrdiv32_fs518_out(.a(arrdiv32_mux2to1470_xor0[0]), .b(b[6]), .bin(arrdiv32_fs517_or0[0]), .fs_xor1(arrdiv32_fs518_xor1), .fs_or0(arrdiv32_fs518_or0));
  fs fs_arrdiv32_fs519_out(.a(arrdiv32_mux2to1471_xor0[0]), .b(b[7]), .bin(arrdiv32_fs518_or0[0]), .fs_xor1(arrdiv32_fs519_xor1), .fs_or0(arrdiv32_fs519_or0));
  fs fs_arrdiv32_fs520_out(.a(arrdiv32_mux2to1472_xor0[0]), .b(b[8]), .bin(arrdiv32_fs519_or0[0]), .fs_xor1(arrdiv32_fs520_xor1), .fs_or0(arrdiv32_fs520_or0));
  fs fs_arrdiv32_fs521_out(.a(arrdiv32_mux2to1473_xor0[0]), .b(b[9]), .bin(arrdiv32_fs520_or0[0]), .fs_xor1(arrdiv32_fs521_xor1), .fs_or0(arrdiv32_fs521_or0));
  fs fs_arrdiv32_fs522_out(.a(arrdiv32_mux2to1474_xor0[0]), .b(b[10]), .bin(arrdiv32_fs521_or0[0]), .fs_xor1(arrdiv32_fs522_xor1), .fs_or0(arrdiv32_fs522_or0));
  fs fs_arrdiv32_fs523_out(.a(arrdiv32_mux2to1475_xor0[0]), .b(b[11]), .bin(arrdiv32_fs522_or0[0]), .fs_xor1(arrdiv32_fs523_xor1), .fs_or0(arrdiv32_fs523_or0));
  fs fs_arrdiv32_fs524_out(.a(arrdiv32_mux2to1476_xor0[0]), .b(b[12]), .bin(arrdiv32_fs523_or0[0]), .fs_xor1(arrdiv32_fs524_xor1), .fs_or0(arrdiv32_fs524_or0));
  fs fs_arrdiv32_fs525_out(.a(arrdiv32_mux2to1477_xor0[0]), .b(b[13]), .bin(arrdiv32_fs524_or0[0]), .fs_xor1(arrdiv32_fs525_xor1), .fs_or0(arrdiv32_fs525_or0));
  fs fs_arrdiv32_fs526_out(.a(arrdiv32_mux2to1478_xor0[0]), .b(b[14]), .bin(arrdiv32_fs525_or0[0]), .fs_xor1(arrdiv32_fs526_xor1), .fs_or0(arrdiv32_fs526_or0));
  fs fs_arrdiv32_fs527_out(.a(arrdiv32_mux2to1479_xor0[0]), .b(b[15]), .bin(arrdiv32_fs526_or0[0]), .fs_xor1(arrdiv32_fs527_xor1), .fs_or0(arrdiv32_fs527_or0));
  fs fs_arrdiv32_fs528_out(.a(arrdiv32_mux2to1480_xor0[0]), .b(b[16]), .bin(arrdiv32_fs527_or0[0]), .fs_xor1(arrdiv32_fs528_xor1), .fs_or0(arrdiv32_fs528_or0));
  fs fs_arrdiv32_fs529_out(.a(arrdiv32_mux2to1481_xor0[0]), .b(b[17]), .bin(arrdiv32_fs528_or0[0]), .fs_xor1(arrdiv32_fs529_xor1), .fs_or0(arrdiv32_fs529_or0));
  fs fs_arrdiv32_fs530_out(.a(arrdiv32_mux2to1482_xor0[0]), .b(b[18]), .bin(arrdiv32_fs529_or0[0]), .fs_xor1(arrdiv32_fs530_xor1), .fs_or0(arrdiv32_fs530_or0));
  fs fs_arrdiv32_fs531_out(.a(arrdiv32_mux2to1483_xor0[0]), .b(b[19]), .bin(arrdiv32_fs530_or0[0]), .fs_xor1(arrdiv32_fs531_xor1), .fs_or0(arrdiv32_fs531_or0));
  fs fs_arrdiv32_fs532_out(.a(arrdiv32_mux2to1484_xor0[0]), .b(b[20]), .bin(arrdiv32_fs531_or0[0]), .fs_xor1(arrdiv32_fs532_xor1), .fs_or0(arrdiv32_fs532_or0));
  fs fs_arrdiv32_fs533_out(.a(arrdiv32_mux2to1485_xor0[0]), .b(b[21]), .bin(arrdiv32_fs532_or0[0]), .fs_xor1(arrdiv32_fs533_xor1), .fs_or0(arrdiv32_fs533_or0));
  fs fs_arrdiv32_fs534_out(.a(arrdiv32_mux2to1486_xor0[0]), .b(b[22]), .bin(arrdiv32_fs533_or0[0]), .fs_xor1(arrdiv32_fs534_xor1), .fs_or0(arrdiv32_fs534_or0));
  fs fs_arrdiv32_fs535_out(.a(arrdiv32_mux2to1487_xor0[0]), .b(b[23]), .bin(arrdiv32_fs534_or0[0]), .fs_xor1(arrdiv32_fs535_xor1), .fs_or0(arrdiv32_fs535_or0));
  fs fs_arrdiv32_fs536_out(.a(arrdiv32_mux2to1488_xor0[0]), .b(b[24]), .bin(arrdiv32_fs535_or0[0]), .fs_xor1(arrdiv32_fs536_xor1), .fs_or0(arrdiv32_fs536_or0));
  fs fs_arrdiv32_fs537_out(.a(arrdiv32_mux2to1489_xor0[0]), .b(b[25]), .bin(arrdiv32_fs536_or0[0]), .fs_xor1(arrdiv32_fs537_xor1), .fs_or0(arrdiv32_fs537_or0));
  fs fs_arrdiv32_fs538_out(.a(arrdiv32_mux2to1490_xor0[0]), .b(b[26]), .bin(arrdiv32_fs537_or0[0]), .fs_xor1(arrdiv32_fs538_xor1), .fs_or0(arrdiv32_fs538_or0));
  fs fs_arrdiv32_fs539_out(.a(arrdiv32_mux2to1491_xor0[0]), .b(b[27]), .bin(arrdiv32_fs538_or0[0]), .fs_xor1(arrdiv32_fs539_xor1), .fs_or0(arrdiv32_fs539_or0));
  fs fs_arrdiv32_fs540_out(.a(arrdiv32_mux2to1492_xor0[0]), .b(b[28]), .bin(arrdiv32_fs539_or0[0]), .fs_xor1(arrdiv32_fs540_xor1), .fs_or0(arrdiv32_fs540_or0));
  fs fs_arrdiv32_fs541_out(.a(arrdiv32_mux2to1493_xor0[0]), .b(b[29]), .bin(arrdiv32_fs540_or0[0]), .fs_xor1(arrdiv32_fs541_xor1), .fs_or0(arrdiv32_fs541_or0));
  fs fs_arrdiv32_fs542_out(.a(arrdiv32_mux2to1494_xor0[0]), .b(b[30]), .bin(arrdiv32_fs541_or0[0]), .fs_xor1(arrdiv32_fs542_xor1), .fs_or0(arrdiv32_fs542_or0));
  fs fs_arrdiv32_fs543_out(.a(arrdiv32_mux2to1495_xor0[0]), .b(b[31]), .bin(arrdiv32_fs542_or0[0]), .fs_xor1(arrdiv32_fs543_xor1), .fs_or0(arrdiv32_fs543_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1496_out(.d0(arrdiv32_fs512_xor0[0]), .d1(a[15]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1496_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1497_out(.d0(arrdiv32_fs513_xor1[0]), .d1(arrdiv32_mux2to1465_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1497_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1498_out(.d0(arrdiv32_fs514_xor1[0]), .d1(arrdiv32_mux2to1466_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1498_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1499_out(.d0(arrdiv32_fs515_xor1[0]), .d1(arrdiv32_mux2to1467_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1499_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1500_out(.d0(arrdiv32_fs516_xor1[0]), .d1(arrdiv32_mux2to1468_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1500_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1501_out(.d0(arrdiv32_fs517_xor1[0]), .d1(arrdiv32_mux2to1469_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1501_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1502_out(.d0(arrdiv32_fs518_xor1[0]), .d1(arrdiv32_mux2to1470_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1502_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1503_out(.d0(arrdiv32_fs519_xor1[0]), .d1(arrdiv32_mux2to1471_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1503_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1504_out(.d0(arrdiv32_fs520_xor1[0]), .d1(arrdiv32_mux2to1472_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1504_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1505_out(.d0(arrdiv32_fs521_xor1[0]), .d1(arrdiv32_mux2to1473_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1505_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1506_out(.d0(arrdiv32_fs522_xor1[0]), .d1(arrdiv32_mux2to1474_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1506_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1507_out(.d0(arrdiv32_fs523_xor1[0]), .d1(arrdiv32_mux2to1475_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1507_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1508_out(.d0(arrdiv32_fs524_xor1[0]), .d1(arrdiv32_mux2to1476_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1508_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1509_out(.d0(arrdiv32_fs525_xor1[0]), .d1(arrdiv32_mux2to1477_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1509_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1510_out(.d0(arrdiv32_fs526_xor1[0]), .d1(arrdiv32_mux2to1478_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1510_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1511_out(.d0(arrdiv32_fs527_xor1[0]), .d1(arrdiv32_mux2to1479_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1511_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1512_out(.d0(arrdiv32_fs528_xor1[0]), .d1(arrdiv32_mux2to1480_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1512_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1513_out(.d0(arrdiv32_fs529_xor1[0]), .d1(arrdiv32_mux2to1481_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1513_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1514_out(.d0(arrdiv32_fs530_xor1[0]), .d1(arrdiv32_mux2to1482_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1514_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1515_out(.d0(arrdiv32_fs531_xor1[0]), .d1(arrdiv32_mux2to1483_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1515_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1516_out(.d0(arrdiv32_fs532_xor1[0]), .d1(arrdiv32_mux2to1484_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1516_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1517_out(.d0(arrdiv32_fs533_xor1[0]), .d1(arrdiv32_mux2to1485_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1517_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1518_out(.d0(arrdiv32_fs534_xor1[0]), .d1(arrdiv32_mux2to1486_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1518_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1519_out(.d0(arrdiv32_fs535_xor1[0]), .d1(arrdiv32_mux2to1487_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1519_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1520_out(.d0(arrdiv32_fs536_xor1[0]), .d1(arrdiv32_mux2to1488_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1520_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1521_out(.d0(arrdiv32_fs537_xor1[0]), .d1(arrdiv32_mux2to1489_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1521_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1522_out(.d0(arrdiv32_fs538_xor1[0]), .d1(arrdiv32_mux2to1490_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1522_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1523_out(.d0(arrdiv32_fs539_xor1[0]), .d1(arrdiv32_mux2to1491_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1523_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1524_out(.d0(arrdiv32_fs540_xor1[0]), .d1(arrdiv32_mux2to1492_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1524_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1525_out(.d0(arrdiv32_fs541_xor1[0]), .d1(arrdiv32_mux2to1493_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1525_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1526_out(.d0(arrdiv32_fs542_xor1[0]), .d1(arrdiv32_mux2to1494_xor0[0]), .sel(arrdiv32_fs543_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1526_xor0));
  not_gate not_gate_arrdiv32_not16(.a(arrdiv32_fs543_or0[0]), .out(arrdiv32_not16));
  fs fs_arrdiv32_fs544_out(.a(a[14]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs544_xor0), .fs_or0(arrdiv32_fs544_and0));
  fs fs_arrdiv32_fs545_out(.a(arrdiv32_mux2to1496_xor0[0]), .b(b[1]), .bin(arrdiv32_fs544_and0[0]), .fs_xor1(arrdiv32_fs545_xor1), .fs_or0(arrdiv32_fs545_or0));
  fs fs_arrdiv32_fs546_out(.a(arrdiv32_mux2to1497_xor0[0]), .b(b[2]), .bin(arrdiv32_fs545_or0[0]), .fs_xor1(arrdiv32_fs546_xor1), .fs_or0(arrdiv32_fs546_or0));
  fs fs_arrdiv32_fs547_out(.a(arrdiv32_mux2to1498_xor0[0]), .b(b[3]), .bin(arrdiv32_fs546_or0[0]), .fs_xor1(arrdiv32_fs547_xor1), .fs_or0(arrdiv32_fs547_or0));
  fs fs_arrdiv32_fs548_out(.a(arrdiv32_mux2to1499_xor0[0]), .b(b[4]), .bin(arrdiv32_fs547_or0[0]), .fs_xor1(arrdiv32_fs548_xor1), .fs_or0(arrdiv32_fs548_or0));
  fs fs_arrdiv32_fs549_out(.a(arrdiv32_mux2to1500_xor0[0]), .b(b[5]), .bin(arrdiv32_fs548_or0[0]), .fs_xor1(arrdiv32_fs549_xor1), .fs_or0(arrdiv32_fs549_or0));
  fs fs_arrdiv32_fs550_out(.a(arrdiv32_mux2to1501_xor0[0]), .b(b[6]), .bin(arrdiv32_fs549_or0[0]), .fs_xor1(arrdiv32_fs550_xor1), .fs_or0(arrdiv32_fs550_or0));
  fs fs_arrdiv32_fs551_out(.a(arrdiv32_mux2to1502_xor0[0]), .b(b[7]), .bin(arrdiv32_fs550_or0[0]), .fs_xor1(arrdiv32_fs551_xor1), .fs_or0(arrdiv32_fs551_or0));
  fs fs_arrdiv32_fs552_out(.a(arrdiv32_mux2to1503_xor0[0]), .b(b[8]), .bin(arrdiv32_fs551_or0[0]), .fs_xor1(arrdiv32_fs552_xor1), .fs_or0(arrdiv32_fs552_or0));
  fs fs_arrdiv32_fs553_out(.a(arrdiv32_mux2to1504_xor0[0]), .b(b[9]), .bin(arrdiv32_fs552_or0[0]), .fs_xor1(arrdiv32_fs553_xor1), .fs_or0(arrdiv32_fs553_or0));
  fs fs_arrdiv32_fs554_out(.a(arrdiv32_mux2to1505_xor0[0]), .b(b[10]), .bin(arrdiv32_fs553_or0[0]), .fs_xor1(arrdiv32_fs554_xor1), .fs_or0(arrdiv32_fs554_or0));
  fs fs_arrdiv32_fs555_out(.a(arrdiv32_mux2to1506_xor0[0]), .b(b[11]), .bin(arrdiv32_fs554_or0[0]), .fs_xor1(arrdiv32_fs555_xor1), .fs_or0(arrdiv32_fs555_or0));
  fs fs_arrdiv32_fs556_out(.a(arrdiv32_mux2to1507_xor0[0]), .b(b[12]), .bin(arrdiv32_fs555_or0[0]), .fs_xor1(arrdiv32_fs556_xor1), .fs_or0(arrdiv32_fs556_or0));
  fs fs_arrdiv32_fs557_out(.a(arrdiv32_mux2to1508_xor0[0]), .b(b[13]), .bin(arrdiv32_fs556_or0[0]), .fs_xor1(arrdiv32_fs557_xor1), .fs_or0(arrdiv32_fs557_or0));
  fs fs_arrdiv32_fs558_out(.a(arrdiv32_mux2to1509_xor0[0]), .b(b[14]), .bin(arrdiv32_fs557_or0[0]), .fs_xor1(arrdiv32_fs558_xor1), .fs_or0(arrdiv32_fs558_or0));
  fs fs_arrdiv32_fs559_out(.a(arrdiv32_mux2to1510_xor0[0]), .b(b[15]), .bin(arrdiv32_fs558_or0[0]), .fs_xor1(arrdiv32_fs559_xor1), .fs_or0(arrdiv32_fs559_or0));
  fs fs_arrdiv32_fs560_out(.a(arrdiv32_mux2to1511_xor0[0]), .b(b[16]), .bin(arrdiv32_fs559_or0[0]), .fs_xor1(arrdiv32_fs560_xor1), .fs_or0(arrdiv32_fs560_or0));
  fs fs_arrdiv32_fs561_out(.a(arrdiv32_mux2to1512_xor0[0]), .b(b[17]), .bin(arrdiv32_fs560_or0[0]), .fs_xor1(arrdiv32_fs561_xor1), .fs_or0(arrdiv32_fs561_or0));
  fs fs_arrdiv32_fs562_out(.a(arrdiv32_mux2to1513_xor0[0]), .b(b[18]), .bin(arrdiv32_fs561_or0[0]), .fs_xor1(arrdiv32_fs562_xor1), .fs_or0(arrdiv32_fs562_or0));
  fs fs_arrdiv32_fs563_out(.a(arrdiv32_mux2to1514_xor0[0]), .b(b[19]), .bin(arrdiv32_fs562_or0[0]), .fs_xor1(arrdiv32_fs563_xor1), .fs_or0(arrdiv32_fs563_or0));
  fs fs_arrdiv32_fs564_out(.a(arrdiv32_mux2to1515_xor0[0]), .b(b[20]), .bin(arrdiv32_fs563_or0[0]), .fs_xor1(arrdiv32_fs564_xor1), .fs_or0(arrdiv32_fs564_or0));
  fs fs_arrdiv32_fs565_out(.a(arrdiv32_mux2to1516_xor0[0]), .b(b[21]), .bin(arrdiv32_fs564_or0[0]), .fs_xor1(arrdiv32_fs565_xor1), .fs_or0(arrdiv32_fs565_or0));
  fs fs_arrdiv32_fs566_out(.a(arrdiv32_mux2to1517_xor0[0]), .b(b[22]), .bin(arrdiv32_fs565_or0[0]), .fs_xor1(arrdiv32_fs566_xor1), .fs_or0(arrdiv32_fs566_or0));
  fs fs_arrdiv32_fs567_out(.a(arrdiv32_mux2to1518_xor0[0]), .b(b[23]), .bin(arrdiv32_fs566_or0[0]), .fs_xor1(arrdiv32_fs567_xor1), .fs_or0(arrdiv32_fs567_or0));
  fs fs_arrdiv32_fs568_out(.a(arrdiv32_mux2to1519_xor0[0]), .b(b[24]), .bin(arrdiv32_fs567_or0[0]), .fs_xor1(arrdiv32_fs568_xor1), .fs_or0(arrdiv32_fs568_or0));
  fs fs_arrdiv32_fs569_out(.a(arrdiv32_mux2to1520_xor0[0]), .b(b[25]), .bin(arrdiv32_fs568_or0[0]), .fs_xor1(arrdiv32_fs569_xor1), .fs_or0(arrdiv32_fs569_or0));
  fs fs_arrdiv32_fs570_out(.a(arrdiv32_mux2to1521_xor0[0]), .b(b[26]), .bin(arrdiv32_fs569_or0[0]), .fs_xor1(arrdiv32_fs570_xor1), .fs_or0(arrdiv32_fs570_or0));
  fs fs_arrdiv32_fs571_out(.a(arrdiv32_mux2to1522_xor0[0]), .b(b[27]), .bin(arrdiv32_fs570_or0[0]), .fs_xor1(arrdiv32_fs571_xor1), .fs_or0(arrdiv32_fs571_or0));
  fs fs_arrdiv32_fs572_out(.a(arrdiv32_mux2to1523_xor0[0]), .b(b[28]), .bin(arrdiv32_fs571_or0[0]), .fs_xor1(arrdiv32_fs572_xor1), .fs_or0(arrdiv32_fs572_or0));
  fs fs_arrdiv32_fs573_out(.a(arrdiv32_mux2to1524_xor0[0]), .b(b[29]), .bin(arrdiv32_fs572_or0[0]), .fs_xor1(arrdiv32_fs573_xor1), .fs_or0(arrdiv32_fs573_or0));
  fs fs_arrdiv32_fs574_out(.a(arrdiv32_mux2to1525_xor0[0]), .b(b[30]), .bin(arrdiv32_fs573_or0[0]), .fs_xor1(arrdiv32_fs574_xor1), .fs_or0(arrdiv32_fs574_or0));
  fs fs_arrdiv32_fs575_out(.a(arrdiv32_mux2to1526_xor0[0]), .b(b[31]), .bin(arrdiv32_fs574_or0[0]), .fs_xor1(arrdiv32_fs575_xor1), .fs_or0(arrdiv32_fs575_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1527_out(.d0(arrdiv32_fs544_xor0[0]), .d1(a[14]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1527_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1528_out(.d0(arrdiv32_fs545_xor1[0]), .d1(arrdiv32_mux2to1496_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1528_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1529_out(.d0(arrdiv32_fs546_xor1[0]), .d1(arrdiv32_mux2to1497_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1529_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1530_out(.d0(arrdiv32_fs547_xor1[0]), .d1(arrdiv32_mux2to1498_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1530_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1531_out(.d0(arrdiv32_fs548_xor1[0]), .d1(arrdiv32_mux2to1499_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1531_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1532_out(.d0(arrdiv32_fs549_xor1[0]), .d1(arrdiv32_mux2to1500_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1532_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1533_out(.d0(arrdiv32_fs550_xor1[0]), .d1(arrdiv32_mux2to1501_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1533_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1534_out(.d0(arrdiv32_fs551_xor1[0]), .d1(arrdiv32_mux2to1502_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1534_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1535_out(.d0(arrdiv32_fs552_xor1[0]), .d1(arrdiv32_mux2to1503_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1535_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1536_out(.d0(arrdiv32_fs553_xor1[0]), .d1(arrdiv32_mux2to1504_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1536_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1537_out(.d0(arrdiv32_fs554_xor1[0]), .d1(arrdiv32_mux2to1505_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1537_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1538_out(.d0(arrdiv32_fs555_xor1[0]), .d1(arrdiv32_mux2to1506_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1538_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1539_out(.d0(arrdiv32_fs556_xor1[0]), .d1(arrdiv32_mux2to1507_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1539_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1540_out(.d0(arrdiv32_fs557_xor1[0]), .d1(arrdiv32_mux2to1508_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1540_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1541_out(.d0(arrdiv32_fs558_xor1[0]), .d1(arrdiv32_mux2to1509_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1541_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1542_out(.d0(arrdiv32_fs559_xor1[0]), .d1(arrdiv32_mux2to1510_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1542_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1543_out(.d0(arrdiv32_fs560_xor1[0]), .d1(arrdiv32_mux2to1511_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1543_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1544_out(.d0(arrdiv32_fs561_xor1[0]), .d1(arrdiv32_mux2to1512_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1544_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1545_out(.d0(arrdiv32_fs562_xor1[0]), .d1(arrdiv32_mux2to1513_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1545_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1546_out(.d0(arrdiv32_fs563_xor1[0]), .d1(arrdiv32_mux2to1514_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1546_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1547_out(.d0(arrdiv32_fs564_xor1[0]), .d1(arrdiv32_mux2to1515_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1547_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1548_out(.d0(arrdiv32_fs565_xor1[0]), .d1(arrdiv32_mux2to1516_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1548_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1549_out(.d0(arrdiv32_fs566_xor1[0]), .d1(arrdiv32_mux2to1517_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1549_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1550_out(.d0(arrdiv32_fs567_xor1[0]), .d1(arrdiv32_mux2to1518_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1550_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1551_out(.d0(arrdiv32_fs568_xor1[0]), .d1(arrdiv32_mux2to1519_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1551_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1552_out(.d0(arrdiv32_fs569_xor1[0]), .d1(arrdiv32_mux2to1520_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1552_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1553_out(.d0(arrdiv32_fs570_xor1[0]), .d1(arrdiv32_mux2to1521_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1553_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1554_out(.d0(arrdiv32_fs571_xor1[0]), .d1(arrdiv32_mux2to1522_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1554_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1555_out(.d0(arrdiv32_fs572_xor1[0]), .d1(arrdiv32_mux2to1523_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1555_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1556_out(.d0(arrdiv32_fs573_xor1[0]), .d1(arrdiv32_mux2to1524_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1556_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1557_out(.d0(arrdiv32_fs574_xor1[0]), .d1(arrdiv32_mux2to1525_xor0[0]), .sel(arrdiv32_fs575_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1557_xor0));
  not_gate not_gate_arrdiv32_not17(.a(arrdiv32_fs575_or0[0]), .out(arrdiv32_not17));
  fs fs_arrdiv32_fs576_out(.a(a[13]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs576_xor0), .fs_or0(arrdiv32_fs576_and0));
  fs fs_arrdiv32_fs577_out(.a(arrdiv32_mux2to1527_xor0[0]), .b(b[1]), .bin(arrdiv32_fs576_and0[0]), .fs_xor1(arrdiv32_fs577_xor1), .fs_or0(arrdiv32_fs577_or0));
  fs fs_arrdiv32_fs578_out(.a(arrdiv32_mux2to1528_xor0[0]), .b(b[2]), .bin(arrdiv32_fs577_or0[0]), .fs_xor1(arrdiv32_fs578_xor1), .fs_or0(arrdiv32_fs578_or0));
  fs fs_arrdiv32_fs579_out(.a(arrdiv32_mux2to1529_xor0[0]), .b(b[3]), .bin(arrdiv32_fs578_or0[0]), .fs_xor1(arrdiv32_fs579_xor1), .fs_or0(arrdiv32_fs579_or0));
  fs fs_arrdiv32_fs580_out(.a(arrdiv32_mux2to1530_xor0[0]), .b(b[4]), .bin(arrdiv32_fs579_or0[0]), .fs_xor1(arrdiv32_fs580_xor1), .fs_or0(arrdiv32_fs580_or0));
  fs fs_arrdiv32_fs581_out(.a(arrdiv32_mux2to1531_xor0[0]), .b(b[5]), .bin(arrdiv32_fs580_or0[0]), .fs_xor1(arrdiv32_fs581_xor1), .fs_or0(arrdiv32_fs581_or0));
  fs fs_arrdiv32_fs582_out(.a(arrdiv32_mux2to1532_xor0[0]), .b(b[6]), .bin(arrdiv32_fs581_or0[0]), .fs_xor1(arrdiv32_fs582_xor1), .fs_or0(arrdiv32_fs582_or0));
  fs fs_arrdiv32_fs583_out(.a(arrdiv32_mux2to1533_xor0[0]), .b(b[7]), .bin(arrdiv32_fs582_or0[0]), .fs_xor1(arrdiv32_fs583_xor1), .fs_or0(arrdiv32_fs583_or0));
  fs fs_arrdiv32_fs584_out(.a(arrdiv32_mux2to1534_xor0[0]), .b(b[8]), .bin(arrdiv32_fs583_or0[0]), .fs_xor1(arrdiv32_fs584_xor1), .fs_or0(arrdiv32_fs584_or0));
  fs fs_arrdiv32_fs585_out(.a(arrdiv32_mux2to1535_xor0[0]), .b(b[9]), .bin(arrdiv32_fs584_or0[0]), .fs_xor1(arrdiv32_fs585_xor1), .fs_or0(arrdiv32_fs585_or0));
  fs fs_arrdiv32_fs586_out(.a(arrdiv32_mux2to1536_xor0[0]), .b(b[10]), .bin(arrdiv32_fs585_or0[0]), .fs_xor1(arrdiv32_fs586_xor1), .fs_or0(arrdiv32_fs586_or0));
  fs fs_arrdiv32_fs587_out(.a(arrdiv32_mux2to1537_xor0[0]), .b(b[11]), .bin(arrdiv32_fs586_or0[0]), .fs_xor1(arrdiv32_fs587_xor1), .fs_or0(arrdiv32_fs587_or0));
  fs fs_arrdiv32_fs588_out(.a(arrdiv32_mux2to1538_xor0[0]), .b(b[12]), .bin(arrdiv32_fs587_or0[0]), .fs_xor1(arrdiv32_fs588_xor1), .fs_or0(arrdiv32_fs588_or0));
  fs fs_arrdiv32_fs589_out(.a(arrdiv32_mux2to1539_xor0[0]), .b(b[13]), .bin(arrdiv32_fs588_or0[0]), .fs_xor1(arrdiv32_fs589_xor1), .fs_or0(arrdiv32_fs589_or0));
  fs fs_arrdiv32_fs590_out(.a(arrdiv32_mux2to1540_xor0[0]), .b(b[14]), .bin(arrdiv32_fs589_or0[0]), .fs_xor1(arrdiv32_fs590_xor1), .fs_or0(arrdiv32_fs590_or0));
  fs fs_arrdiv32_fs591_out(.a(arrdiv32_mux2to1541_xor0[0]), .b(b[15]), .bin(arrdiv32_fs590_or0[0]), .fs_xor1(arrdiv32_fs591_xor1), .fs_or0(arrdiv32_fs591_or0));
  fs fs_arrdiv32_fs592_out(.a(arrdiv32_mux2to1542_xor0[0]), .b(b[16]), .bin(arrdiv32_fs591_or0[0]), .fs_xor1(arrdiv32_fs592_xor1), .fs_or0(arrdiv32_fs592_or0));
  fs fs_arrdiv32_fs593_out(.a(arrdiv32_mux2to1543_xor0[0]), .b(b[17]), .bin(arrdiv32_fs592_or0[0]), .fs_xor1(arrdiv32_fs593_xor1), .fs_or0(arrdiv32_fs593_or0));
  fs fs_arrdiv32_fs594_out(.a(arrdiv32_mux2to1544_xor0[0]), .b(b[18]), .bin(arrdiv32_fs593_or0[0]), .fs_xor1(arrdiv32_fs594_xor1), .fs_or0(arrdiv32_fs594_or0));
  fs fs_arrdiv32_fs595_out(.a(arrdiv32_mux2to1545_xor0[0]), .b(b[19]), .bin(arrdiv32_fs594_or0[0]), .fs_xor1(arrdiv32_fs595_xor1), .fs_or0(arrdiv32_fs595_or0));
  fs fs_arrdiv32_fs596_out(.a(arrdiv32_mux2to1546_xor0[0]), .b(b[20]), .bin(arrdiv32_fs595_or0[0]), .fs_xor1(arrdiv32_fs596_xor1), .fs_or0(arrdiv32_fs596_or0));
  fs fs_arrdiv32_fs597_out(.a(arrdiv32_mux2to1547_xor0[0]), .b(b[21]), .bin(arrdiv32_fs596_or0[0]), .fs_xor1(arrdiv32_fs597_xor1), .fs_or0(arrdiv32_fs597_or0));
  fs fs_arrdiv32_fs598_out(.a(arrdiv32_mux2to1548_xor0[0]), .b(b[22]), .bin(arrdiv32_fs597_or0[0]), .fs_xor1(arrdiv32_fs598_xor1), .fs_or0(arrdiv32_fs598_or0));
  fs fs_arrdiv32_fs599_out(.a(arrdiv32_mux2to1549_xor0[0]), .b(b[23]), .bin(arrdiv32_fs598_or0[0]), .fs_xor1(arrdiv32_fs599_xor1), .fs_or0(arrdiv32_fs599_or0));
  fs fs_arrdiv32_fs600_out(.a(arrdiv32_mux2to1550_xor0[0]), .b(b[24]), .bin(arrdiv32_fs599_or0[0]), .fs_xor1(arrdiv32_fs600_xor1), .fs_or0(arrdiv32_fs600_or0));
  fs fs_arrdiv32_fs601_out(.a(arrdiv32_mux2to1551_xor0[0]), .b(b[25]), .bin(arrdiv32_fs600_or0[0]), .fs_xor1(arrdiv32_fs601_xor1), .fs_or0(arrdiv32_fs601_or0));
  fs fs_arrdiv32_fs602_out(.a(arrdiv32_mux2to1552_xor0[0]), .b(b[26]), .bin(arrdiv32_fs601_or0[0]), .fs_xor1(arrdiv32_fs602_xor1), .fs_or0(arrdiv32_fs602_or0));
  fs fs_arrdiv32_fs603_out(.a(arrdiv32_mux2to1553_xor0[0]), .b(b[27]), .bin(arrdiv32_fs602_or0[0]), .fs_xor1(arrdiv32_fs603_xor1), .fs_or0(arrdiv32_fs603_or0));
  fs fs_arrdiv32_fs604_out(.a(arrdiv32_mux2to1554_xor0[0]), .b(b[28]), .bin(arrdiv32_fs603_or0[0]), .fs_xor1(arrdiv32_fs604_xor1), .fs_or0(arrdiv32_fs604_or0));
  fs fs_arrdiv32_fs605_out(.a(arrdiv32_mux2to1555_xor0[0]), .b(b[29]), .bin(arrdiv32_fs604_or0[0]), .fs_xor1(arrdiv32_fs605_xor1), .fs_or0(arrdiv32_fs605_or0));
  fs fs_arrdiv32_fs606_out(.a(arrdiv32_mux2to1556_xor0[0]), .b(b[30]), .bin(arrdiv32_fs605_or0[0]), .fs_xor1(arrdiv32_fs606_xor1), .fs_or0(arrdiv32_fs606_or0));
  fs fs_arrdiv32_fs607_out(.a(arrdiv32_mux2to1557_xor0[0]), .b(b[31]), .bin(arrdiv32_fs606_or0[0]), .fs_xor1(arrdiv32_fs607_xor1), .fs_or0(arrdiv32_fs607_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1558_out(.d0(arrdiv32_fs576_xor0[0]), .d1(a[13]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1558_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1559_out(.d0(arrdiv32_fs577_xor1[0]), .d1(arrdiv32_mux2to1527_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1559_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1560_out(.d0(arrdiv32_fs578_xor1[0]), .d1(arrdiv32_mux2to1528_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1560_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1561_out(.d0(arrdiv32_fs579_xor1[0]), .d1(arrdiv32_mux2to1529_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1561_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1562_out(.d0(arrdiv32_fs580_xor1[0]), .d1(arrdiv32_mux2to1530_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1562_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1563_out(.d0(arrdiv32_fs581_xor1[0]), .d1(arrdiv32_mux2to1531_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1563_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1564_out(.d0(arrdiv32_fs582_xor1[0]), .d1(arrdiv32_mux2to1532_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1564_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1565_out(.d0(arrdiv32_fs583_xor1[0]), .d1(arrdiv32_mux2to1533_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1565_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1566_out(.d0(arrdiv32_fs584_xor1[0]), .d1(arrdiv32_mux2to1534_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1566_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1567_out(.d0(arrdiv32_fs585_xor1[0]), .d1(arrdiv32_mux2to1535_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1567_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1568_out(.d0(arrdiv32_fs586_xor1[0]), .d1(arrdiv32_mux2to1536_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1568_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1569_out(.d0(arrdiv32_fs587_xor1[0]), .d1(arrdiv32_mux2to1537_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1569_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1570_out(.d0(arrdiv32_fs588_xor1[0]), .d1(arrdiv32_mux2to1538_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1570_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1571_out(.d0(arrdiv32_fs589_xor1[0]), .d1(arrdiv32_mux2to1539_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1571_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1572_out(.d0(arrdiv32_fs590_xor1[0]), .d1(arrdiv32_mux2to1540_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1572_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1573_out(.d0(arrdiv32_fs591_xor1[0]), .d1(arrdiv32_mux2to1541_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1573_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1574_out(.d0(arrdiv32_fs592_xor1[0]), .d1(arrdiv32_mux2to1542_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1574_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1575_out(.d0(arrdiv32_fs593_xor1[0]), .d1(arrdiv32_mux2to1543_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1575_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1576_out(.d0(arrdiv32_fs594_xor1[0]), .d1(arrdiv32_mux2to1544_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1576_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1577_out(.d0(arrdiv32_fs595_xor1[0]), .d1(arrdiv32_mux2to1545_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1577_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1578_out(.d0(arrdiv32_fs596_xor1[0]), .d1(arrdiv32_mux2to1546_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1578_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1579_out(.d0(arrdiv32_fs597_xor1[0]), .d1(arrdiv32_mux2to1547_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1579_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1580_out(.d0(arrdiv32_fs598_xor1[0]), .d1(arrdiv32_mux2to1548_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1580_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1581_out(.d0(arrdiv32_fs599_xor1[0]), .d1(arrdiv32_mux2to1549_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1581_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1582_out(.d0(arrdiv32_fs600_xor1[0]), .d1(arrdiv32_mux2to1550_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1582_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1583_out(.d0(arrdiv32_fs601_xor1[0]), .d1(arrdiv32_mux2to1551_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1583_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1584_out(.d0(arrdiv32_fs602_xor1[0]), .d1(arrdiv32_mux2to1552_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1584_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1585_out(.d0(arrdiv32_fs603_xor1[0]), .d1(arrdiv32_mux2to1553_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1585_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1586_out(.d0(arrdiv32_fs604_xor1[0]), .d1(arrdiv32_mux2to1554_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1586_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1587_out(.d0(arrdiv32_fs605_xor1[0]), .d1(arrdiv32_mux2to1555_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1587_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1588_out(.d0(arrdiv32_fs606_xor1[0]), .d1(arrdiv32_mux2to1556_xor0[0]), .sel(arrdiv32_fs607_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1588_xor0));
  not_gate not_gate_arrdiv32_not18(.a(arrdiv32_fs607_or0[0]), .out(arrdiv32_not18));
  fs fs_arrdiv32_fs608_out(.a(a[12]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs608_xor0), .fs_or0(arrdiv32_fs608_and0));
  fs fs_arrdiv32_fs609_out(.a(arrdiv32_mux2to1558_xor0[0]), .b(b[1]), .bin(arrdiv32_fs608_and0[0]), .fs_xor1(arrdiv32_fs609_xor1), .fs_or0(arrdiv32_fs609_or0));
  fs fs_arrdiv32_fs610_out(.a(arrdiv32_mux2to1559_xor0[0]), .b(b[2]), .bin(arrdiv32_fs609_or0[0]), .fs_xor1(arrdiv32_fs610_xor1), .fs_or0(arrdiv32_fs610_or0));
  fs fs_arrdiv32_fs611_out(.a(arrdiv32_mux2to1560_xor0[0]), .b(b[3]), .bin(arrdiv32_fs610_or0[0]), .fs_xor1(arrdiv32_fs611_xor1), .fs_or0(arrdiv32_fs611_or0));
  fs fs_arrdiv32_fs612_out(.a(arrdiv32_mux2to1561_xor0[0]), .b(b[4]), .bin(arrdiv32_fs611_or0[0]), .fs_xor1(arrdiv32_fs612_xor1), .fs_or0(arrdiv32_fs612_or0));
  fs fs_arrdiv32_fs613_out(.a(arrdiv32_mux2to1562_xor0[0]), .b(b[5]), .bin(arrdiv32_fs612_or0[0]), .fs_xor1(arrdiv32_fs613_xor1), .fs_or0(arrdiv32_fs613_or0));
  fs fs_arrdiv32_fs614_out(.a(arrdiv32_mux2to1563_xor0[0]), .b(b[6]), .bin(arrdiv32_fs613_or0[0]), .fs_xor1(arrdiv32_fs614_xor1), .fs_or0(arrdiv32_fs614_or0));
  fs fs_arrdiv32_fs615_out(.a(arrdiv32_mux2to1564_xor0[0]), .b(b[7]), .bin(arrdiv32_fs614_or0[0]), .fs_xor1(arrdiv32_fs615_xor1), .fs_or0(arrdiv32_fs615_or0));
  fs fs_arrdiv32_fs616_out(.a(arrdiv32_mux2to1565_xor0[0]), .b(b[8]), .bin(arrdiv32_fs615_or0[0]), .fs_xor1(arrdiv32_fs616_xor1), .fs_or0(arrdiv32_fs616_or0));
  fs fs_arrdiv32_fs617_out(.a(arrdiv32_mux2to1566_xor0[0]), .b(b[9]), .bin(arrdiv32_fs616_or0[0]), .fs_xor1(arrdiv32_fs617_xor1), .fs_or0(arrdiv32_fs617_or0));
  fs fs_arrdiv32_fs618_out(.a(arrdiv32_mux2to1567_xor0[0]), .b(b[10]), .bin(arrdiv32_fs617_or0[0]), .fs_xor1(arrdiv32_fs618_xor1), .fs_or0(arrdiv32_fs618_or0));
  fs fs_arrdiv32_fs619_out(.a(arrdiv32_mux2to1568_xor0[0]), .b(b[11]), .bin(arrdiv32_fs618_or0[0]), .fs_xor1(arrdiv32_fs619_xor1), .fs_or0(arrdiv32_fs619_or0));
  fs fs_arrdiv32_fs620_out(.a(arrdiv32_mux2to1569_xor0[0]), .b(b[12]), .bin(arrdiv32_fs619_or0[0]), .fs_xor1(arrdiv32_fs620_xor1), .fs_or0(arrdiv32_fs620_or0));
  fs fs_arrdiv32_fs621_out(.a(arrdiv32_mux2to1570_xor0[0]), .b(b[13]), .bin(arrdiv32_fs620_or0[0]), .fs_xor1(arrdiv32_fs621_xor1), .fs_or0(arrdiv32_fs621_or0));
  fs fs_arrdiv32_fs622_out(.a(arrdiv32_mux2to1571_xor0[0]), .b(b[14]), .bin(arrdiv32_fs621_or0[0]), .fs_xor1(arrdiv32_fs622_xor1), .fs_or0(arrdiv32_fs622_or0));
  fs fs_arrdiv32_fs623_out(.a(arrdiv32_mux2to1572_xor0[0]), .b(b[15]), .bin(arrdiv32_fs622_or0[0]), .fs_xor1(arrdiv32_fs623_xor1), .fs_or0(arrdiv32_fs623_or0));
  fs fs_arrdiv32_fs624_out(.a(arrdiv32_mux2to1573_xor0[0]), .b(b[16]), .bin(arrdiv32_fs623_or0[0]), .fs_xor1(arrdiv32_fs624_xor1), .fs_or0(arrdiv32_fs624_or0));
  fs fs_arrdiv32_fs625_out(.a(arrdiv32_mux2to1574_xor0[0]), .b(b[17]), .bin(arrdiv32_fs624_or0[0]), .fs_xor1(arrdiv32_fs625_xor1), .fs_or0(arrdiv32_fs625_or0));
  fs fs_arrdiv32_fs626_out(.a(arrdiv32_mux2to1575_xor0[0]), .b(b[18]), .bin(arrdiv32_fs625_or0[0]), .fs_xor1(arrdiv32_fs626_xor1), .fs_or0(arrdiv32_fs626_or0));
  fs fs_arrdiv32_fs627_out(.a(arrdiv32_mux2to1576_xor0[0]), .b(b[19]), .bin(arrdiv32_fs626_or0[0]), .fs_xor1(arrdiv32_fs627_xor1), .fs_or0(arrdiv32_fs627_or0));
  fs fs_arrdiv32_fs628_out(.a(arrdiv32_mux2to1577_xor0[0]), .b(b[20]), .bin(arrdiv32_fs627_or0[0]), .fs_xor1(arrdiv32_fs628_xor1), .fs_or0(arrdiv32_fs628_or0));
  fs fs_arrdiv32_fs629_out(.a(arrdiv32_mux2to1578_xor0[0]), .b(b[21]), .bin(arrdiv32_fs628_or0[0]), .fs_xor1(arrdiv32_fs629_xor1), .fs_or0(arrdiv32_fs629_or0));
  fs fs_arrdiv32_fs630_out(.a(arrdiv32_mux2to1579_xor0[0]), .b(b[22]), .bin(arrdiv32_fs629_or0[0]), .fs_xor1(arrdiv32_fs630_xor1), .fs_or0(arrdiv32_fs630_or0));
  fs fs_arrdiv32_fs631_out(.a(arrdiv32_mux2to1580_xor0[0]), .b(b[23]), .bin(arrdiv32_fs630_or0[0]), .fs_xor1(arrdiv32_fs631_xor1), .fs_or0(arrdiv32_fs631_or0));
  fs fs_arrdiv32_fs632_out(.a(arrdiv32_mux2to1581_xor0[0]), .b(b[24]), .bin(arrdiv32_fs631_or0[0]), .fs_xor1(arrdiv32_fs632_xor1), .fs_or0(arrdiv32_fs632_or0));
  fs fs_arrdiv32_fs633_out(.a(arrdiv32_mux2to1582_xor0[0]), .b(b[25]), .bin(arrdiv32_fs632_or0[0]), .fs_xor1(arrdiv32_fs633_xor1), .fs_or0(arrdiv32_fs633_or0));
  fs fs_arrdiv32_fs634_out(.a(arrdiv32_mux2to1583_xor0[0]), .b(b[26]), .bin(arrdiv32_fs633_or0[0]), .fs_xor1(arrdiv32_fs634_xor1), .fs_or0(arrdiv32_fs634_or0));
  fs fs_arrdiv32_fs635_out(.a(arrdiv32_mux2to1584_xor0[0]), .b(b[27]), .bin(arrdiv32_fs634_or0[0]), .fs_xor1(arrdiv32_fs635_xor1), .fs_or0(arrdiv32_fs635_or0));
  fs fs_arrdiv32_fs636_out(.a(arrdiv32_mux2to1585_xor0[0]), .b(b[28]), .bin(arrdiv32_fs635_or0[0]), .fs_xor1(arrdiv32_fs636_xor1), .fs_or0(arrdiv32_fs636_or0));
  fs fs_arrdiv32_fs637_out(.a(arrdiv32_mux2to1586_xor0[0]), .b(b[29]), .bin(arrdiv32_fs636_or0[0]), .fs_xor1(arrdiv32_fs637_xor1), .fs_or0(arrdiv32_fs637_or0));
  fs fs_arrdiv32_fs638_out(.a(arrdiv32_mux2to1587_xor0[0]), .b(b[30]), .bin(arrdiv32_fs637_or0[0]), .fs_xor1(arrdiv32_fs638_xor1), .fs_or0(arrdiv32_fs638_or0));
  fs fs_arrdiv32_fs639_out(.a(arrdiv32_mux2to1588_xor0[0]), .b(b[31]), .bin(arrdiv32_fs638_or0[0]), .fs_xor1(arrdiv32_fs639_xor1), .fs_or0(arrdiv32_fs639_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1589_out(.d0(arrdiv32_fs608_xor0[0]), .d1(a[12]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1589_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1590_out(.d0(arrdiv32_fs609_xor1[0]), .d1(arrdiv32_mux2to1558_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1590_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1591_out(.d0(arrdiv32_fs610_xor1[0]), .d1(arrdiv32_mux2to1559_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1591_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1592_out(.d0(arrdiv32_fs611_xor1[0]), .d1(arrdiv32_mux2to1560_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1592_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1593_out(.d0(arrdiv32_fs612_xor1[0]), .d1(arrdiv32_mux2to1561_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1593_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1594_out(.d0(arrdiv32_fs613_xor1[0]), .d1(arrdiv32_mux2to1562_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1594_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1595_out(.d0(arrdiv32_fs614_xor1[0]), .d1(arrdiv32_mux2to1563_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1595_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1596_out(.d0(arrdiv32_fs615_xor1[0]), .d1(arrdiv32_mux2to1564_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1596_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1597_out(.d0(arrdiv32_fs616_xor1[0]), .d1(arrdiv32_mux2to1565_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1597_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1598_out(.d0(arrdiv32_fs617_xor1[0]), .d1(arrdiv32_mux2to1566_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1598_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1599_out(.d0(arrdiv32_fs618_xor1[0]), .d1(arrdiv32_mux2to1567_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1599_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1600_out(.d0(arrdiv32_fs619_xor1[0]), .d1(arrdiv32_mux2to1568_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1600_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1601_out(.d0(arrdiv32_fs620_xor1[0]), .d1(arrdiv32_mux2to1569_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1601_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1602_out(.d0(arrdiv32_fs621_xor1[0]), .d1(arrdiv32_mux2to1570_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1602_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1603_out(.d0(arrdiv32_fs622_xor1[0]), .d1(arrdiv32_mux2to1571_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1603_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1604_out(.d0(arrdiv32_fs623_xor1[0]), .d1(arrdiv32_mux2to1572_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1604_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1605_out(.d0(arrdiv32_fs624_xor1[0]), .d1(arrdiv32_mux2to1573_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1605_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1606_out(.d0(arrdiv32_fs625_xor1[0]), .d1(arrdiv32_mux2to1574_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1606_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1607_out(.d0(arrdiv32_fs626_xor1[0]), .d1(arrdiv32_mux2to1575_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1607_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1608_out(.d0(arrdiv32_fs627_xor1[0]), .d1(arrdiv32_mux2to1576_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1608_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1609_out(.d0(arrdiv32_fs628_xor1[0]), .d1(arrdiv32_mux2to1577_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1609_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1610_out(.d0(arrdiv32_fs629_xor1[0]), .d1(arrdiv32_mux2to1578_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1610_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1611_out(.d0(arrdiv32_fs630_xor1[0]), .d1(arrdiv32_mux2to1579_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1611_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1612_out(.d0(arrdiv32_fs631_xor1[0]), .d1(arrdiv32_mux2to1580_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1612_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1613_out(.d0(arrdiv32_fs632_xor1[0]), .d1(arrdiv32_mux2to1581_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1613_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1614_out(.d0(arrdiv32_fs633_xor1[0]), .d1(arrdiv32_mux2to1582_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1614_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1615_out(.d0(arrdiv32_fs634_xor1[0]), .d1(arrdiv32_mux2to1583_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1615_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1616_out(.d0(arrdiv32_fs635_xor1[0]), .d1(arrdiv32_mux2to1584_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1616_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1617_out(.d0(arrdiv32_fs636_xor1[0]), .d1(arrdiv32_mux2to1585_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1617_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1618_out(.d0(arrdiv32_fs637_xor1[0]), .d1(arrdiv32_mux2to1586_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1618_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1619_out(.d0(arrdiv32_fs638_xor1[0]), .d1(arrdiv32_mux2to1587_xor0[0]), .sel(arrdiv32_fs639_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1619_xor0));
  not_gate not_gate_arrdiv32_not19(.a(arrdiv32_fs639_or0[0]), .out(arrdiv32_not19));
  fs fs_arrdiv32_fs640_out(.a(a[11]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs640_xor0), .fs_or0(arrdiv32_fs640_and0));
  fs fs_arrdiv32_fs641_out(.a(arrdiv32_mux2to1589_xor0[0]), .b(b[1]), .bin(arrdiv32_fs640_and0[0]), .fs_xor1(arrdiv32_fs641_xor1), .fs_or0(arrdiv32_fs641_or0));
  fs fs_arrdiv32_fs642_out(.a(arrdiv32_mux2to1590_xor0[0]), .b(b[2]), .bin(arrdiv32_fs641_or0[0]), .fs_xor1(arrdiv32_fs642_xor1), .fs_or0(arrdiv32_fs642_or0));
  fs fs_arrdiv32_fs643_out(.a(arrdiv32_mux2to1591_xor0[0]), .b(b[3]), .bin(arrdiv32_fs642_or0[0]), .fs_xor1(arrdiv32_fs643_xor1), .fs_or0(arrdiv32_fs643_or0));
  fs fs_arrdiv32_fs644_out(.a(arrdiv32_mux2to1592_xor0[0]), .b(b[4]), .bin(arrdiv32_fs643_or0[0]), .fs_xor1(arrdiv32_fs644_xor1), .fs_or0(arrdiv32_fs644_or0));
  fs fs_arrdiv32_fs645_out(.a(arrdiv32_mux2to1593_xor0[0]), .b(b[5]), .bin(arrdiv32_fs644_or0[0]), .fs_xor1(arrdiv32_fs645_xor1), .fs_or0(arrdiv32_fs645_or0));
  fs fs_arrdiv32_fs646_out(.a(arrdiv32_mux2to1594_xor0[0]), .b(b[6]), .bin(arrdiv32_fs645_or0[0]), .fs_xor1(arrdiv32_fs646_xor1), .fs_or0(arrdiv32_fs646_or0));
  fs fs_arrdiv32_fs647_out(.a(arrdiv32_mux2to1595_xor0[0]), .b(b[7]), .bin(arrdiv32_fs646_or0[0]), .fs_xor1(arrdiv32_fs647_xor1), .fs_or0(arrdiv32_fs647_or0));
  fs fs_arrdiv32_fs648_out(.a(arrdiv32_mux2to1596_xor0[0]), .b(b[8]), .bin(arrdiv32_fs647_or0[0]), .fs_xor1(arrdiv32_fs648_xor1), .fs_or0(arrdiv32_fs648_or0));
  fs fs_arrdiv32_fs649_out(.a(arrdiv32_mux2to1597_xor0[0]), .b(b[9]), .bin(arrdiv32_fs648_or0[0]), .fs_xor1(arrdiv32_fs649_xor1), .fs_or0(arrdiv32_fs649_or0));
  fs fs_arrdiv32_fs650_out(.a(arrdiv32_mux2to1598_xor0[0]), .b(b[10]), .bin(arrdiv32_fs649_or0[0]), .fs_xor1(arrdiv32_fs650_xor1), .fs_or0(arrdiv32_fs650_or0));
  fs fs_arrdiv32_fs651_out(.a(arrdiv32_mux2to1599_xor0[0]), .b(b[11]), .bin(arrdiv32_fs650_or0[0]), .fs_xor1(arrdiv32_fs651_xor1), .fs_or0(arrdiv32_fs651_or0));
  fs fs_arrdiv32_fs652_out(.a(arrdiv32_mux2to1600_xor0[0]), .b(b[12]), .bin(arrdiv32_fs651_or0[0]), .fs_xor1(arrdiv32_fs652_xor1), .fs_or0(arrdiv32_fs652_or0));
  fs fs_arrdiv32_fs653_out(.a(arrdiv32_mux2to1601_xor0[0]), .b(b[13]), .bin(arrdiv32_fs652_or0[0]), .fs_xor1(arrdiv32_fs653_xor1), .fs_or0(arrdiv32_fs653_or0));
  fs fs_arrdiv32_fs654_out(.a(arrdiv32_mux2to1602_xor0[0]), .b(b[14]), .bin(arrdiv32_fs653_or0[0]), .fs_xor1(arrdiv32_fs654_xor1), .fs_or0(arrdiv32_fs654_or0));
  fs fs_arrdiv32_fs655_out(.a(arrdiv32_mux2to1603_xor0[0]), .b(b[15]), .bin(arrdiv32_fs654_or0[0]), .fs_xor1(arrdiv32_fs655_xor1), .fs_or0(arrdiv32_fs655_or0));
  fs fs_arrdiv32_fs656_out(.a(arrdiv32_mux2to1604_xor0[0]), .b(b[16]), .bin(arrdiv32_fs655_or0[0]), .fs_xor1(arrdiv32_fs656_xor1), .fs_or0(arrdiv32_fs656_or0));
  fs fs_arrdiv32_fs657_out(.a(arrdiv32_mux2to1605_xor0[0]), .b(b[17]), .bin(arrdiv32_fs656_or0[0]), .fs_xor1(arrdiv32_fs657_xor1), .fs_or0(arrdiv32_fs657_or0));
  fs fs_arrdiv32_fs658_out(.a(arrdiv32_mux2to1606_xor0[0]), .b(b[18]), .bin(arrdiv32_fs657_or0[0]), .fs_xor1(arrdiv32_fs658_xor1), .fs_or0(arrdiv32_fs658_or0));
  fs fs_arrdiv32_fs659_out(.a(arrdiv32_mux2to1607_xor0[0]), .b(b[19]), .bin(arrdiv32_fs658_or0[0]), .fs_xor1(arrdiv32_fs659_xor1), .fs_or0(arrdiv32_fs659_or0));
  fs fs_arrdiv32_fs660_out(.a(arrdiv32_mux2to1608_xor0[0]), .b(b[20]), .bin(arrdiv32_fs659_or0[0]), .fs_xor1(arrdiv32_fs660_xor1), .fs_or0(arrdiv32_fs660_or0));
  fs fs_arrdiv32_fs661_out(.a(arrdiv32_mux2to1609_xor0[0]), .b(b[21]), .bin(arrdiv32_fs660_or0[0]), .fs_xor1(arrdiv32_fs661_xor1), .fs_or0(arrdiv32_fs661_or0));
  fs fs_arrdiv32_fs662_out(.a(arrdiv32_mux2to1610_xor0[0]), .b(b[22]), .bin(arrdiv32_fs661_or0[0]), .fs_xor1(arrdiv32_fs662_xor1), .fs_or0(arrdiv32_fs662_or0));
  fs fs_arrdiv32_fs663_out(.a(arrdiv32_mux2to1611_xor0[0]), .b(b[23]), .bin(arrdiv32_fs662_or0[0]), .fs_xor1(arrdiv32_fs663_xor1), .fs_or0(arrdiv32_fs663_or0));
  fs fs_arrdiv32_fs664_out(.a(arrdiv32_mux2to1612_xor0[0]), .b(b[24]), .bin(arrdiv32_fs663_or0[0]), .fs_xor1(arrdiv32_fs664_xor1), .fs_or0(arrdiv32_fs664_or0));
  fs fs_arrdiv32_fs665_out(.a(arrdiv32_mux2to1613_xor0[0]), .b(b[25]), .bin(arrdiv32_fs664_or0[0]), .fs_xor1(arrdiv32_fs665_xor1), .fs_or0(arrdiv32_fs665_or0));
  fs fs_arrdiv32_fs666_out(.a(arrdiv32_mux2to1614_xor0[0]), .b(b[26]), .bin(arrdiv32_fs665_or0[0]), .fs_xor1(arrdiv32_fs666_xor1), .fs_or0(arrdiv32_fs666_or0));
  fs fs_arrdiv32_fs667_out(.a(arrdiv32_mux2to1615_xor0[0]), .b(b[27]), .bin(arrdiv32_fs666_or0[0]), .fs_xor1(arrdiv32_fs667_xor1), .fs_or0(arrdiv32_fs667_or0));
  fs fs_arrdiv32_fs668_out(.a(arrdiv32_mux2to1616_xor0[0]), .b(b[28]), .bin(arrdiv32_fs667_or0[0]), .fs_xor1(arrdiv32_fs668_xor1), .fs_or0(arrdiv32_fs668_or0));
  fs fs_arrdiv32_fs669_out(.a(arrdiv32_mux2to1617_xor0[0]), .b(b[29]), .bin(arrdiv32_fs668_or0[0]), .fs_xor1(arrdiv32_fs669_xor1), .fs_or0(arrdiv32_fs669_or0));
  fs fs_arrdiv32_fs670_out(.a(arrdiv32_mux2to1618_xor0[0]), .b(b[30]), .bin(arrdiv32_fs669_or0[0]), .fs_xor1(arrdiv32_fs670_xor1), .fs_or0(arrdiv32_fs670_or0));
  fs fs_arrdiv32_fs671_out(.a(arrdiv32_mux2to1619_xor0[0]), .b(b[31]), .bin(arrdiv32_fs670_or0[0]), .fs_xor1(arrdiv32_fs671_xor1), .fs_or0(arrdiv32_fs671_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1620_out(.d0(arrdiv32_fs640_xor0[0]), .d1(a[11]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1620_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1621_out(.d0(arrdiv32_fs641_xor1[0]), .d1(arrdiv32_mux2to1589_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1621_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1622_out(.d0(arrdiv32_fs642_xor1[0]), .d1(arrdiv32_mux2to1590_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1622_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1623_out(.d0(arrdiv32_fs643_xor1[0]), .d1(arrdiv32_mux2to1591_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1623_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1624_out(.d0(arrdiv32_fs644_xor1[0]), .d1(arrdiv32_mux2to1592_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1624_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1625_out(.d0(arrdiv32_fs645_xor1[0]), .d1(arrdiv32_mux2to1593_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1625_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1626_out(.d0(arrdiv32_fs646_xor1[0]), .d1(arrdiv32_mux2to1594_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1626_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1627_out(.d0(arrdiv32_fs647_xor1[0]), .d1(arrdiv32_mux2to1595_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1627_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1628_out(.d0(arrdiv32_fs648_xor1[0]), .d1(arrdiv32_mux2to1596_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1628_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1629_out(.d0(arrdiv32_fs649_xor1[0]), .d1(arrdiv32_mux2to1597_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1629_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1630_out(.d0(arrdiv32_fs650_xor1[0]), .d1(arrdiv32_mux2to1598_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1630_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1631_out(.d0(arrdiv32_fs651_xor1[0]), .d1(arrdiv32_mux2to1599_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1631_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1632_out(.d0(arrdiv32_fs652_xor1[0]), .d1(arrdiv32_mux2to1600_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1632_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1633_out(.d0(arrdiv32_fs653_xor1[0]), .d1(arrdiv32_mux2to1601_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1633_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1634_out(.d0(arrdiv32_fs654_xor1[0]), .d1(arrdiv32_mux2to1602_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1634_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1635_out(.d0(arrdiv32_fs655_xor1[0]), .d1(arrdiv32_mux2to1603_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1635_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1636_out(.d0(arrdiv32_fs656_xor1[0]), .d1(arrdiv32_mux2to1604_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1636_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1637_out(.d0(arrdiv32_fs657_xor1[0]), .d1(arrdiv32_mux2to1605_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1637_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1638_out(.d0(arrdiv32_fs658_xor1[0]), .d1(arrdiv32_mux2to1606_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1638_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1639_out(.d0(arrdiv32_fs659_xor1[0]), .d1(arrdiv32_mux2to1607_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1639_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1640_out(.d0(arrdiv32_fs660_xor1[0]), .d1(arrdiv32_mux2to1608_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1640_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1641_out(.d0(arrdiv32_fs661_xor1[0]), .d1(arrdiv32_mux2to1609_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1641_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1642_out(.d0(arrdiv32_fs662_xor1[0]), .d1(arrdiv32_mux2to1610_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1642_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1643_out(.d0(arrdiv32_fs663_xor1[0]), .d1(arrdiv32_mux2to1611_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1643_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1644_out(.d0(arrdiv32_fs664_xor1[0]), .d1(arrdiv32_mux2to1612_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1644_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1645_out(.d0(arrdiv32_fs665_xor1[0]), .d1(arrdiv32_mux2to1613_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1645_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1646_out(.d0(arrdiv32_fs666_xor1[0]), .d1(arrdiv32_mux2to1614_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1646_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1647_out(.d0(arrdiv32_fs667_xor1[0]), .d1(arrdiv32_mux2to1615_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1647_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1648_out(.d0(arrdiv32_fs668_xor1[0]), .d1(arrdiv32_mux2to1616_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1648_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1649_out(.d0(arrdiv32_fs669_xor1[0]), .d1(arrdiv32_mux2to1617_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1649_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1650_out(.d0(arrdiv32_fs670_xor1[0]), .d1(arrdiv32_mux2to1618_xor0[0]), .sel(arrdiv32_fs671_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1650_xor0));
  not_gate not_gate_arrdiv32_not20(.a(arrdiv32_fs671_or0[0]), .out(arrdiv32_not20));
  fs fs_arrdiv32_fs672_out(.a(a[10]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs672_xor0), .fs_or0(arrdiv32_fs672_and0));
  fs fs_arrdiv32_fs673_out(.a(arrdiv32_mux2to1620_xor0[0]), .b(b[1]), .bin(arrdiv32_fs672_and0[0]), .fs_xor1(arrdiv32_fs673_xor1), .fs_or0(arrdiv32_fs673_or0));
  fs fs_arrdiv32_fs674_out(.a(arrdiv32_mux2to1621_xor0[0]), .b(b[2]), .bin(arrdiv32_fs673_or0[0]), .fs_xor1(arrdiv32_fs674_xor1), .fs_or0(arrdiv32_fs674_or0));
  fs fs_arrdiv32_fs675_out(.a(arrdiv32_mux2to1622_xor0[0]), .b(b[3]), .bin(arrdiv32_fs674_or0[0]), .fs_xor1(arrdiv32_fs675_xor1), .fs_or0(arrdiv32_fs675_or0));
  fs fs_arrdiv32_fs676_out(.a(arrdiv32_mux2to1623_xor0[0]), .b(b[4]), .bin(arrdiv32_fs675_or0[0]), .fs_xor1(arrdiv32_fs676_xor1), .fs_or0(arrdiv32_fs676_or0));
  fs fs_arrdiv32_fs677_out(.a(arrdiv32_mux2to1624_xor0[0]), .b(b[5]), .bin(arrdiv32_fs676_or0[0]), .fs_xor1(arrdiv32_fs677_xor1), .fs_or0(arrdiv32_fs677_or0));
  fs fs_arrdiv32_fs678_out(.a(arrdiv32_mux2to1625_xor0[0]), .b(b[6]), .bin(arrdiv32_fs677_or0[0]), .fs_xor1(arrdiv32_fs678_xor1), .fs_or0(arrdiv32_fs678_or0));
  fs fs_arrdiv32_fs679_out(.a(arrdiv32_mux2to1626_xor0[0]), .b(b[7]), .bin(arrdiv32_fs678_or0[0]), .fs_xor1(arrdiv32_fs679_xor1), .fs_or0(arrdiv32_fs679_or0));
  fs fs_arrdiv32_fs680_out(.a(arrdiv32_mux2to1627_xor0[0]), .b(b[8]), .bin(arrdiv32_fs679_or0[0]), .fs_xor1(arrdiv32_fs680_xor1), .fs_or0(arrdiv32_fs680_or0));
  fs fs_arrdiv32_fs681_out(.a(arrdiv32_mux2to1628_xor0[0]), .b(b[9]), .bin(arrdiv32_fs680_or0[0]), .fs_xor1(arrdiv32_fs681_xor1), .fs_or0(arrdiv32_fs681_or0));
  fs fs_arrdiv32_fs682_out(.a(arrdiv32_mux2to1629_xor0[0]), .b(b[10]), .bin(arrdiv32_fs681_or0[0]), .fs_xor1(arrdiv32_fs682_xor1), .fs_or0(arrdiv32_fs682_or0));
  fs fs_arrdiv32_fs683_out(.a(arrdiv32_mux2to1630_xor0[0]), .b(b[11]), .bin(arrdiv32_fs682_or0[0]), .fs_xor1(arrdiv32_fs683_xor1), .fs_or0(arrdiv32_fs683_or0));
  fs fs_arrdiv32_fs684_out(.a(arrdiv32_mux2to1631_xor0[0]), .b(b[12]), .bin(arrdiv32_fs683_or0[0]), .fs_xor1(arrdiv32_fs684_xor1), .fs_or0(arrdiv32_fs684_or0));
  fs fs_arrdiv32_fs685_out(.a(arrdiv32_mux2to1632_xor0[0]), .b(b[13]), .bin(arrdiv32_fs684_or0[0]), .fs_xor1(arrdiv32_fs685_xor1), .fs_or0(arrdiv32_fs685_or0));
  fs fs_arrdiv32_fs686_out(.a(arrdiv32_mux2to1633_xor0[0]), .b(b[14]), .bin(arrdiv32_fs685_or0[0]), .fs_xor1(arrdiv32_fs686_xor1), .fs_or0(arrdiv32_fs686_or0));
  fs fs_arrdiv32_fs687_out(.a(arrdiv32_mux2to1634_xor0[0]), .b(b[15]), .bin(arrdiv32_fs686_or0[0]), .fs_xor1(arrdiv32_fs687_xor1), .fs_or0(arrdiv32_fs687_or0));
  fs fs_arrdiv32_fs688_out(.a(arrdiv32_mux2to1635_xor0[0]), .b(b[16]), .bin(arrdiv32_fs687_or0[0]), .fs_xor1(arrdiv32_fs688_xor1), .fs_or0(arrdiv32_fs688_or0));
  fs fs_arrdiv32_fs689_out(.a(arrdiv32_mux2to1636_xor0[0]), .b(b[17]), .bin(arrdiv32_fs688_or0[0]), .fs_xor1(arrdiv32_fs689_xor1), .fs_or0(arrdiv32_fs689_or0));
  fs fs_arrdiv32_fs690_out(.a(arrdiv32_mux2to1637_xor0[0]), .b(b[18]), .bin(arrdiv32_fs689_or0[0]), .fs_xor1(arrdiv32_fs690_xor1), .fs_or0(arrdiv32_fs690_or0));
  fs fs_arrdiv32_fs691_out(.a(arrdiv32_mux2to1638_xor0[0]), .b(b[19]), .bin(arrdiv32_fs690_or0[0]), .fs_xor1(arrdiv32_fs691_xor1), .fs_or0(arrdiv32_fs691_or0));
  fs fs_arrdiv32_fs692_out(.a(arrdiv32_mux2to1639_xor0[0]), .b(b[20]), .bin(arrdiv32_fs691_or0[0]), .fs_xor1(arrdiv32_fs692_xor1), .fs_or0(arrdiv32_fs692_or0));
  fs fs_arrdiv32_fs693_out(.a(arrdiv32_mux2to1640_xor0[0]), .b(b[21]), .bin(arrdiv32_fs692_or0[0]), .fs_xor1(arrdiv32_fs693_xor1), .fs_or0(arrdiv32_fs693_or0));
  fs fs_arrdiv32_fs694_out(.a(arrdiv32_mux2to1641_xor0[0]), .b(b[22]), .bin(arrdiv32_fs693_or0[0]), .fs_xor1(arrdiv32_fs694_xor1), .fs_or0(arrdiv32_fs694_or0));
  fs fs_arrdiv32_fs695_out(.a(arrdiv32_mux2to1642_xor0[0]), .b(b[23]), .bin(arrdiv32_fs694_or0[0]), .fs_xor1(arrdiv32_fs695_xor1), .fs_or0(arrdiv32_fs695_or0));
  fs fs_arrdiv32_fs696_out(.a(arrdiv32_mux2to1643_xor0[0]), .b(b[24]), .bin(arrdiv32_fs695_or0[0]), .fs_xor1(arrdiv32_fs696_xor1), .fs_or0(arrdiv32_fs696_or0));
  fs fs_arrdiv32_fs697_out(.a(arrdiv32_mux2to1644_xor0[0]), .b(b[25]), .bin(arrdiv32_fs696_or0[0]), .fs_xor1(arrdiv32_fs697_xor1), .fs_or0(arrdiv32_fs697_or0));
  fs fs_arrdiv32_fs698_out(.a(arrdiv32_mux2to1645_xor0[0]), .b(b[26]), .bin(arrdiv32_fs697_or0[0]), .fs_xor1(arrdiv32_fs698_xor1), .fs_or0(arrdiv32_fs698_or0));
  fs fs_arrdiv32_fs699_out(.a(arrdiv32_mux2to1646_xor0[0]), .b(b[27]), .bin(arrdiv32_fs698_or0[0]), .fs_xor1(arrdiv32_fs699_xor1), .fs_or0(arrdiv32_fs699_or0));
  fs fs_arrdiv32_fs700_out(.a(arrdiv32_mux2to1647_xor0[0]), .b(b[28]), .bin(arrdiv32_fs699_or0[0]), .fs_xor1(arrdiv32_fs700_xor1), .fs_or0(arrdiv32_fs700_or0));
  fs fs_arrdiv32_fs701_out(.a(arrdiv32_mux2to1648_xor0[0]), .b(b[29]), .bin(arrdiv32_fs700_or0[0]), .fs_xor1(arrdiv32_fs701_xor1), .fs_or0(arrdiv32_fs701_or0));
  fs fs_arrdiv32_fs702_out(.a(arrdiv32_mux2to1649_xor0[0]), .b(b[30]), .bin(arrdiv32_fs701_or0[0]), .fs_xor1(arrdiv32_fs702_xor1), .fs_or0(arrdiv32_fs702_or0));
  fs fs_arrdiv32_fs703_out(.a(arrdiv32_mux2to1650_xor0[0]), .b(b[31]), .bin(arrdiv32_fs702_or0[0]), .fs_xor1(arrdiv32_fs703_xor1), .fs_or0(arrdiv32_fs703_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1651_out(.d0(arrdiv32_fs672_xor0[0]), .d1(a[10]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1651_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1652_out(.d0(arrdiv32_fs673_xor1[0]), .d1(arrdiv32_mux2to1620_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1652_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1653_out(.d0(arrdiv32_fs674_xor1[0]), .d1(arrdiv32_mux2to1621_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1653_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1654_out(.d0(arrdiv32_fs675_xor1[0]), .d1(arrdiv32_mux2to1622_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1654_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1655_out(.d0(arrdiv32_fs676_xor1[0]), .d1(arrdiv32_mux2to1623_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1655_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1656_out(.d0(arrdiv32_fs677_xor1[0]), .d1(arrdiv32_mux2to1624_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1656_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1657_out(.d0(arrdiv32_fs678_xor1[0]), .d1(arrdiv32_mux2to1625_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1657_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1658_out(.d0(arrdiv32_fs679_xor1[0]), .d1(arrdiv32_mux2to1626_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1658_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1659_out(.d0(arrdiv32_fs680_xor1[0]), .d1(arrdiv32_mux2to1627_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1659_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1660_out(.d0(arrdiv32_fs681_xor1[0]), .d1(arrdiv32_mux2to1628_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1660_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1661_out(.d0(arrdiv32_fs682_xor1[0]), .d1(arrdiv32_mux2to1629_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1661_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1662_out(.d0(arrdiv32_fs683_xor1[0]), .d1(arrdiv32_mux2to1630_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1662_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1663_out(.d0(arrdiv32_fs684_xor1[0]), .d1(arrdiv32_mux2to1631_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1663_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1664_out(.d0(arrdiv32_fs685_xor1[0]), .d1(arrdiv32_mux2to1632_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1664_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1665_out(.d0(arrdiv32_fs686_xor1[0]), .d1(arrdiv32_mux2to1633_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1665_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1666_out(.d0(arrdiv32_fs687_xor1[0]), .d1(arrdiv32_mux2to1634_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1666_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1667_out(.d0(arrdiv32_fs688_xor1[0]), .d1(arrdiv32_mux2to1635_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1667_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1668_out(.d0(arrdiv32_fs689_xor1[0]), .d1(arrdiv32_mux2to1636_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1668_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1669_out(.d0(arrdiv32_fs690_xor1[0]), .d1(arrdiv32_mux2to1637_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1669_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1670_out(.d0(arrdiv32_fs691_xor1[0]), .d1(arrdiv32_mux2to1638_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1670_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1671_out(.d0(arrdiv32_fs692_xor1[0]), .d1(arrdiv32_mux2to1639_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1671_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1672_out(.d0(arrdiv32_fs693_xor1[0]), .d1(arrdiv32_mux2to1640_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1672_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1673_out(.d0(arrdiv32_fs694_xor1[0]), .d1(arrdiv32_mux2to1641_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1673_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1674_out(.d0(arrdiv32_fs695_xor1[0]), .d1(arrdiv32_mux2to1642_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1674_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1675_out(.d0(arrdiv32_fs696_xor1[0]), .d1(arrdiv32_mux2to1643_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1675_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1676_out(.d0(arrdiv32_fs697_xor1[0]), .d1(arrdiv32_mux2to1644_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1676_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1677_out(.d0(arrdiv32_fs698_xor1[0]), .d1(arrdiv32_mux2to1645_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1677_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1678_out(.d0(arrdiv32_fs699_xor1[0]), .d1(arrdiv32_mux2to1646_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1678_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1679_out(.d0(arrdiv32_fs700_xor1[0]), .d1(arrdiv32_mux2to1647_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1679_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1680_out(.d0(arrdiv32_fs701_xor1[0]), .d1(arrdiv32_mux2to1648_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1680_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1681_out(.d0(arrdiv32_fs702_xor1[0]), .d1(arrdiv32_mux2to1649_xor0[0]), .sel(arrdiv32_fs703_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1681_xor0));
  not_gate not_gate_arrdiv32_not21(.a(arrdiv32_fs703_or0[0]), .out(arrdiv32_not21));
  fs fs_arrdiv32_fs704_out(.a(a[9]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs704_xor0), .fs_or0(arrdiv32_fs704_and0));
  fs fs_arrdiv32_fs705_out(.a(arrdiv32_mux2to1651_xor0[0]), .b(b[1]), .bin(arrdiv32_fs704_and0[0]), .fs_xor1(arrdiv32_fs705_xor1), .fs_or0(arrdiv32_fs705_or0));
  fs fs_arrdiv32_fs706_out(.a(arrdiv32_mux2to1652_xor0[0]), .b(b[2]), .bin(arrdiv32_fs705_or0[0]), .fs_xor1(arrdiv32_fs706_xor1), .fs_or0(arrdiv32_fs706_or0));
  fs fs_arrdiv32_fs707_out(.a(arrdiv32_mux2to1653_xor0[0]), .b(b[3]), .bin(arrdiv32_fs706_or0[0]), .fs_xor1(arrdiv32_fs707_xor1), .fs_or0(arrdiv32_fs707_or0));
  fs fs_arrdiv32_fs708_out(.a(arrdiv32_mux2to1654_xor0[0]), .b(b[4]), .bin(arrdiv32_fs707_or0[0]), .fs_xor1(arrdiv32_fs708_xor1), .fs_or0(arrdiv32_fs708_or0));
  fs fs_arrdiv32_fs709_out(.a(arrdiv32_mux2to1655_xor0[0]), .b(b[5]), .bin(arrdiv32_fs708_or0[0]), .fs_xor1(arrdiv32_fs709_xor1), .fs_or0(arrdiv32_fs709_or0));
  fs fs_arrdiv32_fs710_out(.a(arrdiv32_mux2to1656_xor0[0]), .b(b[6]), .bin(arrdiv32_fs709_or0[0]), .fs_xor1(arrdiv32_fs710_xor1), .fs_or0(arrdiv32_fs710_or0));
  fs fs_arrdiv32_fs711_out(.a(arrdiv32_mux2to1657_xor0[0]), .b(b[7]), .bin(arrdiv32_fs710_or0[0]), .fs_xor1(arrdiv32_fs711_xor1), .fs_or0(arrdiv32_fs711_or0));
  fs fs_arrdiv32_fs712_out(.a(arrdiv32_mux2to1658_xor0[0]), .b(b[8]), .bin(arrdiv32_fs711_or0[0]), .fs_xor1(arrdiv32_fs712_xor1), .fs_or0(arrdiv32_fs712_or0));
  fs fs_arrdiv32_fs713_out(.a(arrdiv32_mux2to1659_xor0[0]), .b(b[9]), .bin(arrdiv32_fs712_or0[0]), .fs_xor1(arrdiv32_fs713_xor1), .fs_or0(arrdiv32_fs713_or0));
  fs fs_arrdiv32_fs714_out(.a(arrdiv32_mux2to1660_xor0[0]), .b(b[10]), .bin(arrdiv32_fs713_or0[0]), .fs_xor1(arrdiv32_fs714_xor1), .fs_or0(arrdiv32_fs714_or0));
  fs fs_arrdiv32_fs715_out(.a(arrdiv32_mux2to1661_xor0[0]), .b(b[11]), .bin(arrdiv32_fs714_or0[0]), .fs_xor1(arrdiv32_fs715_xor1), .fs_or0(arrdiv32_fs715_or0));
  fs fs_arrdiv32_fs716_out(.a(arrdiv32_mux2to1662_xor0[0]), .b(b[12]), .bin(arrdiv32_fs715_or0[0]), .fs_xor1(arrdiv32_fs716_xor1), .fs_or0(arrdiv32_fs716_or0));
  fs fs_arrdiv32_fs717_out(.a(arrdiv32_mux2to1663_xor0[0]), .b(b[13]), .bin(arrdiv32_fs716_or0[0]), .fs_xor1(arrdiv32_fs717_xor1), .fs_or0(arrdiv32_fs717_or0));
  fs fs_arrdiv32_fs718_out(.a(arrdiv32_mux2to1664_xor0[0]), .b(b[14]), .bin(arrdiv32_fs717_or0[0]), .fs_xor1(arrdiv32_fs718_xor1), .fs_or0(arrdiv32_fs718_or0));
  fs fs_arrdiv32_fs719_out(.a(arrdiv32_mux2to1665_xor0[0]), .b(b[15]), .bin(arrdiv32_fs718_or0[0]), .fs_xor1(arrdiv32_fs719_xor1), .fs_or0(arrdiv32_fs719_or0));
  fs fs_arrdiv32_fs720_out(.a(arrdiv32_mux2to1666_xor0[0]), .b(b[16]), .bin(arrdiv32_fs719_or0[0]), .fs_xor1(arrdiv32_fs720_xor1), .fs_or0(arrdiv32_fs720_or0));
  fs fs_arrdiv32_fs721_out(.a(arrdiv32_mux2to1667_xor0[0]), .b(b[17]), .bin(arrdiv32_fs720_or0[0]), .fs_xor1(arrdiv32_fs721_xor1), .fs_or0(arrdiv32_fs721_or0));
  fs fs_arrdiv32_fs722_out(.a(arrdiv32_mux2to1668_xor0[0]), .b(b[18]), .bin(arrdiv32_fs721_or0[0]), .fs_xor1(arrdiv32_fs722_xor1), .fs_or0(arrdiv32_fs722_or0));
  fs fs_arrdiv32_fs723_out(.a(arrdiv32_mux2to1669_xor0[0]), .b(b[19]), .bin(arrdiv32_fs722_or0[0]), .fs_xor1(arrdiv32_fs723_xor1), .fs_or0(arrdiv32_fs723_or0));
  fs fs_arrdiv32_fs724_out(.a(arrdiv32_mux2to1670_xor0[0]), .b(b[20]), .bin(arrdiv32_fs723_or0[0]), .fs_xor1(arrdiv32_fs724_xor1), .fs_or0(arrdiv32_fs724_or0));
  fs fs_arrdiv32_fs725_out(.a(arrdiv32_mux2to1671_xor0[0]), .b(b[21]), .bin(arrdiv32_fs724_or0[0]), .fs_xor1(arrdiv32_fs725_xor1), .fs_or0(arrdiv32_fs725_or0));
  fs fs_arrdiv32_fs726_out(.a(arrdiv32_mux2to1672_xor0[0]), .b(b[22]), .bin(arrdiv32_fs725_or0[0]), .fs_xor1(arrdiv32_fs726_xor1), .fs_or0(arrdiv32_fs726_or0));
  fs fs_arrdiv32_fs727_out(.a(arrdiv32_mux2to1673_xor0[0]), .b(b[23]), .bin(arrdiv32_fs726_or0[0]), .fs_xor1(arrdiv32_fs727_xor1), .fs_or0(arrdiv32_fs727_or0));
  fs fs_arrdiv32_fs728_out(.a(arrdiv32_mux2to1674_xor0[0]), .b(b[24]), .bin(arrdiv32_fs727_or0[0]), .fs_xor1(arrdiv32_fs728_xor1), .fs_or0(arrdiv32_fs728_or0));
  fs fs_arrdiv32_fs729_out(.a(arrdiv32_mux2to1675_xor0[0]), .b(b[25]), .bin(arrdiv32_fs728_or0[0]), .fs_xor1(arrdiv32_fs729_xor1), .fs_or0(arrdiv32_fs729_or0));
  fs fs_arrdiv32_fs730_out(.a(arrdiv32_mux2to1676_xor0[0]), .b(b[26]), .bin(arrdiv32_fs729_or0[0]), .fs_xor1(arrdiv32_fs730_xor1), .fs_or0(arrdiv32_fs730_or0));
  fs fs_arrdiv32_fs731_out(.a(arrdiv32_mux2to1677_xor0[0]), .b(b[27]), .bin(arrdiv32_fs730_or0[0]), .fs_xor1(arrdiv32_fs731_xor1), .fs_or0(arrdiv32_fs731_or0));
  fs fs_arrdiv32_fs732_out(.a(arrdiv32_mux2to1678_xor0[0]), .b(b[28]), .bin(arrdiv32_fs731_or0[0]), .fs_xor1(arrdiv32_fs732_xor1), .fs_or0(arrdiv32_fs732_or0));
  fs fs_arrdiv32_fs733_out(.a(arrdiv32_mux2to1679_xor0[0]), .b(b[29]), .bin(arrdiv32_fs732_or0[0]), .fs_xor1(arrdiv32_fs733_xor1), .fs_or0(arrdiv32_fs733_or0));
  fs fs_arrdiv32_fs734_out(.a(arrdiv32_mux2to1680_xor0[0]), .b(b[30]), .bin(arrdiv32_fs733_or0[0]), .fs_xor1(arrdiv32_fs734_xor1), .fs_or0(arrdiv32_fs734_or0));
  fs fs_arrdiv32_fs735_out(.a(arrdiv32_mux2to1681_xor0[0]), .b(b[31]), .bin(arrdiv32_fs734_or0[0]), .fs_xor1(arrdiv32_fs735_xor1), .fs_or0(arrdiv32_fs735_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1682_out(.d0(arrdiv32_fs704_xor0[0]), .d1(a[9]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1682_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1683_out(.d0(arrdiv32_fs705_xor1[0]), .d1(arrdiv32_mux2to1651_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1683_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1684_out(.d0(arrdiv32_fs706_xor1[0]), .d1(arrdiv32_mux2to1652_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1684_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1685_out(.d0(arrdiv32_fs707_xor1[0]), .d1(arrdiv32_mux2to1653_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1685_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1686_out(.d0(arrdiv32_fs708_xor1[0]), .d1(arrdiv32_mux2to1654_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1686_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1687_out(.d0(arrdiv32_fs709_xor1[0]), .d1(arrdiv32_mux2to1655_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1687_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1688_out(.d0(arrdiv32_fs710_xor1[0]), .d1(arrdiv32_mux2to1656_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1688_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1689_out(.d0(arrdiv32_fs711_xor1[0]), .d1(arrdiv32_mux2to1657_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1689_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1690_out(.d0(arrdiv32_fs712_xor1[0]), .d1(arrdiv32_mux2to1658_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1690_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1691_out(.d0(arrdiv32_fs713_xor1[0]), .d1(arrdiv32_mux2to1659_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1691_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1692_out(.d0(arrdiv32_fs714_xor1[0]), .d1(arrdiv32_mux2to1660_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1692_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1693_out(.d0(arrdiv32_fs715_xor1[0]), .d1(arrdiv32_mux2to1661_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1693_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1694_out(.d0(arrdiv32_fs716_xor1[0]), .d1(arrdiv32_mux2to1662_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1694_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1695_out(.d0(arrdiv32_fs717_xor1[0]), .d1(arrdiv32_mux2to1663_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1695_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1696_out(.d0(arrdiv32_fs718_xor1[0]), .d1(arrdiv32_mux2to1664_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1696_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1697_out(.d0(arrdiv32_fs719_xor1[0]), .d1(arrdiv32_mux2to1665_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1697_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1698_out(.d0(arrdiv32_fs720_xor1[0]), .d1(arrdiv32_mux2to1666_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1698_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1699_out(.d0(arrdiv32_fs721_xor1[0]), .d1(arrdiv32_mux2to1667_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1699_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1700_out(.d0(arrdiv32_fs722_xor1[0]), .d1(arrdiv32_mux2to1668_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1700_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1701_out(.d0(arrdiv32_fs723_xor1[0]), .d1(arrdiv32_mux2to1669_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1701_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1702_out(.d0(arrdiv32_fs724_xor1[0]), .d1(arrdiv32_mux2to1670_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1702_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1703_out(.d0(arrdiv32_fs725_xor1[0]), .d1(arrdiv32_mux2to1671_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1703_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1704_out(.d0(arrdiv32_fs726_xor1[0]), .d1(arrdiv32_mux2to1672_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1704_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1705_out(.d0(arrdiv32_fs727_xor1[0]), .d1(arrdiv32_mux2to1673_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1705_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1706_out(.d0(arrdiv32_fs728_xor1[0]), .d1(arrdiv32_mux2to1674_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1706_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1707_out(.d0(arrdiv32_fs729_xor1[0]), .d1(arrdiv32_mux2to1675_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1707_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1708_out(.d0(arrdiv32_fs730_xor1[0]), .d1(arrdiv32_mux2to1676_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1708_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1709_out(.d0(arrdiv32_fs731_xor1[0]), .d1(arrdiv32_mux2to1677_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1709_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1710_out(.d0(arrdiv32_fs732_xor1[0]), .d1(arrdiv32_mux2to1678_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1710_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1711_out(.d0(arrdiv32_fs733_xor1[0]), .d1(arrdiv32_mux2to1679_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1711_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1712_out(.d0(arrdiv32_fs734_xor1[0]), .d1(arrdiv32_mux2to1680_xor0[0]), .sel(arrdiv32_fs735_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1712_xor0));
  not_gate not_gate_arrdiv32_not22(.a(arrdiv32_fs735_or0[0]), .out(arrdiv32_not22));
  fs fs_arrdiv32_fs736_out(.a(a[8]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs736_xor0), .fs_or0(arrdiv32_fs736_and0));
  fs fs_arrdiv32_fs737_out(.a(arrdiv32_mux2to1682_xor0[0]), .b(b[1]), .bin(arrdiv32_fs736_and0[0]), .fs_xor1(arrdiv32_fs737_xor1), .fs_or0(arrdiv32_fs737_or0));
  fs fs_arrdiv32_fs738_out(.a(arrdiv32_mux2to1683_xor0[0]), .b(b[2]), .bin(arrdiv32_fs737_or0[0]), .fs_xor1(arrdiv32_fs738_xor1), .fs_or0(arrdiv32_fs738_or0));
  fs fs_arrdiv32_fs739_out(.a(arrdiv32_mux2to1684_xor0[0]), .b(b[3]), .bin(arrdiv32_fs738_or0[0]), .fs_xor1(arrdiv32_fs739_xor1), .fs_or0(arrdiv32_fs739_or0));
  fs fs_arrdiv32_fs740_out(.a(arrdiv32_mux2to1685_xor0[0]), .b(b[4]), .bin(arrdiv32_fs739_or0[0]), .fs_xor1(arrdiv32_fs740_xor1), .fs_or0(arrdiv32_fs740_or0));
  fs fs_arrdiv32_fs741_out(.a(arrdiv32_mux2to1686_xor0[0]), .b(b[5]), .bin(arrdiv32_fs740_or0[0]), .fs_xor1(arrdiv32_fs741_xor1), .fs_or0(arrdiv32_fs741_or0));
  fs fs_arrdiv32_fs742_out(.a(arrdiv32_mux2to1687_xor0[0]), .b(b[6]), .bin(arrdiv32_fs741_or0[0]), .fs_xor1(arrdiv32_fs742_xor1), .fs_or0(arrdiv32_fs742_or0));
  fs fs_arrdiv32_fs743_out(.a(arrdiv32_mux2to1688_xor0[0]), .b(b[7]), .bin(arrdiv32_fs742_or0[0]), .fs_xor1(arrdiv32_fs743_xor1), .fs_or0(arrdiv32_fs743_or0));
  fs fs_arrdiv32_fs744_out(.a(arrdiv32_mux2to1689_xor0[0]), .b(b[8]), .bin(arrdiv32_fs743_or0[0]), .fs_xor1(arrdiv32_fs744_xor1), .fs_or0(arrdiv32_fs744_or0));
  fs fs_arrdiv32_fs745_out(.a(arrdiv32_mux2to1690_xor0[0]), .b(b[9]), .bin(arrdiv32_fs744_or0[0]), .fs_xor1(arrdiv32_fs745_xor1), .fs_or0(arrdiv32_fs745_or0));
  fs fs_arrdiv32_fs746_out(.a(arrdiv32_mux2to1691_xor0[0]), .b(b[10]), .bin(arrdiv32_fs745_or0[0]), .fs_xor1(arrdiv32_fs746_xor1), .fs_or0(arrdiv32_fs746_or0));
  fs fs_arrdiv32_fs747_out(.a(arrdiv32_mux2to1692_xor0[0]), .b(b[11]), .bin(arrdiv32_fs746_or0[0]), .fs_xor1(arrdiv32_fs747_xor1), .fs_or0(arrdiv32_fs747_or0));
  fs fs_arrdiv32_fs748_out(.a(arrdiv32_mux2to1693_xor0[0]), .b(b[12]), .bin(arrdiv32_fs747_or0[0]), .fs_xor1(arrdiv32_fs748_xor1), .fs_or0(arrdiv32_fs748_or0));
  fs fs_arrdiv32_fs749_out(.a(arrdiv32_mux2to1694_xor0[0]), .b(b[13]), .bin(arrdiv32_fs748_or0[0]), .fs_xor1(arrdiv32_fs749_xor1), .fs_or0(arrdiv32_fs749_or0));
  fs fs_arrdiv32_fs750_out(.a(arrdiv32_mux2to1695_xor0[0]), .b(b[14]), .bin(arrdiv32_fs749_or0[0]), .fs_xor1(arrdiv32_fs750_xor1), .fs_or0(arrdiv32_fs750_or0));
  fs fs_arrdiv32_fs751_out(.a(arrdiv32_mux2to1696_xor0[0]), .b(b[15]), .bin(arrdiv32_fs750_or0[0]), .fs_xor1(arrdiv32_fs751_xor1), .fs_or0(arrdiv32_fs751_or0));
  fs fs_arrdiv32_fs752_out(.a(arrdiv32_mux2to1697_xor0[0]), .b(b[16]), .bin(arrdiv32_fs751_or0[0]), .fs_xor1(arrdiv32_fs752_xor1), .fs_or0(arrdiv32_fs752_or0));
  fs fs_arrdiv32_fs753_out(.a(arrdiv32_mux2to1698_xor0[0]), .b(b[17]), .bin(arrdiv32_fs752_or0[0]), .fs_xor1(arrdiv32_fs753_xor1), .fs_or0(arrdiv32_fs753_or0));
  fs fs_arrdiv32_fs754_out(.a(arrdiv32_mux2to1699_xor0[0]), .b(b[18]), .bin(arrdiv32_fs753_or0[0]), .fs_xor1(arrdiv32_fs754_xor1), .fs_or0(arrdiv32_fs754_or0));
  fs fs_arrdiv32_fs755_out(.a(arrdiv32_mux2to1700_xor0[0]), .b(b[19]), .bin(arrdiv32_fs754_or0[0]), .fs_xor1(arrdiv32_fs755_xor1), .fs_or0(arrdiv32_fs755_or0));
  fs fs_arrdiv32_fs756_out(.a(arrdiv32_mux2to1701_xor0[0]), .b(b[20]), .bin(arrdiv32_fs755_or0[0]), .fs_xor1(arrdiv32_fs756_xor1), .fs_or0(arrdiv32_fs756_or0));
  fs fs_arrdiv32_fs757_out(.a(arrdiv32_mux2to1702_xor0[0]), .b(b[21]), .bin(arrdiv32_fs756_or0[0]), .fs_xor1(arrdiv32_fs757_xor1), .fs_or0(arrdiv32_fs757_or0));
  fs fs_arrdiv32_fs758_out(.a(arrdiv32_mux2to1703_xor0[0]), .b(b[22]), .bin(arrdiv32_fs757_or0[0]), .fs_xor1(arrdiv32_fs758_xor1), .fs_or0(arrdiv32_fs758_or0));
  fs fs_arrdiv32_fs759_out(.a(arrdiv32_mux2to1704_xor0[0]), .b(b[23]), .bin(arrdiv32_fs758_or0[0]), .fs_xor1(arrdiv32_fs759_xor1), .fs_or0(arrdiv32_fs759_or0));
  fs fs_arrdiv32_fs760_out(.a(arrdiv32_mux2to1705_xor0[0]), .b(b[24]), .bin(arrdiv32_fs759_or0[0]), .fs_xor1(arrdiv32_fs760_xor1), .fs_or0(arrdiv32_fs760_or0));
  fs fs_arrdiv32_fs761_out(.a(arrdiv32_mux2to1706_xor0[0]), .b(b[25]), .bin(arrdiv32_fs760_or0[0]), .fs_xor1(arrdiv32_fs761_xor1), .fs_or0(arrdiv32_fs761_or0));
  fs fs_arrdiv32_fs762_out(.a(arrdiv32_mux2to1707_xor0[0]), .b(b[26]), .bin(arrdiv32_fs761_or0[0]), .fs_xor1(arrdiv32_fs762_xor1), .fs_or0(arrdiv32_fs762_or0));
  fs fs_arrdiv32_fs763_out(.a(arrdiv32_mux2to1708_xor0[0]), .b(b[27]), .bin(arrdiv32_fs762_or0[0]), .fs_xor1(arrdiv32_fs763_xor1), .fs_or0(arrdiv32_fs763_or0));
  fs fs_arrdiv32_fs764_out(.a(arrdiv32_mux2to1709_xor0[0]), .b(b[28]), .bin(arrdiv32_fs763_or0[0]), .fs_xor1(arrdiv32_fs764_xor1), .fs_or0(arrdiv32_fs764_or0));
  fs fs_arrdiv32_fs765_out(.a(arrdiv32_mux2to1710_xor0[0]), .b(b[29]), .bin(arrdiv32_fs764_or0[0]), .fs_xor1(arrdiv32_fs765_xor1), .fs_or0(arrdiv32_fs765_or0));
  fs fs_arrdiv32_fs766_out(.a(arrdiv32_mux2to1711_xor0[0]), .b(b[30]), .bin(arrdiv32_fs765_or0[0]), .fs_xor1(arrdiv32_fs766_xor1), .fs_or0(arrdiv32_fs766_or0));
  fs fs_arrdiv32_fs767_out(.a(arrdiv32_mux2to1712_xor0[0]), .b(b[31]), .bin(arrdiv32_fs766_or0[0]), .fs_xor1(arrdiv32_fs767_xor1), .fs_or0(arrdiv32_fs767_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1713_out(.d0(arrdiv32_fs736_xor0[0]), .d1(a[8]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1713_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1714_out(.d0(arrdiv32_fs737_xor1[0]), .d1(arrdiv32_mux2to1682_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1714_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1715_out(.d0(arrdiv32_fs738_xor1[0]), .d1(arrdiv32_mux2to1683_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1715_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1716_out(.d0(arrdiv32_fs739_xor1[0]), .d1(arrdiv32_mux2to1684_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1716_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1717_out(.d0(arrdiv32_fs740_xor1[0]), .d1(arrdiv32_mux2to1685_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1717_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1718_out(.d0(arrdiv32_fs741_xor1[0]), .d1(arrdiv32_mux2to1686_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1718_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1719_out(.d0(arrdiv32_fs742_xor1[0]), .d1(arrdiv32_mux2to1687_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1719_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1720_out(.d0(arrdiv32_fs743_xor1[0]), .d1(arrdiv32_mux2to1688_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1720_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1721_out(.d0(arrdiv32_fs744_xor1[0]), .d1(arrdiv32_mux2to1689_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1721_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1722_out(.d0(arrdiv32_fs745_xor1[0]), .d1(arrdiv32_mux2to1690_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1722_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1723_out(.d0(arrdiv32_fs746_xor1[0]), .d1(arrdiv32_mux2to1691_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1723_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1724_out(.d0(arrdiv32_fs747_xor1[0]), .d1(arrdiv32_mux2to1692_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1724_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1725_out(.d0(arrdiv32_fs748_xor1[0]), .d1(arrdiv32_mux2to1693_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1725_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1726_out(.d0(arrdiv32_fs749_xor1[0]), .d1(arrdiv32_mux2to1694_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1726_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1727_out(.d0(arrdiv32_fs750_xor1[0]), .d1(arrdiv32_mux2to1695_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1727_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1728_out(.d0(arrdiv32_fs751_xor1[0]), .d1(arrdiv32_mux2to1696_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1728_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1729_out(.d0(arrdiv32_fs752_xor1[0]), .d1(arrdiv32_mux2to1697_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1729_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1730_out(.d0(arrdiv32_fs753_xor1[0]), .d1(arrdiv32_mux2to1698_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1730_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1731_out(.d0(arrdiv32_fs754_xor1[0]), .d1(arrdiv32_mux2to1699_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1731_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1732_out(.d0(arrdiv32_fs755_xor1[0]), .d1(arrdiv32_mux2to1700_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1732_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1733_out(.d0(arrdiv32_fs756_xor1[0]), .d1(arrdiv32_mux2to1701_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1733_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1734_out(.d0(arrdiv32_fs757_xor1[0]), .d1(arrdiv32_mux2to1702_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1734_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1735_out(.d0(arrdiv32_fs758_xor1[0]), .d1(arrdiv32_mux2to1703_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1735_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1736_out(.d0(arrdiv32_fs759_xor1[0]), .d1(arrdiv32_mux2to1704_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1736_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1737_out(.d0(arrdiv32_fs760_xor1[0]), .d1(arrdiv32_mux2to1705_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1737_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1738_out(.d0(arrdiv32_fs761_xor1[0]), .d1(arrdiv32_mux2to1706_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1738_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1739_out(.d0(arrdiv32_fs762_xor1[0]), .d1(arrdiv32_mux2to1707_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1739_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1740_out(.d0(arrdiv32_fs763_xor1[0]), .d1(arrdiv32_mux2to1708_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1740_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1741_out(.d0(arrdiv32_fs764_xor1[0]), .d1(arrdiv32_mux2to1709_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1741_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1742_out(.d0(arrdiv32_fs765_xor1[0]), .d1(arrdiv32_mux2to1710_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1742_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1743_out(.d0(arrdiv32_fs766_xor1[0]), .d1(arrdiv32_mux2to1711_xor0[0]), .sel(arrdiv32_fs767_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1743_xor0));
  not_gate not_gate_arrdiv32_not23(.a(arrdiv32_fs767_or0[0]), .out(arrdiv32_not23));
  fs fs_arrdiv32_fs768_out(.a(a[7]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs768_xor0), .fs_or0(arrdiv32_fs768_and0));
  fs fs_arrdiv32_fs769_out(.a(arrdiv32_mux2to1713_xor0[0]), .b(b[1]), .bin(arrdiv32_fs768_and0[0]), .fs_xor1(arrdiv32_fs769_xor1), .fs_or0(arrdiv32_fs769_or0));
  fs fs_arrdiv32_fs770_out(.a(arrdiv32_mux2to1714_xor0[0]), .b(b[2]), .bin(arrdiv32_fs769_or0[0]), .fs_xor1(arrdiv32_fs770_xor1), .fs_or0(arrdiv32_fs770_or0));
  fs fs_arrdiv32_fs771_out(.a(arrdiv32_mux2to1715_xor0[0]), .b(b[3]), .bin(arrdiv32_fs770_or0[0]), .fs_xor1(arrdiv32_fs771_xor1), .fs_or0(arrdiv32_fs771_or0));
  fs fs_arrdiv32_fs772_out(.a(arrdiv32_mux2to1716_xor0[0]), .b(b[4]), .bin(arrdiv32_fs771_or0[0]), .fs_xor1(arrdiv32_fs772_xor1), .fs_or0(arrdiv32_fs772_or0));
  fs fs_arrdiv32_fs773_out(.a(arrdiv32_mux2to1717_xor0[0]), .b(b[5]), .bin(arrdiv32_fs772_or0[0]), .fs_xor1(arrdiv32_fs773_xor1), .fs_or0(arrdiv32_fs773_or0));
  fs fs_arrdiv32_fs774_out(.a(arrdiv32_mux2to1718_xor0[0]), .b(b[6]), .bin(arrdiv32_fs773_or0[0]), .fs_xor1(arrdiv32_fs774_xor1), .fs_or0(arrdiv32_fs774_or0));
  fs fs_arrdiv32_fs775_out(.a(arrdiv32_mux2to1719_xor0[0]), .b(b[7]), .bin(arrdiv32_fs774_or0[0]), .fs_xor1(arrdiv32_fs775_xor1), .fs_or0(arrdiv32_fs775_or0));
  fs fs_arrdiv32_fs776_out(.a(arrdiv32_mux2to1720_xor0[0]), .b(b[8]), .bin(arrdiv32_fs775_or0[0]), .fs_xor1(arrdiv32_fs776_xor1), .fs_or0(arrdiv32_fs776_or0));
  fs fs_arrdiv32_fs777_out(.a(arrdiv32_mux2to1721_xor0[0]), .b(b[9]), .bin(arrdiv32_fs776_or0[0]), .fs_xor1(arrdiv32_fs777_xor1), .fs_or0(arrdiv32_fs777_or0));
  fs fs_arrdiv32_fs778_out(.a(arrdiv32_mux2to1722_xor0[0]), .b(b[10]), .bin(arrdiv32_fs777_or0[0]), .fs_xor1(arrdiv32_fs778_xor1), .fs_or0(arrdiv32_fs778_or0));
  fs fs_arrdiv32_fs779_out(.a(arrdiv32_mux2to1723_xor0[0]), .b(b[11]), .bin(arrdiv32_fs778_or0[0]), .fs_xor1(arrdiv32_fs779_xor1), .fs_or0(arrdiv32_fs779_or0));
  fs fs_arrdiv32_fs780_out(.a(arrdiv32_mux2to1724_xor0[0]), .b(b[12]), .bin(arrdiv32_fs779_or0[0]), .fs_xor1(arrdiv32_fs780_xor1), .fs_or0(arrdiv32_fs780_or0));
  fs fs_arrdiv32_fs781_out(.a(arrdiv32_mux2to1725_xor0[0]), .b(b[13]), .bin(arrdiv32_fs780_or0[0]), .fs_xor1(arrdiv32_fs781_xor1), .fs_or0(arrdiv32_fs781_or0));
  fs fs_arrdiv32_fs782_out(.a(arrdiv32_mux2to1726_xor0[0]), .b(b[14]), .bin(arrdiv32_fs781_or0[0]), .fs_xor1(arrdiv32_fs782_xor1), .fs_or0(arrdiv32_fs782_or0));
  fs fs_arrdiv32_fs783_out(.a(arrdiv32_mux2to1727_xor0[0]), .b(b[15]), .bin(arrdiv32_fs782_or0[0]), .fs_xor1(arrdiv32_fs783_xor1), .fs_or0(arrdiv32_fs783_or0));
  fs fs_arrdiv32_fs784_out(.a(arrdiv32_mux2to1728_xor0[0]), .b(b[16]), .bin(arrdiv32_fs783_or0[0]), .fs_xor1(arrdiv32_fs784_xor1), .fs_or0(arrdiv32_fs784_or0));
  fs fs_arrdiv32_fs785_out(.a(arrdiv32_mux2to1729_xor0[0]), .b(b[17]), .bin(arrdiv32_fs784_or0[0]), .fs_xor1(arrdiv32_fs785_xor1), .fs_or0(arrdiv32_fs785_or0));
  fs fs_arrdiv32_fs786_out(.a(arrdiv32_mux2to1730_xor0[0]), .b(b[18]), .bin(arrdiv32_fs785_or0[0]), .fs_xor1(arrdiv32_fs786_xor1), .fs_or0(arrdiv32_fs786_or0));
  fs fs_arrdiv32_fs787_out(.a(arrdiv32_mux2to1731_xor0[0]), .b(b[19]), .bin(arrdiv32_fs786_or0[0]), .fs_xor1(arrdiv32_fs787_xor1), .fs_or0(arrdiv32_fs787_or0));
  fs fs_arrdiv32_fs788_out(.a(arrdiv32_mux2to1732_xor0[0]), .b(b[20]), .bin(arrdiv32_fs787_or0[0]), .fs_xor1(arrdiv32_fs788_xor1), .fs_or0(arrdiv32_fs788_or0));
  fs fs_arrdiv32_fs789_out(.a(arrdiv32_mux2to1733_xor0[0]), .b(b[21]), .bin(arrdiv32_fs788_or0[0]), .fs_xor1(arrdiv32_fs789_xor1), .fs_or0(arrdiv32_fs789_or0));
  fs fs_arrdiv32_fs790_out(.a(arrdiv32_mux2to1734_xor0[0]), .b(b[22]), .bin(arrdiv32_fs789_or0[0]), .fs_xor1(arrdiv32_fs790_xor1), .fs_or0(arrdiv32_fs790_or0));
  fs fs_arrdiv32_fs791_out(.a(arrdiv32_mux2to1735_xor0[0]), .b(b[23]), .bin(arrdiv32_fs790_or0[0]), .fs_xor1(arrdiv32_fs791_xor1), .fs_or0(arrdiv32_fs791_or0));
  fs fs_arrdiv32_fs792_out(.a(arrdiv32_mux2to1736_xor0[0]), .b(b[24]), .bin(arrdiv32_fs791_or0[0]), .fs_xor1(arrdiv32_fs792_xor1), .fs_or0(arrdiv32_fs792_or0));
  fs fs_arrdiv32_fs793_out(.a(arrdiv32_mux2to1737_xor0[0]), .b(b[25]), .bin(arrdiv32_fs792_or0[0]), .fs_xor1(arrdiv32_fs793_xor1), .fs_or0(arrdiv32_fs793_or0));
  fs fs_arrdiv32_fs794_out(.a(arrdiv32_mux2to1738_xor0[0]), .b(b[26]), .bin(arrdiv32_fs793_or0[0]), .fs_xor1(arrdiv32_fs794_xor1), .fs_or0(arrdiv32_fs794_or0));
  fs fs_arrdiv32_fs795_out(.a(arrdiv32_mux2to1739_xor0[0]), .b(b[27]), .bin(arrdiv32_fs794_or0[0]), .fs_xor1(arrdiv32_fs795_xor1), .fs_or0(arrdiv32_fs795_or0));
  fs fs_arrdiv32_fs796_out(.a(arrdiv32_mux2to1740_xor0[0]), .b(b[28]), .bin(arrdiv32_fs795_or0[0]), .fs_xor1(arrdiv32_fs796_xor1), .fs_or0(arrdiv32_fs796_or0));
  fs fs_arrdiv32_fs797_out(.a(arrdiv32_mux2to1741_xor0[0]), .b(b[29]), .bin(arrdiv32_fs796_or0[0]), .fs_xor1(arrdiv32_fs797_xor1), .fs_or0(arrdiv32_fs797_or0));
  fs fs_arrdiv32_fs798_out(.a(arrdiv32_mux2to1742_xor0[0]), .b(b[30]), .bin(arrdiv32_fs797_or0[0]), .fs_xor1(arrdiv32_fs798_xor1), .fs_or0(arrdiv32_fs798_or0));
  fs fs_arrdiv32_fs799_out(.a(arrdiv32_mux2to1743_xor0[0]), .b(b[31]), .bin(arrdiv32_fs798_or0[0]), .fs_xor1(arrdiv32_fs799_xor1), .fs_or0(arrdiv32_fs799_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1744_out(.d0(arrdiv32_fs768_xor0[0]), .d1(a[7]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1744_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1745_out(.d0(arrdiv32_fs769_xor1[0]), .d1(arrdiv32_mux2to1713_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1745_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1746_out(.d0(arrdiv32_fs770_xor1[0]), .d1(arrdiv32_mux2to1714_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1746_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1747_out(.d0(arrdiv32_fs771_xor1[0]), .d1(arrdiv32_mux2to1715_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1747_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1748_out(.d0(arrdiv32_fs772_xor1[0]), .d1(arrdiv32_mux2to1716_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1748_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1749_out(.d0(arrdiv32_fs773_xor1[0]), .d1(arrdiv32_mux2to1717_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1749_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1750_out(.d0(arrdiv32_fs774_xor1[0]), .d1(arrdiv32_mux2to1718_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1750_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1751_out(.d0(arrdiv32_fs775_xor1[0]), .d1(arrdiv32_mux2to1719_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1751_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1752_out(.d0(arrdiv32_fs776_xor1[0]), .d1(arrdiv32_mux2to1720_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1752_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1753_out(.d0(arrdiv32_fs777_xor1[0]), .d1(arrdiv32_mux2to1721_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1753_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1754_out(.d0(arrdiv32_fs778_xor1[0]), .d1(arrdiv32_mux2to1722_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1754_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1755_out(.d0(arrdiv32_fs779_xor1[0]), .d1(arrdiv32_mux2to1723_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1755_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1756_out(.d0(arrdiv32_fs780_xor1[0]), .d1(arrdiv32_mux2to1724_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1756_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1757_out(.d0(arrdiv32_fs781_xor1[0]), .d1(arrdiv32_mux2to1725_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1757_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1758_out(.d0(arrdiv32_fs782_xor1[0]), .d1(arrdiv32_mux2to1726_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1758_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1759_out(.d0(arrdiv32_fs783_xor1[0]), .d1(arrdiv32_mux2to1727_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1759_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1760_out(.d0(arrdiv32_fs784_xor1[0]), .d1(arrdiv32_mux2to1728_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1760_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1761_out(.d0(arrdiv32_fs785_xor1[0]), .d1(arrdiv32_mux2to1729_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1761_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1762_out(.d0(arrdiv32_fs786_xor1[0]), .d1(arrdiv32_mux2to1730_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1762_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1763_out(.d0(arrdiv32_fs787_xor1[0]), .d1(arrdiv32_mux2to1731_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1763_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1764_out(.d0(arrdiv32_fs788_xor1[0]), .d1(arrdiv32_mux2to1732_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1764_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1765_out(.d0(arrdiv32_fs789_xor1[0]), .d1(arrdiv32_mux2to1733_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1765_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1766_out(.d0(arrdiv32_fs790_xor1[0]), .d1(arrdiv32_mux2to1734_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1766_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1767_out(.d0(arrdiv32_fs791_xor1[0]), .d1(arrdiv32_mux2to1735_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1767_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1768_out(.d0(arrdiv32_fs792_xor1[0]), .d1(arrdiv32_mux2to1736_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1768_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1769_out(.d0(arrdiv32_fs793_xor1[0]), .d1(arrdiv32_mux2to1737_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1769_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1770_out(.d0(arrdiv32_fs794_xor1[0]), .d1(arrdiv32_mux2to1738_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1770_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1771_out(.d0(arrdiv32_fs795_xor1[0]), .d1(arrdiv32_mux2to1739_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1771_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1772_out(.d0(arrdiv32_fs796_xor1[0]), .d1(arrdiv32_mux2to1740_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1772_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1773_out(.d0(arrdiv32_fs797_xor1[0]), .d1(arrdiv32_mux2to1741_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1773_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1774_out(.d0(arrdiv32_fs798_xor1[0]), .d1(arrdiv32_mux2to1742_xor0[0]), .sel(arrdiv32_fs799_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1774_xor0));
  not_gate not_gate_arrdiv32_not24(.a(arrdiv32_fs799_or0[0]), .out(arrdiv32_not24));
  fs fs_arrdiv32_fs800_out(.a(a[6]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs800_xor0), .fs_or0(arrdiv32_fs800_and0));
  fs fs_arrdiv32_fs801_out(.a(arrdiv32_mux2to1744_xor0[0]), .b(b[1]), .bin(arrdiv32_fs800_and0[0]), .fs_xor1(arrdiv32_fs801_xor1), .fs_or0(arrdiv32_fs801_or0));
  fs fs_arrdiv32_fs802_out(.a(arrdiv32_mux2to1745_xor0[0]), .b(b[2]), .bin(arrdiv32_fs801_or0[0]), .fs_xor1(arrdiv32_fs802_xor1), .fs_or0(arrdiv32_fs802_or0));
  fs fs_arrdiv32_fs803_out(.a(arrdiv32_mux2to1746_xor0[0]), .b(b[3]), .bin(arrdiv32_fs802_or0[0]), .fs_xor1(arrdiv32_fs803_xor1), .fs_or0(arrdiv32_fs803_or0));
  fs fs_arrdiv32_fs804_out(.a(arrdiv32_mux2to1747_xor0[0]), .b(b[4]), .bin(arrdiv32_fs803_or0[0]), .fs_xor1(arrdiv32_fs804_xor1), .fs_or0(arrdiv32_fs804_or0));
  fs fs_arrdiv32_fs805_out(.a(arrdiv32_mux2to1748_xor0[0]), .b(b[5]), .bin(arrdiv32_fs804_or0[0]), .fs_xor1(arrdiv32_fs805_xor1), .fs_or0(arrdiv32_fs805_or0));
  fs fs_arrdiv32_fs806_out(.a(arrdiv32_mux2to1749_xor0[0]), .b(b[6]), .bin(arrdiv32_fs805_or0[0]), .fs_xor1(arrdiv32_fs806_xor1), .fs_or0(arrdiv32_fs806_or0));
  fs fs_arrdiv32_fs807_out(.a(arrdiv32_mux2to1750_xor0[0]), .b(b[7]), .bin(arrdiv32_fs806_or0[0]), .fs_xor1(arrdiv32_fs807_xor1), .fs_or0(arrdiv32_fs807_or0));
  fs fs_arrdiv32_fs808_out(.a(arrdiv32_mux2to1751_xor0[0]), .b(b[8]), .bin(arrdiv32_fs807_or0[0]), .fs_xor1(arrdiv32_fs808_xor1), .fs_or0(arrdiv32_fs808_or0));
  fs fs_arrdiv32_fs809_out(.a(arrdiv32_mux2to1752_xor0[0]), .b(b[9]), .bin(arrdiv32_fs808_or0[0]), .fs_xor1(arrdiv32_fs809_xor1), .fs_or0(arrdiv32_fs809_or0));
  fs fs_arrdiv32_fs810_out(.a(arrdiv32_mux2to1753_xor0[0]), .b(b[10]), .bin(arrdiv32_fs809_or0[0]), .fs_xor1(arrdiv32_fs810_xor1), .fs_or0(arrdiv32_fs810_or0));
  fs fs_arrdiv32_fs811_out(.a(arrdiv32_mux2to1754_xor0[0]), .b(b[11]), .bin(arrdiv32_fs810_or0[0]), .fs_xor1(arrdiv32_fs811_xor1), .fs_or0(arrdiv32_fs811_or0));
  fs fs_arrdiv32_fs812_out(.a(arrdiv32_mux2to1755_xor0[0]), .b(b[12]), .bin(arrdiv32_fs811_or0[0]), .fs_xor1(arrdiv32_fs812_xor1), .fs_or0(arrdiv32_fs812_or0));
  fs fs_arrdiv32_fs813_out(.a(arrdiv32_mux2to1756_xor0[0]), .b(b[13]), .bin(arrdiv32_fs812_or0[0]), .fs_xor1(arrdiv32_fs813_xor1), .fs_or0(arrdiv32_fs813_or0));
  fs fs_arrdiv32_fs814_out(.a(arrdiv32_mux2to1757_xor0[0]), .b(b[14]), .bin(arrdiv32_fs813_or0[0]), .fs_xor1(arrdiv32_fs814_xor1), .fs_or0(arrdiv32_fs814_or0));
  fs fs_arrdiv32_fs815_out(.a(arrdiv32_mux2to1758_xor0[0]), .b(b[15]), .bin(arrdiv32_fs814_or0[0]), .fs_xor1(arrdiv32_fs815_xor1), .fs_or0(arrdiv32_fs815_or0));
  fs fs_arrdiv32_fs816_out(.a(arrdiv32_mux2to1759_xor0[0]), .b(b[16]), .bin(arrdiv32_fs815_or0[0]), .fs_xor1(arrdiv32_fs816_xor1), .fs_or0(arrdiv32_fs816_or0));
  fs fs_arrdiv32_fs817_out(.a(arrdiv32_mux2to1760_xor0[0]), .b(b[17]), .bin(arrdiv32_fs816_or0[0]), .fs_xor1(arrdiv32_fs817_xor1), .fs_or0(arrdiv32_fs817_or0));
  fs fs_arrdiv32_fs818_out(.a(arrdiv32_mux2to1761_xor0[0]), .b(b[18]), .bin(arrdiv32_fs817_or0[0]), .fs_xor1(arrdiv32_fs818_xor1), .fs_or0(arrdiv32_fs818_or0));
  fs fs_arrdiv32_fs819_out(.a(arrdiv32_mux2to1762_xor0[0]), .b(b[19]), .bin(arrdiv32_fs818_or0[0]), .fs_xor1(arrdiv32_fs819_xor1), .fs_or0(arrdiv32_fs819_or0));
  fs fs_arrdiv32_fs820_out(.a(arrdiv32_mux2to1763_xor0[0]), .b(b[20]), .bin(arrdiv32_fs819_or0[0]), .fs_xor1(arrdiv32_fs820_xor1), .fs_or0(arrdiv32_fs820_or0));
  fs fs_arrdiv32_fs821_out(.a(arrdiv32_mux2to1764_xor0[0]), .b(b[21]), .bin(arrdiv32_fs820_or0[0]), .fs_xor1(arrdiv32_fs821_xor1), .fs_or0(arrdiv32_fs821_or0));
  fs fs_arrdiv32_fs822_out(.a(arrdiv32_mux2to1765_xor0[0]), .b(b[22]), .bin(arrdiv32_fs821_or0[0]), .fs_xor1(arrdiv32_fs822_xor1), .fs_or0(arrdiv32_fs822_or0));
  fs fs_arrdiv32_fs823_out(.a(arrdiv32_mux2to1766_xor0[0]), .b(b[23]), .bin(arrdiv32_fs822_or0[0]), .fs_xor1(arrdiv32_fs823_xor1), .fs_or0(arrdiv32_fs823_or0));
  fs fs_arrdiv32_fs824_out(.a(arrdiv32_mux2to1767_xor0[0]), .b(b[24]), .bin(arrdiv32_fs823_or0[0]), .fs_xor1(arrdiv32_fs824_xor1), .fs_or0(arrdiv32_fs824_or0));
  fs fs_arrdiv32_fs825_out(.a(arrdiv32_mux2to1768_xor0[0]), .b(b[25]), .bin(arrdiv32_fs824_or0[0]), .fs_xor1(arrdiv32_fs825_xor1), .fs_or0(arrdiv32_fs825_or0));
  fs fs_arrdiv32_fs826_out(.a(arrdiv32_mux2to1769_xor0[0]), .b(b[26]), .bin(arrdiv32_fs825_or0[0]), .fs_xor1(arrdiv32_fs826_xor1), .fs_or0(arrdiv32_fs826_or0));
  fs fs_arrdiv32_fs827_out(.a(arrdiv32_mux2to1770_xor0[0]), .b(b[27]), .bin(arrdiv32_fs826_or0[0]), .fs_xor1(arrdiv32_fs827_xor1), .fs_or0(arrdiv32_fs827_or0));
  fs fs_arrdiv32_fs828_out(.a(arrdiv32_mux2to1771_xor0[0]), .b(b[28]), .bin(arrdiv32_fs827_or0[0]), .fs_xor1(arrdiv32_fs828_xor1), .fs_or0(arrdiv32_fs828_or0));
  fs fs_arrdiv32_fs829_out(.a(arrdiv32_mux2to1772_xor0[0]), .b(b[29]), .bin(arrdiv32_fs828_or0[0]), .fs_xor1(arrdiv32_fs829_xor1), .fs_or0(arrdiv32_fs829_or0));
  fs fs_arrdiv32_fs830_out(.a(arrdiv32_mux2to1773_xor0[0]), .b(b[30]), .bin(arrdiv32_fs829_or0[0]), .fs_xor1(arrdiv32_fs830_xor1), .fs_or0(arrdiv32_fs830_or0));
  fs fs_arrdiv32_fs831_out(.a(arrdiv32_mux2to1774_xor0[0]), .b(b[31]), .bin(arrdiv32_fs830_or0[0]), .fs_xor1(arrdiv32_fs831_xor1), .fs_or0(arrdiv32_fs831_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1775_out(.d0(arrdiv32_fs800_xor0[0]), .d1(a[6]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1775_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1776_out(.d0(arrdiv32_fs801_xor1[0]), .d1(arrdiv32_mux2to1744_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1776_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1777_out(.d0(arrdiv32_fs802_xor1[0]), .d1(arrdiv32_mux2to1745_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1777_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1778_out(.d0(arrdiv32_fs803_xor1[0]), .d1(arrdiv32_mux2to1746_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1778_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1779_out(.d0(arrdiv32_fs804_xor1[0]), .d1(arrdiv32_mux2to1747_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1779_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1780_out(.d0(arrdiv32_fs805_xor1[0]), .d1(arrdiv32_mux2to1748_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1780_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1781_out(.d0(arrdiv32_fs806_xor1[0]), .d1(arrdiv32_mux2to1749_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1781_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1782_out(.d0(arrdiv32_fs807_xor1[0]), .d1(arrdiv32_mux2to1750_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1782_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1783_out(.d0(arrdiv32_fs808_xor1[0]), .d1(arrdiv32_mux2to1751_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1783_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1784_out(.d0(arrdiv32_fs809_xor1[0]), .d1(arrdiv32_mux2to1752_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1784_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1785_out(.d0(arrdiv32_fs810_xor1[0]), .d1(arrdiv32_mux2to1753_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1785_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1786_out(.d0(arrdiv32_fs811_xor1[0]), .d1(arrdiv32_mux2to1754_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1786_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1787_out(.d0(arrdiv32_fs812_xor1[0]), .d1(arrdiv32_mux2to1755_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1787_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1788_out(.d0(arrdiv32_fs813_xor1[0]), .d1(arrdiv32_mux2to1756_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1788_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1789_out(.d0(arrdiv32_fs814_xor1[0]), .d1(arrdiv32_mux2to1757_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1789_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1790_out(.d0(arrdiv32_fs815_xor1[0]), .d1(arrdiv32_mux2to1758_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1790_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1791_out(.d0(arrdiv32_fs816_xor1[0]), .d1(arrdiv32_mux2to1759_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1791_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1792_out(.d0(arrdiv32_fs817_xor1[0]), .d1(arrdiv32_mux2to1760_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1792_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1793_out(.d0(arrdiv32_fs818_xor1[0]), .d1(arrdiv32_mux2to1761_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1793_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1794_out(.d0(arrdiv32_fs819_xor1[0]), .d1(arrdiv32_mux2to1762_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1794_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1795_out(.d0(arrdiv32_fs820_xor1[0]), .d1(arrdiv32_mux2to1763_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1795_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1796_out(.d0(arrdiv32_fs821_xor1[0]), .d1(arrdiv32_mux2to1764_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1796_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1797_out(.d0(arrdiv32_fs822_xor1[0]), .d1(arrdiv32_mux2to1765_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1797_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1798_out(.d0(arrdiv32_fs823_xor1[0]), .d1(arrdiv32_mux2to1766_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1798_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1799_out(.d0(arrdiv32_fs824_xor1[0]), .d1(arrdiv32_mux2to1767_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1799_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1800_out(.d0(arrdiv32_fs825_xor1[0]), .d1(arrdiv32_mux2to1768_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1800_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1801_out(.d0(arrdiv32_fs826_xor1[0]), .d1(arrdiv32_mux2to1769_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1801_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1802_out(.d0(arrdiv32_fs827_xor1[0]), .d1(arrdiv32_mux2to1770_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1802_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1803_out(.d0(arrdiv32_fs828_xor1[0]), .d1(arrdiv32_mux2to1771_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1803_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1804_out(.d0(arrdiv32_fs829_xor1[0]), .d1(arrdiv32_mux2to1772_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1804_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1805_out(.d0(arrdiv32_fs830_xor1[0]), .d1(arrdiv32_mux2to1773_xor0[0]), .sel(arrdiv32_fs831_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1805_xor0));
  not_gate not_gate_arrdiv32_not25(.a(arrdiv32_fs831_or0[0]), .out(arrdiv32_not25));
  fs fs_arrdiv32_fs832_out(.a(a[5]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs832_xor0), .fs_or0(arrdiv32_fs832_and0));
  fs fs_arrdiv32_fs833_out(.a(arrdiv32_mux2to1775_xor0[0]), .b(b[1]), .bin(arrdiv32_fs832_and0[0]), .fs_xor1(arrdiv32_fs833_xor1), .fs_or0(arrdiv32_fs833_or0));
  fs fs_arrdiv32_fs834_out(.a(arrdiv32_mux2to1776_xor0[0]), .b(b[2]), .bin(arrdiv32_fs833_or0[0]), .fs_xor1(arrdiv32_fs834_xor1), .fs_or0(arrdiv32_fs834_or0));
  fs fs_arrdiv32_fs835_out(.a(arrdiv32_mux2to1777_xor0[0]), .b(b[3]), .bin(arrdiv32_fs834_or0[0]), .fs_xor1(arrdiv32_fs835_xor1), .fs_or0(arrdiv32_fs835_or0));
  fs fs_arrdiv32_fs836_out(.a(arrdiv32_mux2to1778_xor0[0]), .b(b[4]), .bin(arrdiv32_fs835_or0[0]), .fs_xor1(arrdiv32_fs836_xor1), .fs_or0(arrdiv32_fs836_or0));
  fs fs_arrdiv32_fs837_out(.a(arrdiv32_mux2to1779_xor0[0]), .b(b[5]), .bin(arrdiv32_fs836_or0[0]), .fs_xor1(arrdiv32_fs837_xor1), .fs_or0(arrdiv32_fs837_or0));
  fs fs_arrdiv32_fs838_out(.a(arrdiv32_mux2to1780_xor0[0]), .b(b[6]), .bin(arrdiv32_fs837_or0[0]), .fs_xor1(arrdiv32_fs838_xor1), .fs_or0(arrdiv32_fs838_or0));
  fs fs_arrdiv32_fs839_out(.a(arrdiv32_mux2to1781_xor0[0]), .b(b[7]), .bin(arrdiv32_fs838_or0[0]), .fs_xor1(arrdiv32_fs839_xor1), .fs_or0(arrdiv32_fs839_or0));
  fs fs_arrdiv32_fs840_out(.a(arrdiv32_mux2to1782_xor0[0]), .b(b[8]), .bin(arrdiv32_fs839_or0[0]), .fs_xor1(arrdiv32_fs840_xor1), .fs_or0(arrdiv32_fs840_or0));
  fs fs_arrdiv32_fs841_out(.a(arrdiv32_mux2to1783_xor0[0]), .b(b[9]), .bin(arrdiv32_fs840_or0[0]), .fs_xor1(arrdiv32_fs841_xor1), .fs_or0(arrdiv32_fs841_or0));
  fs fs_arrdiv32_fs842_out(.a(arrdiv32_mux2to1784_xor0[0]), .b(b[10]), .bin(arrdiv32_fs841_or0[0]), .fs_xor1(arrdiv32_fs842_xor1), .fs_or0(arrdiv32_fs842_or0));
  fs fs_arrdiv32_fs843_out(.a(arrdiv32_mux2to1785_xor0[0]), .b(b[11]), .bin(arrdiv32_fs842_or0[0]), .fs_xor1(arrdiv32_fs843_xor1), .fs_or0(arrdiv32_fs843_or0));
  fs fs_arrdiv32_fs844_out(.a(arrdiv32_mux2to1786_xor0[0]), .b(b[12]), .bin(arrdiv32_fs843_or0[0]), .fs_xor1(arrdiv32_fs844_xor1), .fs_or0(arrdiv32_fs844_or0));
  fs fs_arrdiv32_fs845_out(.a(arrdiv32_mux2to1787_xor0[0]), .b(b[13]), .bin(arrdiv32_fs844_or0[0]), .fs_xor1(arrdiv32_fs845_xor1), .fs_or0(arrdiv32_fs845_or0));
  fs fs_arrdiv32_fs846_out(.a(arrdiv32_mux2to1788_xor0[0]), .b(b[14]), .bin(arrdiv32_fs845_or0[0]), .fs_xor1(arrdiv32_fs846_xor1), .fs_or0(arrdiv32_fs846_or0));
  fs fs_arrdiv32_fs847_out(.a(arrdiv32_mux2to1789_xor0[0]), .b(b[15]), .bin(arrdiv32_fs846_or0[0]), .fs_xor1(arrdiv32_fs847_xor1), .fs_or0(arrdiv32_fs847_or0));
  fs fs_arrdiv32_fs848_out(.a(arrdiv32_mux2to1790_xor0[0]), .b(b[16]), .bin(arrdiv32_fs847_or0[0]), .fs_xor1(arrdiv32_fs848_xor1), .fs_or0(arrdiv32_fs848_or0));
  fs fs_arrdiv32_fs849_out(.a(arrdiv32_mux2to1791_xor0[0]), .b(b[17]), .bin(arrdiv32_fs848_or0[0]), .fs_xor1(arrdiv32_fs849_xor1), .fs_or0(arrdiv32_fs849_or0));
  fs fs_arrdiv32_fs850_out(.a(arrdiv32_mux2to1792_xor0[0]), .b(b[18]), .bin(arrdiv32_fs849_or0[0]), .fs_xor1(arrdiv32_fs850_xor1), .fs_or0(arrdiv32_fs850_or0));
  fs fs_arrdiv32_fs851_out(.a(arrdiv32_mux2to1793_xor0[0]), .b(b[19]), .bin(arrdiv32_fs850_or0[0]), .fs_xor1(arrdiv32_fs851_xor1), .fs_or0(arrdiv32_fs851_or0));
  fs fs_arrdiv32_fs852_out(.a(arrdiv32_mux2to1794_xor0[0]), .b(b[20]), .bin(arrdiv32_fs851_or0[0]), .fs_xor1(arrdiv32_fs852_xor1), .fs_or0(arrdiv32_fs852_or0));
  fs fs_arrdiv32_fs853_out(.a(arrdiv32_mux2to1795_xor0[0]), .b(b[21]), .bin(arrdiv32_fs852_or0[0]), .fs_xor1(arrdiv32_fs853_xor1), .fs_or0(arrdiv32_fs853_or0));
  fs fs_arrdiv32_fs854_out(.a(arrdiv32_mux2to1796_xor0[0]), .b(b[22]), .bin(arrdiv32_fs853_or0[0]), .fs_xor1(arrdiv32_fs854_xor1), .fs_or0(arrdiv32_fs854_or0));
  fs fs_arrdiv32_fs855_out(.a(arrdiv32_mux2to1797_xor0[0]), .b(b[23]), .bin(arrdiv32_fs854_or0[0]), .fs_xor1(arrdiv32_fs855_xor1), .fs_or0(arrdiv32_fs855_or0));
  fs fs_arrdiv32_fs856_out(.a(arrdiv32_mux2to1798_xor0[0]), .b(b[24]), .bin(arrdiv32_fs855_or0[0]), .fs_xor1(arrdiv32_fs856_xor1), .fs_or0(arrdiv32_fs856_or0));
  fs fs_arrdiv32_fs857_out(.a(arrdiv32_mux2to1799_xor0[0]), .b(b[25]), .bin(arrdiv32_fs856_or0[0]), .fs_xor1(arrdiv32_fs857_xor1), .fs_or0(arrdiv32_fs857_or0));
  fs fs_arrdiv32_fs858_out(.a(arrdiv32_mux2to1800_xor0[0]), .b(b[26]), .bin(arrdiv32_fs857_or0[0]), .fs_xor1(arrdiv32_fs858_xor1), .fs_or0(arrdiv32_fs858_or0));
  fs fs_arrdiv32_fs859_out(.a(arrdiv32_mux2to1801_xor0[0]), .b(b[27]), .bin(arrdiv32_fs858_or0[0]), .fs_xor1(arrdiv32_fs859_xor1), .fs_or0(arrdiv32_fs859_or0));
  fs fs_arrdiv32_fs860_out(.a(arrdiv32_mux2to1802_xor0[0]), .b(b[28]), .bin(arrdiv32_fs859_or0[0]), .fs_xor1(arrdiv32_fs860_xor1), .fs_or0(arrdiv32_fs860_or0));
  fs fs_arrdiv32_fs861_out(.a(arrdiv32_mux2to1803_xor0[0]), .b(b[29]), .bin(arrdiv32_fs860_or0[0]), .fs_xor1(arrdiv32_fs861_xor1), .fs_or0(arrdiv32_fs861_or0));
  fs fs_arrdiv32_fs862_out(.a(arrdiv32_mux2to1804_xor0[0]), .b(b[30]), .bin(arrdiv32_fs861_or0[0]), .fs_xor1(arrdiv32_fs862_xor1), .fs_or0(arrdiv32_fs862_or0));
  fs fs_arrdiv32_fs863_out(.a(arrdiv32_mux2to1805_xor0[0]), .b(b[31]), .bin(arrdiv32_fs862_or0[0]), .fs_xor1(arrdiv32_fs863_xor1), .fs_or0(arrdiv32_fs863_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1806_out(.d0(arrdiv32_fs832_xor0[0]), .d1(a[5]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1806_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1807_out(.d0(arrdiv32_fs833_xor1[0]), .d1(arrdiv32_mux2to1775_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1807_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1808_out(.d0(arrdiv32_fs834_xor1[0]), .d1(arrdiv32_mux2to1776_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1808_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1809_out(.d0(arrdiv32_fs835_xor1[0]), .d1(arrdiv32_mux2to1777_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1809_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1810_out(.d0(arrdiv32_fs836_xor1[0]), .d1(arrdiv32_mux2to1778_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1810_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1811_out(.d0(arrdiv32_fs837_xor1[0]), .d1(arrdiv32_mux2to1779_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1811_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1812_out(.d0(arrdiv32_fs838_xor1[0]), .d1(arrdiv32_mux2to1780_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1812_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1813_out(.d0(arrdiv32_fs839_xor1[0]), .d1(arrdiv32_mux2to1781_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1813_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1814_out(.d0(arrdiv32_fs840_xor1[0]), .d1(arrdiv32_mux2to1782_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1814_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1815_out(.d0(arrdiv32_fs841_xor1[0]), .d1(arrdiv32_mux2to1783_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1815_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1816_out(.d0(arrdiv32_fs842_xor1[0]), .d1(arrdiv32_mux2to1784_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1816_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1817_out(.d0(arrdiv32_fs843_xor1[0]), .d1(arrdiv32_mux2to1785_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1817_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1818_out(.d0(arrdiv32_fs844_xor1[0]), .d1(arrdiv32_mux2to1786_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1818_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1819_out(.d0(arrdiv32_fs845_xor1[0]), .d1(arrdiv32_mux2to1787_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1819_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1820_out(.d0(arrdiv32_fs846_xor1[0]), .d1(arrdiv32_mux2to1788_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1820_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1821_out(.d0(arrdiv32_fs847_xor1[0]), .d1(arrdiv32_mux2to1789_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1821_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1822_out(.d0(arrdiv32_fs848_xor1[0]), .d1(arrdiv32_mux2to1790_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1822_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1823_out(.d0(arrdiv32_fs849_xor1[0]), .d1(arrdiv32_mux2to1791_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1823_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1824_out(.d0(arrdiv32_fs850_xor1[0]), .d1(arrdiv32_mux2to1792_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1824_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1825_out(.d0(arrdiv32_fs851_xor1[0]), .d1(arrdiv32_mux2to1793_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1825_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1826_out(.d0(arrdiv32_fs852_xor1[0]), .d1(arrdiv32_mux2to1794_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1826_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1827_out(.d0(arrdiv32_fs853_xor1[0]), .d1(arrdiv32_mux2to1795_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1827_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1828_out(.d0(arrdiv32_fs854_xor1[0]), .d1(arrdiv32_mux2to1796_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1828_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1829_out(.d0(arrdiv32_fs855_xor1[0]), .d1(arrdiv32_mux2to1797_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1829_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1830_out(.d0(arrdiv32_fs856_xor1[0]), .d1(arrdiv32_mux2to1798_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1830_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1831_out(.d0(arrdiv32_fs857_xor1[0]), .d1(arrdiv32_mux2to1799_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1831_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1832_out(.d0(arrdiv32_fs858_xor1[0]), .d1(arrdiv32_mux2to1800_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1832_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1833_out(.d0(arrdiv32_fs859_xor1[0]), .d1(arrdiv32_mux2to1801_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1833_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1834_out(.d0(arrdiv32_fs860_xor1[0]), .d1(arrdiv32_mux2to1802_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1834_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1835_out(.d0(arrdiv32_fs861_xor1[0]), .d1(arrdiv32_mux2to1803_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1835_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1836_out(.d0(arrdiv32_fs862_xor1[0]), .d1(arrdiv32_mux2to1804_xor0[0]), .sel(arrdiv32_fs863_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1836_xor0));
  not_gate not_gate_arrdiv32_not26(.a(arrdiv32_fs863_or0[0]), .out(arrdiv32_not26));
  fs fs_arrdiv32_fs864_out(.a(a[4]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs864_xor0), .fs_or0(arrdiv32_fs864_and0));
  fs fs_arrdiv32_fs865_out(.a(arrdiv32_mux2to1806_xor0[0]), .b(b[1]), .bin(arrdiv32_fs864_and0[0]), .fs_xor1(arrdiv32_fs865_xor1), .fs_or0(arrdiv32_fs865_or0));
  fs fs_arrdiv32_fs866_out(.a(arrdiv32_mux2to1807_xor0[0]), .b(b[2]), .bin(arrdiv32_fs865_or0[0]), .fs_xor1(arrdiv32_fs866_xor1), .fs_or0(arrdiv32_fs866_or0));
  fs fs_arrdiv32_fs867_out(.a(arrdiv32_mux2to1808_xor0[0]), .b(b[3]), .bin(arrdiv32_fs866_or0[0]), .fs_xor1(arrdiv32_fs867_xor1), .fs_or0(arrdiv32_fs867_or0));
  fs fs_arrdiv32_fs868_out(.a(arrdiv32_mux2to1809_xor0[0]), .b(b[4]), .bin(arrdiv32_fs867_or0[0]), .fs_xor1(arrdiv32_fs868_xor1), .fs_or0(arrdiv32_fs868_or0));
  fs fs_arrdiv32_fs869_out(.a(arrdiv32_mux2to1810_xor0[0]), .b(b[5]), .bin(arrdiv32_fs868_or0[0]), .fs_xor1(arrdiv32_fs869_xor1), .fs_or0(arrdiv32_fs869_or0));
  fs fs_arrdiv32_fs870_out(.a(arrdiv32_mux2to1811_xor0[0]), .b(b[6]), .bin(arrdiv32_fs869_or0[0]), .fs_xor1(arrdiv32_fs870_xor1), .fs_or0(arrdiv32_fs870_or0));
  fs fs_arrdiv32_fs871_out(.a(arrdiv32_mux2to1812_xor0[0]), .b(b[7]), .bin(arrdiv32_fs870_or0[0]), .fs_xor1(arrdiv32_fs871_xor1), .fs_or0(arrdiv32_fs871_or0));
  fs fs_arrdiv32_fs872_out(.a(arrdiv32_mux2to1813_xor0[0]), .b(b[8]), .bin(arrdiv32_fs871_or0[0]), .fs_xor1(arrdiv32_fs872_xor1), .fs_or0(arrdiv32_fs872_or0));
  fs fs_arrdiv32_fs873_out(.a(arrdiv32_mux2to1814_xor0[0]), .b(b[9]), .bin(arrdiv32_fs872_or0[0]), .fs_xor1(arrdiv32_fs873_xor1), .fs_or0(arrdiv32_fs873_or0));
  fs fs_arrdiv32_fs874_out(.a(arrdiv32_mux2to1815_xor0[0]), .b(b[10]), .bin(arrdiv32_fs873_or0[0]), .fs_xor1(arrdiv32_fs874_xor1), .fs_or0(arrdiv32_fs874_or0));
  fs fs_arrdiv32_fs875_out(.a(arrdiv32_mux2to1816_xor0[0]), .b(b[11]), .bin(arrdiv32_fs874_or0[0]), .fs_xor1(arrdiv32_fs875_xor1), .fs_or0(arrdiv32_fs875_or0));
  fs fs_arrdiv32_fs876_out(.a(arrdiv32_mux2to1817_xor0[0]), .b(b[12]), .bin(arrdiv32_fs875_or0[0]), .fs_xor1(arrdiv32_fs876_xor1), .fs_or0(arrdiv32_fs876_or0));
  fs fs_arrdiv32_fs877_out(.a(arrdiv32_mux2to1818_xor0[0]), .b(b[13]), .bin(arrdiv32_fs876_or0[0]), .fs_xor1(arrdiv32_fs877_xor1), .fs_or0(arrdiv32_fs877_or0));
  fs fs_arrdiv32_fs878_out(.a(arrdiv32_mux2to1819_xor0[0]), .b(b[14]), .bin(arrdiv32_fs877_or0[0]), .fs_xor1(arrdiv32_fs878_xor1), .fs_or0(arrdiv32_fs878_or0));
  fs fs_arrdiv32_fs879_out(.a(arrdiv32_mux2to1820_xor0[0]), .b(b[15]), .bin(arrdiv32_fs878_or0[0]), .fs_xor1(arrdiv32_fs879_xor1), .fs_or0(arrdiv32_fs879_or0));
  fs fs_arrdiv32_fs880_out(.a(arrdiv32_mux2to1821_xor0[0]), .b(b[16]), .bin(arrdiv32_fs879_or0[0]), .fs_xor1(arrdiv32_fs880_xor1), .fs_or0(arrdiv32_fs880_or0));
  fs fs_arrdiv32_fs881_out(.a(arrdiv32_mux2to1822_xor0[0]), .b(b[17]), .bin(arrdiv32_fs880_or0[0]), .fs_xor1(arrdiv32_fs881_xor1), .fs_or0(arrdiv32_fs881_or0));
  fs fs_arrdiv32_fs882_out(.a(arrdiv32_mux2to1823_xor0[0]), .b(b[18]), .bin(arrdiv32_fs881_or0[0]), .fs_xor1(arrdiv32_fs882_xor1), .fs_or0(arrdiv32_fs882_or0));
  fs fs_arrdiv32_fs883_out(.a(arrdiv32_mux2to1824_xor0[0]), .b(b[19]), .bin(arrdiv32_fs882_or0[0]), .fs_xor1(arrdiv32_fs883_xor1), .fs_or0(arrdiv32_fs883_or0));
  fs fs_arrdiv32_fs884_out(.a(arrdiv32_mux2to1825_xor0[0]), .b(b[20]), .bin(arrdiv32_fs883_or0[0]), .fs_xor1(arrdiv32_fs884_xor1), .fs_or0(arrdiv32_fs884_or0));
  fs fs_arrdiv32_fs885_out(.a(arrdiv32_mux2to1826_xor0[0]), .b(b[21]), .bin(arrdiv32_fs884_or0[0]), .fs_xor1(arrdiv32_fs885_xor1), .fs_or0(arrdiv32_fs885_or0));
  fs fs_arrdiv32_fs886_out(.a(arrdiv32_mux2to1827_xor0[0]), .b(b[22]), .bin(arrdiv32_fs885_or0[0]), .fs_xor1(arrdiv32_fs886_xor1), .fs_or0(arrdiv32_fs886_or0));
  fs fs_arrdiv32_fs887_out(.a(arrdiv32_mux2to1828_xor0[0]), .b(b[23]), .bin(arrdiv32_fs886_or0[0]), .fs_xor1(arrdiv32_fs887_xor1), .fs_or0(arrdiv32_fs887_or0));
  fs fs_arrdiv32_fs888_out(.a(arrdiv32_mux2to1829_xor0[0]), .b(b[24]), .bin(arrdiv32_fs887_or0[0]), .fs_xor1(arrdiv32_fs888_xor1), .fs_or0(arrdiv32_fs888_or0));
  fs fs_arrdiv32_fs889_out(.a(arrdiv32_mux2to1830_xor0[0]), .b(b[25]), .bin(arrdiv32_fs888_or0[0]), .fs_xor1(arrdiv32_fs889_xor1), .fs_or0(arrdiv32_fs889_or0));
  fs fs_arrdiv32_fs890_out(.a(arrdiv32_mux2to1831_xor0[0]), .b(b[26]), .bin(arrdiv32_fs889_or0[0]), .fs_xor1(arrdiv32_fs890_xor1), .fs_or0(arrdiv32_fs890_or0));
  fs fs_arrdiv32_fs891_out(.a(arrdiv32_mux2to1832_xor0[0]), .b(b[27]), .bin(arrdiv32_fs890_or0[0]), .fs_xor1(arrdiv32_fs891_xor1), .fs_or0(arrdiv32_fs891_or0));
  fs fs_arrdiv32_fs892_out(.a(arrdiv32_mux2to1833_xor0[0]), .b(b[28]), .bin(arrdiv32_fs891_or0[0]), .fs_xor1(arrdiv32_fs892_xor1), .fs_or0(arrdiv32_fs892_or0));
  fs fs_arrdiv32_fs893_out(.a(arrdiv32_mux2to1834_xor0[0]), .b(b[29]), .bin(arrdiv32_fs892_or0[0]), .fs_xor1(arrdiv32_fs893_xor1), .fs_or0(arrdiv32_fs893_or0));
  fs fs_arrdiv32_fs894_out(.a(arrdiv32_mux2to1835_xor0[0]), .b(b[30]), .bin(arrdiv32_fs893_or0[0]), .fs_xor1(arrdiv32_fs894_xor1), .fs_or0(arrdiv32_fs894_or0));
  fs fs_arrdiv32_fs895_out(.a(arrdiv32_mux2to1836_xor0[0]), .b(b[31]), .bin(arrdiv32_fs894_or0[0]), .fs_xor1(arrdiv32_fs895_xor1), .fs_or0(arrdiv32_fs895_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1837_out(.d0(arrdiv32_fs864_xor0[0]), .d1(a[4]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1837_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1838_out(.d0(arrdiv32_fs865_xor1[0]), .d1(arrdiv32_mux2to1806_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1838_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1839_out(.d0(arrdiv32_fs866_xor1[0]), .d1(arrdiv32_mux2to1807_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1839_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1840_out(.d0(arrdiv32_fs867_xor1[0]), .d1(arrdiv32_mux2to1808_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1840_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1841_out(.d0(arrdiv32_fs868_xor1[0]), .d1(arrdiv32_mux2to1809_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1841_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1842_out(.d0(arrdiv32_fs869_xor1[0]), .d1(arrdiv32_mux2to1810_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1842_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1843_out(.d0(arrdiv32_fs870_xor1[0]), .d1(arrdiv32_mux2to1811_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1843_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1844_out(.d0(arrdiv32_fs871_xor1[0]), .d1(arrdiv32_mux2to1812_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1844_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1845_out(.d0(arrdiv32_fs872_xor1[0]), .d1(arrdiv32_mux2to1813_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1845_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1846_out(.d0(arrdiv32_fs873_xor1[0]), .d1(arrdiv32_mux2to1814_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1846_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1847_out(.d0(arrdiv32_fs874_xor1[0]), .d1(arrdiv32_mux2to1815_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1847_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1848_out(.d0(arrdiv32_fs875_xor1[0]), .d1(arrdiv32_mux2to1816_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1848_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1849_out(.d0(arrdiv32_fs876_xor1[0]), .d1(arrdiv32_mux2to1817_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1849_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1850_out(.d0(arrdiv32_fs877_xor1[0]), .d1(arrdiv32_mux2to1818_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1850_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1851_out(.d0(arrdiv32_fs878_xor1[0]), .d1(arrdiv32_mux2to1819_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1851_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1852_out(.d0(arrdiv32_fs879_xor1[0]), .d1(arrdiv32_mux2to1820_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1852_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1853_out(.d0(arrdiv32_fs880_xor1[0]), .d1(arrdiv32_mux2to1821_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1853_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1854_out(.d0(arrdiv32_fs881_xor1[0]), .d1(arrdiv32_mux2to1822_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1854_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1855_out(.d0(arrdiv32_fs882_xor1[0]), .d1(arrdiv32_mux2to1823_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1855_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1856_out(.d0(arrdiv32_fs883_xor1[0]), .d1(arrdiv32_mux2to1824_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1856_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1857_out(.d0(arrdiv32_fs884_xor1[0]), .d1(arrdiv32_mux2to1825_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1857_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1858_out(.d0(arrdiv32_fs885_xor1[0]), .d1(arrdiv32_mux2to1826_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1858_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1859_out(.d0(arrdiv32_fs886_xor1[0]), .d1(arrdiv32_mux2to1827_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1859_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1860_out(.d0(arrdiv32_fs887_xor1[0]), .d1(arrdiv32_mux2to1828_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1860_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1861_out(.d0(arrdiv32_fs888_xor1[0]), .d1(arrdiv32_mux2to1829_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1861_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1862_out(.d0(arrdiv32_fs889_xor1[0]), .d1(arrdiv32_mux2to1830_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1862_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1863_out(.d0(arrdiv32_fs890_xor1[0]), .d1(arrdiv32_mux2to1831_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1863_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1864_out(.d0(arrdiv32_fs891_xor1[0]), .d1(arrdiv32_mux2to1832_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1864_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1865_out(.d0(arrdiv32_fs892_xor1[0]), .d1(arrdiv32_mux2to1833_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1865_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1866_out(.d0(arrdiv32_fs893_xor1[0]), .d1(arrdiv32_mux2to1834_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1866_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1867_out(.d0(arrdiv32_fs894_xor1[0]), .d1(arrdiv32_mux2to1835_xor0[0]), .sel(arrdiv32_fs895_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1867_xor0));
  not_gate not_gate_arrdiv32_not27(.a(arrdiv32_fs895_or0[0]), .out(arrdiv32_not27));
  fs fs_arrdiv32_fs896_out(.a(a[3]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs896_xor0), .fs_or0(arrdiv32_fs896_and0));
  fs fs_arrdiv32_fs897_out(.a(arrdiv32_mux2to1837_xor0[0]), .b(b[1]), .bin(arrdiv32_fs896_and0[0]), .fs_xor1(arrdiv32_fs897_xor1), .fs_or0(arrdiv32_fs897_or0));
  fs fs_arrdiv32_fs898_out(.a(arrdiv32_mux2to1838_xor0[0]), .b(b[2]), .bin(arrdiv32_fs897_or0[0]), .fs_xor1(arrdiv32_fs898_xor1), .fs_or0(arrdiv32_fs898_or0));
  fs fs_arrdiv32_fs899_out(.a(arrdiv32_mux2to1839_xor0[0]), .b(b[3]), .bin(arrdiv32_fs898_or0[0]), .fs_xor1(arrdiv32_fs899_xor1), .fs_or0(arrdiv32_fs899_or0));
  fs fs_arrdiv32_fs900_out(.a(arrdiv32_mux2to1840_xor0[0]), .b(b[4]), .bin(arrdiv32_fs899_or0[0]), .fs_xor1(arrdiv32_fs900_xor1), .fs_or0(arrdiv32_fs900_or0));
  fs fs_arrdiv32_fs901_out(.a(arrdiv32_mux2to1841_xor0[0]), .b(b[5]), .bin(arrdiv32_fs900_or0[0]), .fs_xor1(arrdiv32_fs901_xor1), .fs_or0(arrdiv32_fs901_or0));
  fs fs_arrdiv32_fs902_out(.a(arrdiv32_mux2to1842_xor0[0]), .b(b[6]), .bin(arrdiv32_fs901_or0[0]), .fs_xor1(arrdiv32_fs902_xor1), .fs_or0(arrdiv32_fs902_or0));
  fs fs_arrdiv32_fs903_out(.a(arrdiv32_mux2to1843_xor0[0]), .b(b[7]), .bin(arrdiv32_fs902_or0[0]), .fs_xor1(arrdiv32_fs903_xor1), .fs_or0(arrdiv32_fs903_or0));
  fs fs_arrdiv32_fs904_out(.a(arrdiv32_mux2to1844_xor0[0]), .b(b[8]), .bin(arrdiv32_fs903_or0[0]), .fs_xor1(arrdiv32_fs904_xor1), .fs_or0(arrdiv32_fs904_or0));
  fs fs_arrdiv32_fs905_out(.a(arrdiv32_mux2to1845_xor0[0]), .b(b[9]), .bin(arrdiv32_fs904_or0[0]), .fs_xor1(arrdiv32_fs905_xor1), .fs_or0(arrdiv32_fs905_or0));
  fs fs_arrdiv32_fs906_out(.a(arrdiv32_mux2to1846_xor0[0]), .b(b[10]), .bin(arrdiv32_fs905_or0[0]), .fs_xor1(arrdiv32_fs906_xor1), .fs_or0(arrdiv32_fs906_or0));
  fs fs_arrdiv32_fs907_out(.a(arrdiv32_mux2to1847_xor0[0]), .b(b[11]), .bin(arrdiv32_fs906_or0[0]), .fs_xor1(arrdiv32_fs907_xor1), .fs_or0(arrdiv32_fs907_or0));
  fs fs_arrdiv32_fs908_out(.a(arrdiv32_mux2to1848_xor0[0]), .b(b[12]), .bin(arrdiv32_fs907_or0[0]), .fs_xor1(arrdiv32_fs908_xor1), .fs_or0(arrdiv32_fs908_or0));
  fs fs_arrdiv32_fs909_out(.a(arrdiv32_mux2to1849_xor0[0]), .b(b[13]), .bin(arrdiv32_fs908_or0[0]), .fs_xor1(arrdiv32_fs909_xor1), .fs_or0(arrdiv32_fs909_or0));
  fs fs_arrdiv32_fs910_out(.a(arrdiv32_mux2to1850_xor0[0]), .b(b[14]), .bin(arrdiv32_fs909_or0[0]), .fs_xor1(arrdiv32_fs910_xor1), .fs_or0(arrdiv32_fs910_or0));
  fs fs_arrdiv32_fs911_out(.a(arrdiv32_mux2to1851_xor0[0]), .b(b[15]), .bin(arrdiv32_fs910_or0[0]), .fs_xor1(arrdiv32_fs911_xor1), .fs_or0(arrdiv32_fs911_or0));
  fs fs_arrdiv32_fs912_out(.a(arrdiv32_mux2to1852_xor0[0]), .b(b[16]), .bin(arrdiv32_fs911_or0[0]), .fs_xor1(arrdiv32_fs912_xor1), .fs_or0(arrdiv32_fs912_or0));
  fs fs_arrdiv32_fs913_out(.a(arrdiv32_mux2to1853_xor0[0]), .b(b[17]), .bin(arrdiv32_fs912_or0[0]), .fs_xor1(arrdiv32_fs913_xor1), .fs_or0(arrdiv32_fs913_or0));
  fs fs_arrdiv32_fs914_out(.a(arrdiv32_mux2to1854_xor0[0]), .b(b[18]), .bin(arrdiv32_fs913_or0[0]), .fs_xor1(arrdiv32_fs914_xor1), .fs_or0(arrdiv32_fs914_or0));
  fs fs_arrdiv32_fs915_out(.a(arrdiv32_mux2to1855_xor0[0]), .b(b[19]), .bin(arrdiv32_fs914_or0[0]), .fs_xor1(arrdiv32_fs915_xor1), .fs_or0(arrdiv32_fs915_or0));
  fs fs_arrdiv32_fs916_out(.a(arrdiv32_mux2to1856_xor0[0]), .b(b[20]), .bin(arrdiv32_fs915_or0[0]), .fs_xor1(arrdiv32_fs916_xor1), .fs_or0(arrdiv32_fs916_or0));
  fs fs_arrdiv32_fs917_out(.a(arrdiv32_mux2to1857_xor0[0]), .b(b[21]), .bin(arrdiv32_fs916_or0[0]), .fs_xor1(arrdiv32_fs917_xor1), .fs_or0(arrdiv32_fs917_or0));
  fs fs_arrdiv32_fs918_out(.a(arrdiv32_mux2to1858_xor0[0]), .b(b[22]), .bin(arrdiv32_fs917_or0[0]), .fs_xor1(arrdiv32_fs918_xor1), .fs_or0(arrdiv32_fs918_or0));
  fs fs_arrdiv32_fs919_out(.a(arrdiv32_mux2to1859_xor0[0]), .b(b[23]), .bin(arrdiv32_fs918_or0[0]), .fs_xor1(arrdiv32_fs919_xor1), .fs_or0(arrdiv32_fs919_or0));
  fs fs_arrdiv32_fs920_out(.a(arrdiv32_mux2to1860_xor0[0]), .b(b[24]), .bin(arrdiv32_fs919_or0[0]), .fs_xor1(arrdiv32_fs920_xor1), .fs_or0(arrdiv32_fs920_or0));
  fs fs_arrdiv32_fs921_out(.a(arrdiv32_mux2to1861_xor0[0]), .b(b[25]), .bin(arrdiv32_fs920_or0[0]), .fs_xor1(arrdiv32_fs921_xor1), .fs_or0(arrdiv32_fs921_or0));
  fs fs_arrdiv32_fs922_out(.a(arrdiv32_mux2to1862_xor0[0]), .b(b[26]), .bin(arrdiv32_fs921_or0[0]), .fs_xor1(arrdiv32_fs922_xor1), .fs_or0(arrdiv32_fs922_or0));
  fs fs_arrdiv32_fs923_out(.a(arrdiv32_mux2to1863_xor0[0]), .b(b[27]), .bin(arrdiv32_fs922_or0[0]), .fs_xor1(arrdiv32_fs923_xor1), .fs_or0(arrdiv32_fs923_or0));
  fs fs_arrdiv32_fs924_out(.a(arrdiv32_mux2to1864_xor0[0]), .b(b[28]), .bin(arrdiv32_fs923_or0[0]), .fs_xor1(arrdiv32_fs924_xor1), .fs_or0(arrdiv32_fs924_or0));
  fs fs_arrdiv32_fs925_out(.a(arrdiv32_mux2to1865_xor0[0]), .b(b[29]), .bin(arrdiv32_fs924_or0[0]), .fs_xor1(arrdiv32_fs925_xor1), .fs_or0(arrdiv32_fs925_or0));
  fs fs_arrdiv32_fs926_out(.a(arrdiv32_mux2to1866_xor0[0]), .b(b[30]), .bin(arrdiv32_fs925_or0[0]), .fs_xor1(arrdiv32_fs926_xor1), .fs_or0(arrdiv32_fs926_or0));
  fs fs_arrdiv32_fs927_out(.a(arrdiv32_mux2to1867_xor0[0]), .b(b[31]), .bin(arrdiv32_fs926_or0[0]), .fs_xor1(arrdiv32_fs927_xor1), .fs_or0(arrdiv32_fs927_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1868_out(.d0(arrdiv32_fs896_xor0[0]), .d1(a[3]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1868_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1869_out(.d0(arrdiv32_fs897_xor1[0]), .d1(arrdiv32_mux2to1837_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1869_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1870_out(.d0(arrdiv32_fs898_xor1[0]), .d1(arrdiv32_mux2to1838_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1870_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1871_out(.d0(arrdiv32_fs899_xor1[0]), .d1(arrdiv32_mux2to1839_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1871_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1872_out(.d0(arrdiv32_fs900_xor1[0]), .d1(arrdiv32_mux2to1840_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1872_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1873_out(.d0(arrdiv32_fs901_xor1[0]), .d1(arrdiv32_mux2to1841_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1873_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1874_out(.d0(arrdiv32_fs902_xor1[0]), .d1(arrdiv32_mux2to1842_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1874_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1875_out(.d0(arrdiv32_fs903_xor1[0]), .d1(arrdiv32_mux2to1843_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1875_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1876_out(.d0(arrdiv32_fs904_xor1[0]), .d1(arrdiv32_mux2to1844_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1876_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1877_out(.d0(arrdiv32_fs905_xor1[0]), .d1(arrdiv32_mux2to1845_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1877_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1878_out(.d0(arrdiv32_fs906_xor1[0]), .d1(arrdiv32_mux2to1846_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1878_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1879_out(.d0(arrdiv32_fs907_xor1[0]), .d1(arrdiv32_mux2to1847_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1879_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1880_out(.d0(arrdiv32_fs908_xor1[0]), .d1(arrdiv32_mux2to1848_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1880_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1881_out(.d0(arrdiv32_fs909_xor1[0]), .d1(arrdiv32_mux2to1849_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1881_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1882_out(.d0(arrdiv32_fs910_xor1[0]), .d1(arrdiv32_mux2to1850_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1882_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1883_out(.d0(arrdiv32_fs911_xor1[0]), .d1(arrdiv32_mux2to1851_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1883_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1884_out(.d0(arrdiv32_fs912_xor1[0]), .d1(arrdiv32_mux2to1852_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1884_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1885_out(.d0(arrdiv32_fs913_xor1[0]), .d1(arrdiv32_mux2to1853_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1885_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1886_out(.d0(arrdiv32_fs914_xor1[0]), .d1(arrdiv32_mux2to1854_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1886_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1887_out(.d0(arrdiv32_fs915_xor1[0]), .d1(arrdiv32_mux2to1855_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1887_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1888_out(.d0(arrdiv32_fs916_xor1[0]), .d1(arrdiv32_mux2to1856_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1888_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1889_out(.d0(arrdiv32_fs917_xor1[0]), .d1(arrdiv32_mux2to1857_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1889_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1890_out(.d0(arrdiv32_fs918_xor1[0]), .d1(arrdiv32_mux2to1858_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1890_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1891_out(.d0(arrdiv32_fs919_xor1[0]), .d1(arrdiv32_mux2to1859_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1891_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1892_out(.d0(arrdiv32_fs920_xor1[0]), .d1(arrdiv32_mux2to1860_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1892_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1893_out(.d0(arrdiv32_fs921_xor1[0]), .d1(arrdiv32_mux2to1861_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1893_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1894_out(.d0(arrdiv32_fs922_xor1[0]), .d1(arrdiv32_mux2to1862_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1894_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1895_out(.d0(arrdiv32_fs923_xor1[0]), .d1(arrdiv32_mux2to1863_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1895_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1896_out(.d0(arrdiv32_fs924_xor1[0]), .d1(arrdiv32_mux2to1864_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1896_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1897_out(.d0(arrdiv32_fs925_xor1[0]), .d1(arrdiv32_mux2to1865_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1897_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1898_out(.d0(arrdiv32_fs926_xor1[0]), .d1(arrdiv32_mux2to1866_xor0[0]), .sel(arrdiv32_fs927_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1898_xor0));
  not_gate not_gate_arrdiv32_not28(.a(arrdiv32_fs927_or0[0]), .out(arrdiv32_not28));
  fs fs_arrdiv32_fs928_out(.a(a[2]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs928_xor0), .fs_or0(arrdiv32_fs928_and0));
  fs fs_arrdiv32_fs929_out(.a(arrdiv32_mux2to1868_xor0[0]), .b(b[1]), .bin(arrdiv32_fs928_and0[0]), .fs_xor1(arrdiv32_fs929_xor1), .fs_or0(arrdiv32_fs929_or0));
  fs fs_arrdiv32_fs930_out(.a(arrdiv32_mux2to1869_xor0[0]), .b(b[2]), .bin(arrdiv32_fs929_or0[0]), .fs_xor1(arrdiv32_fs930_xor1), .fs_or0(arrdiv32_fs930_or0));
  fs fs_arrdiv32_fs931_out(.a(arrdiv32_mux2to1870_xor0[0]), .b(b[3]), .bin(arrdiv32_fs930_or0[0]), .fs_xor1(arrdiv32_fs931_xor1), .fs_or0(arrdiv32_fs931_or0));
  fs fs_arrdiv32_fs932_out(.a(arrdiv32_mux2to1871_xor0[0]), .b(b[4]), .bin(arrdiv32_fs931_or0[0]), .fs_xor1(arrdiv32_fs932_xor1), .fs_or0(arrdiv32_fs932_or0));
  fs fs_arrdiv32_fs933_out(.a(arrdiv32_mux2to1872_xor0[0]), .b(b[5]), .bin(arrdiv32_fs932_or0[0]), .fs_xor1(arrdiv32_fs933_xor1), .fs_or0(arrdiv32_fs933_or0));
  fs fs_arrdiv32_fs934_out(.a(arrdiv32_mux2to1873_xor0[0]), .b(b[6]), .bin(arrdiv32_fs933_or0[0]), .fs_xor1(arrdiv32_fs934_xor1), .fs_or0(arrdiv32_fs934_or0));
  fs fs_arrdiv32_fs935_out(.a(arrdiv32_mux2to1874_xor0[0]), .b(b[7]), .bin(arrdiv32_fs934_or0[0]), .fs_xor1(arrdiv32_fs935_xor1), .fs_or0(arrdiv32_fs935_or0));
  fs fs_arrdiv32_fs936_out(.a(arrdiv32_mux2to1875_xor0[0]), .b(b[8]), .bin(arrdiv32_fs935_or0[0]), .fs_xor1(arrdiv32_fs936_xor1), .fs_or0(arrdiv32_fs936_or0));
  fs fs_arrdiv32_fs937_out(.a(arrdiv32_mux2to1876_xor0[0]), .b(b[9]), .bin(arrdiv32_fs936_or0[0]), .fs_xor1(arrdiv32_fs937_xor1), .fs_or0(arrdiv32_fs937_or0));
  fs fs_arrdiv32_fs938_out(.a(arrdiv32_mux2to1877_xor0[0]), .b(b[10]), .bin(arrdiv32_fs937_or0[0]), .fs_xor1(arrdiv32_fs938_xor1), .fs_or0(arrdiv32_fs938_or0));
  fs fs_arrdiv32_fs939_out(.a(arrdiv32_mux2to1878_xor0[0]), .b(b[11]), .bin(arrdiv32_fs938_or0[0]), .fs_xor1(arrdiv32_fs939_xor1), .fs_or0(arrdiv32_fs939_or0));
  fs fs_arrdiv32_fs940_out(.a(arrdiv32_mux2to1879_xor0[0]), .b(b[12]), .bin(arrdiv32_fs939_or0[0]), .fs_xor1(arrdiv32_fs940_xor1), .fs_or0(arrdiv32_fs940_or0));
  fs fs_arrdiv32_fs941_out(.a(arrdiv32_mux2to1880_xor0[0]), .b(b[13]), .bin(arrdiv32_fs940_or0[0]), .fs_xor1(arrdiv32_fs941_xor1), .fs_or0(arrdiv32_fs941_or0));
  fs fs_arrdiv32_fs942_out(.a(arrdiv32_mux2to1881_xor0[0]), .b(b[14]), .bin(arrdiv32_fs941_or0[0]), .fs_xor1(arrdiv32_fs942_xor1), .fs_or0(arrdiv32_fs942_or0));
  fs fs_arrdiv32_fs943_out(.a(arrdiv32_mux2to1882_xor0[0]), .b(b[15]), .bin(arrdiv32_fs942_or0[0]), .fs_xor1(arrdiv32_fs943_xor1), .fs_or0(arrdiv32_fs943_or0));
  fs fs_arrdiv32_fs944_out(.a(arrdiv32_mux2to1883_xor0[0]), .b(b[16]), .bin(arrdiv32_fs943_or0[0]), .fs_xor1(arrdiv32_fs944_xor1), .fs_or0(arrdiv32_fs944_or0));
  fs fs_arrdiv32_fs945_out(.a(arrdiv32_mux2to1884_xor0[0]), .b(b[17]), .bin(arrdiv32_fs944_or0[0]), .fs_xor1(arrdiv32_fs945_xor1), .fs_or0(arrdiv32_fs945_or0));
  fs fs_arrdiv32_fs946_out(.a(arrdiv32_mux2to1885_xor0[0]), .b(b[18]), .bin(arrdiv32_fs945_or0[0]), .fs_xor1(arrdiv32_fs946_xor1), .fs_or0(arrdiv32_fs946_or0));
  fs fs_arrdiv32_fs947_out(.a(arrdiv32_mux2to1886_xor0[0]), .b(b[19]), .bin(arrdiv32_fs946_or0[0]), .fs_xor1(arrdiv32_fs947_xor1), .fs_or0(arrdiv32_fs947_or0));
  fs fs_arrdiv32_fs948_out(.a(arrdiv32_mux2to1887_xor0[0]), .b(b[20]), .bin(arrdiv32_fs947_or0[0]), .fs_xor1(arrdiv32_fs948_xor1), .fs_or0(arrdiv32_fs948_or0));
  fs fs_arrdiv32_fs949_out(.a(arrdiv32_mux2to1888_xor0[0]), .b(b[21]), .bin(arrdiv32_fs948_or0[0]), .fs_xor1(arrdiv32_fs949_xor1), .fs_or0(arrdiv32_fs949_or0));
  fs fs_arrdiv32_fs950_out(.a(arrdiv32_mux2to1889_xor0[0]), .b(b[22]), .bin(arrdiv32_fs949_or0[0]), .fs_xor1(arrdiv32_fs950_xor1), .fs_or0(arrdiv32_fs950_or0));
  fs fs_arrdiv32_fs951_out(.a(arrdiv32_mux2to1890_xor0[0]), .b(b[23]), .bin(arrdiv32_fs950_or0[0]), .fs_xor1(arrdiv32_fs951_xor1), .fs_or0(arrdiv32_fs951_or0));
  fs fs_arrdiv32_fs952_out(.a(arrdiv32_mux2to1891_xor0[0]), .b(b[24]), .bin(arrdiv32_fs951_or0[0]), .fs_xor1(arrdiv32_fs952_xor1), .fs_or0(arrdiv32_fs952_or0));
  fs fs_arrdiv32_fs953_out(.a(arrdiv32_mux2to1892_xor0[0]), .b(b[25]), .bin(arrdiv32_fs952_or0[0]), .fs_xor1(arrdiv32_fs953_xor1), .fs_or0(arrdiv32_fs953_or0));
  fs fs_arrdiv32_fs954_out(.a(arrdiv32_mux2to1893_xor0[0]), .b(b[26]), .bin(arrdiv32_fs953_or0[0]), .fs_xor1(arrdiv32_fs954_xor1), .fs_or0(arrdiv32_fs954_or0));
  fs fs_arrdiv32_fs955_out(.a(arrdiv32_mux2to1894_xor0[0]), .b(b[27]), .bin(arrdiv32_fs954_or0[0]), .fs_xor1(arrdiv32_fs955_xor1), .fs_or0(arrdiv32_fs955_or0));
  fs fs_arrdiv32_fs956_out(.a(arrdiv32_mux2to1895_xor0[0]), .b(b[28]), .bin(arrdiv32_fs955_or0[0]), .fs_xor1(arrdiv32_fs956_xor1), .fs_or0(arrdiv32_fs956_or0));
  fs fs_arrdiv32_fs957_out(.a(arrdiv32_mux2to1896_xor0[0]), .b(b[29]), .bin(arrdiv32_fs956_or0[0]), .fs_xor1(arrdiv32_fs957_xor1), .fs_or0(arrdiv32_fs957_or0));
  fs fs_arrdiv32_fs958_out(.a(arrdiv32_mux2to1897_xor0[0]), .b(b[30]), .bin(arrdiv32_fs957_or0[0]), .fs_xor1(arrdiv32_fs958_xor1), .fs_or0(arrdiv32_fs958_or0));
  fs fs_arrdiv32_fs959_out(.a(arrdiv32_mux2to1898_xor0[0]), .b(b[31]), .bin(arrdiv32_fs958_or0[0]), .fs_xor1(arrdiv32_fs959_xor1), .fs_or0(arrdiv32_fs959_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1899_out(.d0(arrdiv32_fs928_xor0[0]), .d1(a[2]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1899_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1900_out(.d0(arrdiv32_fs929_xor1[0]), .d1(arrdiv32_mux2to1868_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1900_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1901_out(.d0(arrdiv32_fs930_xor1[0]), .d1(arrdiv32_mux2to1869_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1901_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1902_out(.d0(arrdiv32_fs931_xor1[0]), .d1(arrdiv32_mux2to1870_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1902_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1903_out(.d0(arrdiv32_fs932_xor1[0]), .d1(arrdiv32_mux2to1871_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1903_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1904_out(.d0(arrdiv32_fs933_xor1[0]), .d1(arrdiv32_mux2to1872_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1904_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1905_out(.d0(arrdiv32_fs934_xor1[0]), .d1(arrdiv32_mux2to1873_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1905_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1906_out(.d0(arrdiv32_fs935_xor1[0]), .d1(arrdiv32_mux2to1874_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1906_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1907_out(.d0(arrdiv32_fs936_xor1[0]), .d1(arrdiv32_mux2to1875_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1907_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1908_out(.d0(arrdiv32_fs937_xor1[0]), .d1(arrdiv32_mux2to1876_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1908_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1909_out(.d0(arrdiv32_fs938_xor1[0]), .d1(arrdiv32_mux2to1877_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1909_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1910_out(.d0(arrdiv32_fs939_xor1[0]), .d1(arrdiv32_mux2to1878_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1910_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1911_out(.d0(arrdiv32_fs940_xor1[0]), .d1(arrdiv32_mux2to1879_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1911_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1912_out(.d0(arrdiv32_fs941_xor1[0]), .d1(arrdiv32_mux2to1880_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1912_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1913_out(.d0(arrdiv32_fs942_xor1[0]), .d1(arrdiv32_mux2to1881_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1913_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1914_out(.d0(arrdiv32_fs943_xor1[0]), .d1(arrdiv32_mux2to1882_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1914_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1915_out(.d0(arrdiv32_fs944_xor1[0]), .d1(arrdiv32_mux2to1883_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1915_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1916_out(.d0(arrdiv32_fs945_xor1[0]), .d1(arrdiv32_mux2to1884_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1916_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1917_out(.d0(arrdiv32_fs946_xor1[0]), .d1(arrdiv32_mux2to1885_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1917_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1918_out(.d0(arrdiv32_fs947_xor1[0]), .d1(arrdiv32_mux2to1886_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1918_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1919_out(.d0(arrdiv32_fs948_xor1[0]), .d1(arrdiv32_mux2to1887_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1919_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1920_out(.d0(arrdiv32_fs949_xor1[0]), .d1(arrdiv32_mux2to1888_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1920_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1921_out(.d0(arrdiv32_fs950_xor1[0]), .d1(arrdiv32_mux2to1889_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1921_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1922_out(.d0(arrdiv32_fs951_xor1[0]), .d1(arrdiv32_mux2to1890_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1922_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1923_out(.d0(arrdiv32_fs952_xor1[0]), .d1(arrdiv32_mux2to1891_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1923_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1924_out(.d0(arrdiv32_fs953_xor1[0]), .d1(arrdiv32_mux2to1892_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1924_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1925_out(.d0(arrdiv32_fs954_xor1[0]), .d1(arrdiv32_mux2to1893_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1925_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1926_out(.d0(arrdiv32_fs955_xor1[0]), .d1(arrdiv32_mux2to1894_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1926_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1927_out(.d0(arrdiv32_fs956_xor1[0]), .d1(arrdiv32_mux2to1895_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1927_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1928_out(.d0(arrdiv32_fs957_xor1[0]), .d1(arrdiv32_mux2to1896_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1928_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1929_out(.d0(arrdiv32_fs958_xor1[0]), .d1(arrdiv32_mux2to1897_xor0[0]), .sel(arrdiv32_fs959_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1929_xor0));
  not_gate not_gate_arrdiv32_not29(.a(arrdiv32_fs959_or0[0]), .out(arrdiv32_not29));
  fs fs_arrdiv32_fs960_out(.a(a[1]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs960_xor0), .fs_or0(arrdiv32_fs960_and0));
  fs fs_arrdiv32_fs961_out(.a(arrdiv32_mux2to1899_xor0[0]), .b(b[1]), .bin(arrdiv32_fs960_and0[0]), .fs_xor1(arrdiv32_fs961_xor1), .fs_or0(arrdiv32_fs961_or0));
  fs fs_arrdiv32_fs962_out(.a(arrdiv32_mux2to1900_xor0[0]), .b(b[2]), .bin(arrdiv32_fs961_or0[0]), .fs_xor1(arrdiv32_fs962_xor1), .fs_or0(arrdiv32_fs962_or0));
  fs fs_arrdiv32_fs963_out(.a(arrdiv32_mux2to1901_xor0[0]), .b(b[3]), .bin(arrdiv32_fs962_or0[0]), .fs_xor1(arrdiv32_fs963_xor1), .fs_or0(arrdiv32_fs963_or0));
  fs fs_arrdiv32_fs964_out(.a(arrdiv32_mux2to1902_xor0[0]), .b(b[4]), .bin(arrdiv32_fs963_or0[0]), .fs_xor1(arrdiv32_fs964_xor1), .fs_or0(arrdiv32_fs964_or0));
  fs fs_arrdiv32_fs965_out(.a(arrdiv32_mux2to1903_xor0[0]), .b(b[5]), .bin(arrdiv32_fs964_or0[0]), .fs_xor1(arrdiv32_fs965_xor1), .fs_or0(arrdiv32_fs965_or0));
  fs fs_arrdiv32_fs966_out(.a(arrdiv32_mux2to1904_xor0[0]), .b(b[6]), .bin(arrdiv32_fs965_or0[0]), .fs_xor1(arrdiv32_fs966_xor1), .fs_or0(arrdiv32_fs966_or0));
  fs fs_arrdiv32_fs967_out(.a(arrdiv32_mux2to1905_xor0[0]), .b(b[7]), .bin(arrdiv32_fs966_or0[0]), .fs_xor1(arrdiv32_fs967_xor1), .fs_or0(arrdiv32_fs967_or0));
  fs fs_arrdiv32_fs968_out(.a(arrdiv32_mux2to1906_xor0[0]), .b(b[8]), .bin(arrdiv32_fs967_or0[0]), .fs_xor1(arrdiv32_fs968_xor1), .fs_or0(arrdiv32_fs968_or0));
  fs fs_arrdiv32_fs969_out(.a(arrdiv32_mux2to1907_xor0[0]), .b(b[9]), .bin(arrdiv32_fs968_or0[0]), .fs_xor1(arrdiv32_fs969_xor1), .fs_or0(arrdiv32_fs969_or0));
  fs fs_arrdiv32_fs970_out(.a(arrdiv32_mux2to1908_xor0[0]), .b(b[10]), .bin(arrdiv32_fs969_or0[0]), .fs_xor1(arrdiv32_fs970_xor1), .fs_or0(arrdiv32_fs970_or0));
  fs fs_arrdiv32_fs971_out(.a(arrdiv32_mux2to1909_xor0[0]), .b(b[11]), .bin(arrdiv32_fs970_or0[0]), .fs_xor1(arrdiv32_fs971_xor1), .fs_or0(arrdiv32_fs971_or0));
  fs fs_arrdiv32_fs972_out(.a(arrdiv32_mux2to1910_xor0[0]), .b(b[12]), .bin(arrdiv32_fs971_or0[0]), .fs_xor1(arrdiv32_fs972_xor1), .fs_or0(arrdiv32_fs972_or0));
  fs fs_arrdiv32_fs973_out(.a(arrdiv32_mux2to1911_xor0[0]), .b(b[13]), .bin(arrdiv32_fs972_or0[0]), .fs_xor1(arrdiv32_fs973_xor1), .fs_or0(arrdiv32_fs973_or0));
  fs fs_arrdiv32_fs974_out(.a(arrdiv32_mux2to1912_xor0[0]), .b(b[14]), .bin(arrdiv32_fs973_or0[0]), .fs_xor1(arrdiv32_fs974_xor1), .fs_or0(arrdiv32_fs974_or0));
  fs fs_arrdiv32_fs975_out(.a(arrdiv32_mux2to1913_xor0[0]), .b(b[15]), .bin(arrdiv32_fs974_or0[0]), .fs_xor1(arrdiv32_fs975_xor1), .fs_or0(arrdiv32_fs975_or0));
  fs fs_arrdiv32_fs976_out(.a(arrdiv32_mux2to1914_xor0[0]), .b(b[16]), .bin(arrdiv32_fs975_or0[0]), .fs_xor1(arrdiv32_fs976_xor1), .fs_or0(arrdiv32_fs976_or0));
  fs fs_arrdiv32_fs977_out(.a(arrdiv32_mux2to1915_xor0[0]), .b(b[17]), .bin(arrdiv32_fs976_or0[0]), .fs_xor1(arrdiv32_fs977_xor1), .fs_or0(arrdiv32_fs977_or0));
  fs fs_arrdiv32_fs978_out(.a(arrdiv32_mux2to1916_xor0[0]), .b(b[18]), .bin(arrdiv32_fs977_or0[0]), .fs_xor1(arrdiv32_fs978_xor1), .fs_or0(arrdiv32_fs978_or0));
  fs fs_arrdiv32_fs979_out(.a(arrdiv32_mux2to1917_xor0[0]), .b(b[19]), .bin(arrdiv32_fs978_or0[0]), .fs_xor1(arrdiv32_fs979_xor1), .fs_or0(arrdiv32_fs979_or0));
  fs fs_arrdiv32_fs980_out(.a(arrdiv32_mux2to1918_xor0[0]), .b(b[20]), .bin(arrdiv32_fs979_or0[0]), .fs_xor1(arrdiv32_fs980_xor1), .fs_or0(arrdiv32_fs980_or0));
  fs fs_arrdiv32_fs981_out(.a(arrdiv32_mux2to1919_xor0[0]), .b(b[21]), .bin(arrdiv32_fs980_or0[0]), .fs_xor1(arrdiv32_fs981_xor1), .fs_or0(arrdiv32_fs981_or0));
  fs fs_arrdiv32_fs982_out(.a(arrdiv32_mux2to1920_xor0[0]), .b(b[22]), .bin(arrdiv32_fs981_or0[0]), .fs_xor1(arrdiv32_fs982_xor1), .fs_or0(arrdiv32_fs982_or0));
  fs fs_arrdiv32_fs983_out(.a(arrdiv32_mux2to1921_xor0[0]), .b(b[23]), .bin(arrdiv32_fs982_or0[0]), .fs_xor1(arrdiv32_fs983_xor1), .fs_or0(arrdiv32_fs983_or0));
  fs fs_arrdiv32_fs984_out(.a(arrdiv32_mux2to1922_xor0[0]), .b(b[24]), .bin(arrdiv32_fs983_or0[0]), .fs_xor1(arrdiv32_fs984_xor1), .fs_or0(arrdiv32_fs984_or0));
  fs fs_arrdiv32_fs985_out(.a(arrdiv32_mux2to1923_xor0[0]), .b(b[25]), .bin(arrdiv32_fs984_or0[0]), .fs_xor1(arrdiv32_fs985_xor1), .fs_or0(arrdiv32_fs985_or0));
  fs fs_arrdiv32_fs986_out(.a(arrdiv32_mux2to1924_xor0[0]), .b(b[26]), .bin(arrdiv32_fs985_or0[0]), .fs_xor1(arrdiv32_fs986_xor1), .fs_or0(arrdiv32_fs986_or0));
  fs fs_arrdiv32_fs987_out(.a(arrdiv32_mux2to1925_xor0[0]), .b(b[27]), .bin(arrdiv32_fs986_or0[0]), .fs_xor1(arrdiv32_fs987_xor1), .fs_or0(arrdiv32_fs987_or0));
  fs fs_arrdiv32_fs988_out(.a(arrdiv32_mux2to1926_xor0[0]), .b(b[28]), .bin(arrdiv32_fs987_or0[0]), .fs_xor1(arrdiv32_fs988_xor1), .fs_or0(arrdiv32_fs988_or0));
  fs fs_arrdiv32_fs989_out(.a(arrdiv32_mux2to1927_xor0[0]), .b(b[29]), .bin(arrdiv32_fs988_or0[0]), .fs_xor1(arrdiv32_fs989_xor1), .fs_or0(arrdiv32_fs989_or0));
  fs fs_arrdiv32_fs990_out(.a(arrdiv32_mux2to1928_xor0[0]), .b(b[30]), .bin(arrdiv32_fs989_or0[0]), .fs_xor1(arrdiv32_fs990_xor1), .fs_or0(arrdiv32_fs990_or0));
  fs fs_arrdiv32_fs991_out(.a(arrdiv32_mux2to1929_xor0[0]), .b(b[31]), .bin(arrdiv32_fs990_or0[0]), .fs_xor1(arrdiv32_fs991_xor1), .fs_or0(arrdiv32_fs991_or0));
  mux2to1 mux2to1_arrdiv32_mux2to1930_out(.d0(arrdiv32_fs960_xor0[0]), .d1(a[1]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1930_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1931_out(.d0(arrdiv32_fs961_xor1[0]), .d1(arrdiv32_mux2to1899_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1931_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1932_out(.d0(arrdiv32_fs962_xor1[0]), .d1(arrdiv32_mux2to1900_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1932_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1933_out(.d0(arrdiv32_fs963_xor1[0]), .d1(arrdiv32_mux2to1901_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1933_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1934_out(.d0(arrdiv32_fs964_xor1[0]), .d1(arrdiv32_mux2to1902_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1934_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1935_out(.d0(arrdiv32_fs965_xor1[0]), .d1(arrdiv32_mux2to1903_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1935_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1936_out(.d0(arrdiv32_fs966_xor1[0]), .d1(arrdiv32_mux2to1904_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1936_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1937_out(.d0(arrdiv32_fs967_xor1[0]), .d1(arrdiv32_mux2to1905_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1937_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1938_out(.d0(arrdiv32_fs968_xor1[0]), .d1(arrdiv32_mux2to1906_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1938_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1939_out(.d0(arrdiv32_fs969_xor1[0]), .d1(arrdiv32_mux2to1907_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1939_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1940_out(.d0(arrdiv32_fs970_xor1[0]), .d1(arrdiv32_mux2to1908_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1940_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1941_out(.d0(arrdiv32_fs971_xor1[0]), .d1(arrdiv32_mux2to1909_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1941_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1942_out(.d0(arrdiv32_fs972_xor1[0]), .d1(arrdiv32_mux2to1910_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1942_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1943_out(.d0(arrdiv32_fs973_xor1[0]), .d1(arrdiv32_mux2to1911_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1943_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1944_out(.d0(arrdiv32_fs974_xor1[0]), .d1(arrdiv32_mux2to1912_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1944_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1945_out(.d0(arrdiv32_fs975_xor1[0]), .d1(arrdiv32_mux2to1913_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1945_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1946_out(.d0(arrdiv32_fs976_xor1[0]), .d1(arrdiv32_mux2to1914_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1946_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1947_out(.d0(arrdiv32_fs977_xor1[0]), .d1(arrdiv32_mux2to1915_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1947_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1948_out(.d0(arrdiv32_fs978_xor1[0]), .d1(arrdiv32_mux2to1916_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1948_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1949_out(.d0(arrdiv32_fs979_xor1[0]), .d1(arrdiv32_mux2to1917_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1949_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1950_out(.d0(arrdiv32_fs980_xor1[0]), .d1(arrdiv32_mux2to1918_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1950_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1951_out(.d0(arrdiv32_fs981_xor1[0]), .d1(arrdiv32_mux2to1919_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1951_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1952_out(.d0(arrdiv32_fs982_xor1[0]), .d1(arrdiv32_mux2to1920_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1952_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1953_out(.d0(arrdiv32_fs983_xor1[0]), .d1(arrdiv32_mux2to1921_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1953_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1954_out(.d0(arrdiv32_fs984_xor1[0]), .d1(arrdiv32_mux2to1922_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1954_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1955_out(.d0(arrdiv32_fs985_xor1[0]), .d1(arrdiv32_mux2to1923_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1955_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1956_out(.d0(arrdiv32_fs986_xor1[0]), .d1(arrdiv32_mux2to1924_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1956_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1957_out(.d0(arrdiv32_fs987_xor1[0]), .d1(arrdiv32_mux2to1925_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1957_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1958_out(.d0(arrdiv32_fs988_xor1[0]), .d1(arrdiv32_mux2to1926_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1958_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1959_out(.d0(arrdiv32_fs989_xor1[0]), .d1(arrdiv32_mux2to1927_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1959_xor0));
  mux2to1 mux2to1_arrdiv32_mux2to1960_out(.d0(arrdiv32_fs990_xor1[0]), .d1(arrdiv32_mux2to1928_xor0[0]), .sel(arrdiv32_fs991_or0[0]), .mux2to1_xor0(arrdiv32_mux2to1960_xor0));
  not_gate not_gate_arrdiv32_not30(.a(arrdiv32_fs991_or0[0]), .out(arrdiv32_not30));
  fs fs_arrdiv32_fs992_out(.a(a[0]), .b(b[0]), .bin(1'b0), .fs_xor1(arrdiv32_fs992_xor0), .fs_or0(arrdiv32_fs992_and0));
  fs fs_arrdiv32_fs993_out(.a(arrdiv32_mux2to1930_xor0[0]), .b(b[1]), .bin(arrdiv32_fs992_and0[0]), .fs_xor1(arrdiv32_fs993_xor1), .fs_or0(arrdiv32_fs993_or0));
  fs fs_arrdiv32_fs994_out(.a(arrdiv32_mux2to1931_xor0[0]), .b(b[2]), .bin(arrdiv32_fs993_or0[0]), .fs_xor1(arrdiv32_fs994_xor1), .fs_or0(arrdiv32_fs994_or0));
  fs fs_arrdiv32_fs995_out(.a(arrdiv32_mux2to1932_xor0[0]), .b(b[3]), .bin(arrdiv32_fs994_or0[0]), .fs_xor1(arrdiv32_fs995_xor1), .fs_or0(arrdiv32_fs995_or0));
  fs fs_arrdiv32_fs996_out(.a(arrdiv32_mux2to1933_xor0[0]), .b(b[4]), .bin(arrdiv32_fs995_or0[0]), .fs_xor1(arrdiv32_fs996_xor1), .fs_or0(arrdiv32_fs996_or0));
  fs fs_arrdiv32_fs997_out(.a(arrdiv32_mux2to1934_xor0[0]), .b(b[5]), .bin(arrdiv32_fs996_or0[0]), .fs_xor1(arrdiv32_fs997_xor1), .fs_or0(arrdiv32_fs997_or0));
  fs fs_arrdiv32_fs998_out(.a(arrdiv32_mux2to1935_xor0[0]), .b(b[6]), .bin(arrdiv32_fs997_or0[0]), .fs_xor1(arrdiv32_fs998_xor1), .fs_or0(arrdiv32_fs998_or0));
  fs fs_arrdiv32_fs999_out(.a(arrdiv32_mux2to1936_xor0[0]), .b(b[7]), .bin(arrdiv32_fs998_or0[0]), .fs_xor1(arrdiv32_fs999_xor1), .fs_or0(arrdiv32_fs999_or0));
  fs fs_arrdiv32_fs1000_out(.a(arrdiv32_mux2to1937_xor0[0]), .b(b[8]), .bin(arrdiv32_fs999_or0[0]), .fs_xor1(arrdiv32_fs1000_xor1), .fs_or0(arrdiv32_fs1000_or0));
  fs fs_arrdiv32_fs1001_out(.a(arrdiv32_mux2to1938_xor0[0]), .b(b[9]), .bin(arrdiv32_fs1000_or0[0]), .fs_xor1(arrdiv32_fs1001_xor1), .fs_or0(arrdiv32_fs1001_or0));
  fs fs_arrdiv32_fs1002_out(.a(arrdiv32_mux2to1939_xor0[0]), .b(b[10]), .bin(arrdiv32_fs1001_or0[0]), .fs_xor1(arrdiv32_fs1002_xor1), .fs_or0(arrdiv32_fs1002_or0));
  fs fs_arrdiv32_fs1003_out(.a(arrdiv32_mux2to1940_xor0[0]), .b(b[11]), .bin(arrdiv32_fs1002_or0[0]), .fs_xor1(arrdiv32_fs1003_xor1), .fs_or0(arrdiv32_fs1003_or0));
  fs fs_arrdiv32_fs1004_out(.a(arrdiv32_mux2to1941_xor0[0]), .b(b[12]), .bin(arrdiv32_fs1003_or0[0]), .fs_xor1(arrdiv32_fs1004_xor1), .fs_or0(arrdiv32_fs1004_or0));
  fs fs_arrdiv32_fs1005_out(.a(arrdiv32_mux2to1942_xor0[0]), .b(b[13]), .bin(arrdiv32_fs1004_or0[0]), .fs_xor1(arrdiv32_fs1005_xor1), .fs_or0(arrdiv32_fs1005_or0));
  fs fs_arrdiv32_fs1006_out(.a(arrdiv32_mux2to1943_xor0[0]), .b(b[14]), .bin(arrdiv32_fs1005_or0[0]), .fs_xor1(arrdiv32_fs1006_xor1), .fs_or0(arrdiv32_fs1006_or0));
  fs fs_arrdiv32_fs1007_out(.a(arrdiv32_mux2to1944_xor0[0]), .b(b[15]), .bin(arrdiv32_fs1006_or0[0]), .fs_xor1(arrdiv32_fs1007_xor1), .fs_or0(arrdiv32_fs1007_or0));
  fs fs_arrdiv32_fs1008_out(.a(arrdiv32_mux2to1945_xor0[0]), .b(b[16]), .bin(arrdiv32_fs1007_or0[0]), .fs_xor1(arrdiv32_fs1008_xor1), .fs_or0(arrdiv32_fs1008_or0));
  fs fs_arrdiv32_fs1009_out(.a(arrdiv32_mux2to1946_xor0[0]), .b(b[17]), .bin(arrdiv32_fs1008_or0[0]), .fs_xor1(arrdiv32_fs1009_xor1), .fs_or0(arrdiv32_fs1009_or0));
  fs fs_arrdiv32_fs1010_out(.a(arrdiv32_mux2to1947_xor0[0]), .b(b[18]), .bin(arrdiv32_fs1009_or0[0]), .fs_xor1(arrdiv32_fs1010_xor1), .fs_or0(arrdiv32_fs1010_or0));
  fs fs_arrdiv32_fs1011_out(.a(arrdiv32_mux2to1948_xor0[0]), .b(b[19]), .bin(arrdiv32_fs1010_or0[0]), .fs_xor1(arrdiv32_fs1011_xor1), .fs_or0(arrdiv32_fs1011_or0));
  fs fs_arrdiv32_fs1012_out(.a(arrdiv32_mux2to1949_xor0[0]), .b(b[20]), .bin(arrdiv32_fs1011_or0[0]), .fs_xor1(arrdiv32_fs1012_xor1), .fs_or0(arrdiv32_fs1012_or0));
  fs fs_arrdiv32_fs1013_out(.a(arrdiv32_mux2to1950_xor0[0]), .b(b[21]), .bin(arrdiv32_fs1012_or0[0]), .fs_xor1(arrdiv32_fs1013_xor1), .fs_or0(arrdiv32_fs1013_or0));
  fs fs_arrdiv32_fs1014_out(.a(arrdiv32_mux2to1951_xor0[0]), .b(b[22]), .bin(arrdiv32_fs1013_or0[0]), .fs_xor1(arrdiv32_fs1014_xor1), .fs_or0(arrdiv32_fs1014_or0));
  fs fs_arrdiv32_fs1015_out(.a(arrdiv32_mux2to1952_xor0[0]), .b(b[23]), .bin(arrdiv32_fs1014_or0[0]), .fs_xor1(arrdiv32_fs1015_xor1), .fs_or0(arrdiv32_fs1015_or0));
  fs fs_arrdiv32_fs1016_out(.a(arrdiv32_mux2to1953_xor0[0]), .b(b[24]), .bin(arrdiv32_fs1015_or0[0]), .fs_xor1(arrdiv32_fs1016_xor1), .fs_or0(arrdiv32_fs1016_or0));
  fs fs_arrdiv32_fs1017_out(.a(arrdiv32_mux2to1954_xor0[0]), .b(b[25]), .bin(arrdiv32_fs1016_or0[0]), .fs_xor1(arrdiv32_fs1017_xor1), .fs_or0(arrdiv32_fs1017_or0));
  fs fs_arrdiv32_fs1018_out(.a(arrdiv32_mux2to1955_xor0[0]), .b(b[26]), .bin(arrdiv32_fs1017_or0[0]), .fs_xor1(arrdiv32_fs1018_xor1), .fs_or0(arrdiv32_fs1018_or0));
  fs fs_arrdiv32_fs1019_out(.a(arrdiv32_mux2to1956_xor0[0]), .b(b[27]), .bin(arrdiv32_fs1018_or0[0]), .fs_xor1(arrdiv32_fs1019_xor1), .fs_or0(arrdiv32_fs1019_or0));
  fs fs_arrdiv32_fs1020_out(.a(arrdiv32_mux2to1957_xor0[0]), .b(b[28]), .bin(arrdiv32_fs1019_or0[0]), .fs_xor1(arrdiv32_fs1020_xor1), .fs_or0(arrdiv32_fs1020_or0));
  fs fs_arrdiv32_fs1021_out(.a(arrdiv32_mux2to1958_xor0[0]), .b(b[29]), .bin(arrdiv32_fs1020_or0[0]), .fs_xor1(arrdiv32_fs1021_xor1), .fs_or0(arrdiv32_fs1021_or0));
  fs fs_arrdiv32_fs1022_out(.a(arrdiv32_mux2to1959_xor0[0]), .b(b[30]), .bin(arrdiv32_fs1021_or0[0]), .fs_xor1(arrdiv32_fs1022_xor1), .fs_or0(arrdiv32_fs1022_or0));
  fs fs_arrdiv32_fs1023_out(.a(arrdiv32_mux2to1960_xor0[0]), .b(b[31]), .bin(arrdiv32_fs1022_or0[0]), .fs_xor1(arrdiv32_fs1023_xor1), .fs_or0(arrdiv32_fs1023_or0));
  not_gate not_gate_arrdiv32_not31(.a(arrdiv32_fs1023_or0[0]), .out(arrdiv32_not31));

  assign arrdiv32_out[0] = arrdiv32_not31[0];
  assign arrdiv32_out[1] = arrdiv32_not30[0];
  assign arrdiv32_out[2] = arrdiv32_not29[0];
  assign arrdiv32_out[3] = arrdiv32_not28[0];
  assign arrdiv32_out[4] = arrdiv32_not27[0];
  assign arrdiv32_out[5] = arrdiv32_not26[0];
  assign arrdiv32_out[6] = arrdiv32_not25[0];
  assign arrdiv32_out[7] = arrdiv32_not24[0];
  assign arrdiv32_out[8] = arrdiv32_not23[0];
  assign arrdiv32_out[9] = arrdiv32_not22[0];
  assign arrdiv32_out[10] = arrdiv32_not21[0];
  assign arrdiv32_out[11] = arrdiv32_not20[0];
  assign arrdiv32_out[12] = arrdiv32_not19[0];
  assign arrdiv32_out[13] = arrdiv32_not18[0];
  assign arrdiv32_out[14] = arrdiv32_not17[0];
  assign arrdiv32_out[15] = arrdiv32_not16[0];
  assign arrdiv32_out[16] = arrdiv32_not15[0];
  assign arrdiv32_out[17] = arrdiv32_not14[0];
  assign arrdiv32_out[18] = arrdiv32_not13[0];
  assign arrdiv32_out[19] = arrdiv32_not12[0];
  assign arrdiv32_out[20] = arrdiv32_not11[0];
  assign arrdiv32_out[21] = arrdiv32_not10[0];
  assign arrdiv32_out[22] = arrdiv32_not9[0];
  assign arrdiv32_out[23] = arrdiv32_not8[0];
  assign arrdiv32_out[24] = arrdiv32_not7[0];
  assign arrdiv32_out[25] = arrdiv32_not6[0];
  assign arrdiv32_out[26] = arrdiv32_not5[0];
  assign arrdiv32_out[27] = arrdiv32_not4[0];
  assign arrdiv32_out[28] = arrdiv32_not3[0];
  assign arrdiv32_out[29] = arrdiv32_not2[0];
  assign arrdiv32_out[30] = arrdiv32_not1[0];
  assign arrdiv32_out[31] = arrdiv32_not0[0];
endmodule