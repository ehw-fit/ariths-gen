module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(a[0], b[0], ha_xor0);
  and_gate and_gate_ha_and0(a[0], b[0], ha_and0);
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(a[0], b[0], fa_xor0);
  and_gate and_gate_fa_and0(a[0], b[0], fa_and0);
  xor_gate xor_gate_fa_xor1(fa_xor0[0], cin[0], fa_xor1);
  and_gate and_gate_fa_and1(fa_xor0[0], cin[0], fa_and1);
  or_gate or_gate_fa_or0(fa_and0[0], fa_and1[0], fa_or0);
endmodule

module h_u_arrmul24(input [23:0] a, input [23:0] b, output [47:0] h_u_arrmul24_out);
  wire [0:0] h_u_arrmul24_and0_0;
  wire [0:0] h_u_arrmul24_and1_0;
  wire [0:0] h_u_arrmul24_and2_0;
  wire [0:0] h_u_arrmul24_and3_0;
  wire [0:0] h_u_arrmul24_and4_0;
  wire [0:0] h_u_arrmul24_and5_0;
  wire [0:0] h_u_arrmul24_and6_0;
  wire [0:0] h_u_arrmul24_and7_0;
  wire [0:0] h_u_arrmul24_and8_0;
  wire [0:0] h_u_arrmul24_and9_0;
  wire [0:0] h_u_arrmul24_and10_0;
  wire [0:0] h_u_arrmul24_and11_0;
  wire [0:0] h_u_arrmul24_and12_0;
  wire [0:0] h_u_arrmul24_and13_0;
  wire [0:0] h_u_arrmul24_and14_0;
  wire [0:0] h_u_arrmul24_and15_0;
  wire [0:0] h_u_arrmul24_and16_0;
  wire [0:0] h_u_arrmul24_and17_0;
  wire [0:0] h_u_arrmul24_and18_0;
  wire [0:0] h_u_arrmul24_and19_0;
  wire [0:0] h_u_arrmul24_and20_0;
  wire [0:0] h_u_arrmul24_and21_0;
  wire [0:0] h_u_arrmul24_and22_0;
  wire [0:0] h_u_arrmul24_and23_0;
  wire [0:0] h_u_arrmul24_and0_1;
  wire [0:0] h_u_arrmul24_ha0_1_xor0;
  wire [0:0] h_u_arrmul24_ha0_1_and0;
  wire [0:0] h_u_arrmul24_and1_1;
  wire [0:0] h_u_arrmul24_fa1_1_xor1;
  wire [0:0] h_u_arrmul24_fa1_1_or0;
  wire [0:0] h_u_arrmul24_and2_1;
  wire [0:0] h_u_arrmul24_fa2_1_xor1;
  wire [0:0] h_u_arrmul24_fa2_1_or0;
  wire [0:0] h_u_arrmul24_and3_1;
  wire [0:0] h_u_arrmul24_fa3_1_xor1;
  wire [0:0] h_u_arrmul24_fa3_1_or0;
  wire [0:0] h_u_arrmul24_and4_1;
  wire [0:0] h_u_arrmul24_fa4_1_xor1;
  wire [0:0] h_u_arrmul24_fa4_1_or0;
  wire [0:0] h_u_arrmul24_and5_1;
  wire [0:0] h_u_arrmul24_fa5_1_xor1;
  wire [0:0] h_u_arrmul24_fa5_1_or0;
  wire [0:0] h_u_arrmul24_and6_1;
  wire [0:0] h_u_arrmul24_fa6_1_xor1;
  wire [0:0] h_u_arrmul24_fa6_1_or0;
  wire [0:0] h_u_arrmul24_and7_1;
  wire [0:0] h_u_arrmul24_fa7_1_xor1;
  wire [0:0] h_u_arrmul24_fa7_1_or0;
  wire [0:0] h_u_arrmul24_and8_1;
  wire [0:0] h_u_arrmul24_fa8_1_xor1;
  wire [0:0] h_u_arrmul24_fa8_1_or0;
  wire [0:0] h_u_arrmul24_and9_1;
  wire [0:0] h_u_arrmul24_fa9_1_xor1;
  wire [0:0] h_u_arrmul24_fa9_1_or0;
  wire [0:0] h_u_arrmul24_and10_1;
  wire [0:0] h_u_arrmul24_fa10_1_xor1;
  wire [0:0] h_u_arrmul24_fa10_1_or0;
  wire [0:0] h_u_arrmul24_and11_1;
  wire [0:0] h_u_arrmul24_fa11_1_xor1;
  wire [0:0] h_u_arrmul24_fa11_1_or0;
  wire [0:0] h_u_arrmul24_and12_1;
  wire [0:0] h_u_arrmul24_fa12_1_xor1;
  wire [0:0] h_u_arrmul24_fa12_1_or0;
  wire [0:0] h_u_arrmul24_and13_1;
  wire [0:0] h_u_arrmul24_fa13_1_xor1;
  wire [0:0] h_u_arrmul24_fa13_1_or0;
  wire [0:0] h_u_arrmul24_and14_1;
  wire [0:0] h_u_arrmul24_fa14_1_xor1;
  wire [0:0] h_u_arrmul24_fa14_1_or0;
  wire [0:0] h_u_arrmul24_and15_1;
  wire [0:0] h_u_arrmul24_fa15_1_xor1;
  wire [0:0] h_u_arrmul24_fa15_1_or0;
  wire [0:0] h_u_arrmul24_and16_1;
  wire [0:0] h_u_arrmul24_fa16_1_xor1;
  wire [0:0] h_u_arrmul24_fa16_1_or0;
  wire [0:0] h_u_arrmul24_and17_1;
  wire [0:0] h_u_arrmul24_fa17_1_xor1;
  wire [0:0] h_u_arrmul24_fa17_1_or0;
  wire [0:0] h_u_arrmul24_and18_1;
  wire [0:0] h_u_arrmul24_fa18_1_xor1;
  wire [0:0] h_u_arrmul24_fa18_1_or0;
  wire [0:0] h_u_arrmul24_and19_1;
  wire [0:0] h_u_arrmul24_fa19_1_xor1;
  wire [0:0] h_u_arrmul24_fa19_1_or0;
  wire [0:0] h_u_arrmul24_and20_1;
  wire [0:0] h_u_arrmul24_fa20_1_xor1;
  wire [0:0] h_u_arrmul24_fa20_1_or0;
  wire [0:0] h_u_arrmul24_and21_1;
  wire [0:0] h_u_arrmul24_fa21_1_xor1;
  wire [0:0] h_u_arrmul24_fa21_1_or0;
  wire [0:0] h_u_arrmul24_and22_1;
  wire [0:0] h_u_arrmul24_fa22_1_xor1;
  wire [0:0] h_u_arrmul24_fa22_1_or0;
  wire [0:0] h_u_arrmul24_and23_1;
  wire [0:0] h_u_arrmul24_ha23_1_xor0;
  wire [0:0] h_u_arrmul24_ha23_1_and0;
  wire [0:0] h_u_arrmul24_and0_2;
  wire [0:0] h_u_arrmul24_ha0_2_xor0;
  wire [0:0] h_u_arrmul24_ha0_2_and0;
  wire [0:0] h_u_arrmul24_and1_2;
  wire [0:0] h_u_arrmul24_fa1_2_xor1;
  wire [0:0] h_u_arrmul24_fa1_2_or0;
  wire [0:0] h_u_arrmul24_and2_2;
  wire [0:0] h_u_arrmul24_fa2_2_xor1;
  wire [0:0] h_u_arrmul24_fa2_2_or0;
  wire [0:0] h_u_arrmul24_and3_2;
  wire [0:0] h_u_arrmul24_fa3_2_xor1;
  wire [0:0] h_u_arrmul24_fa3_2_or0;
  wire [0:0] h_u_arrmul24_and4_2;
  wire [0:0] h_u_arrmul24_fa4_2_xor1;
  wire [0:0] h_u_arrmul24_fa4_2_or0;
  wire [0:0] h_u_arrmul24_and5_2;
  wire [0:0] h_u_arrmul24_fa5_2_xor1;
  wire [0:0] h_u_arrmul24_fa5_2_or0;
  wire [0:0] h_u_arrmul24_and6_2;
  wire [0:0] h_u_arrmul24_fa6_2_xor1;
  wire [0:0] h_u_arrmul24_fa6_2_or0;
  wire [0:0] h_u_arrmul24_and7_2;
  wire [0:0] h_u_arrmul24_fa7_2_xor1;
  wire [0:0] h_u_arrmul24_fa7_2_or0;
  wire [0:0] h_u_arrmul24_and8_2;
  wire [0:0] h_u_arrmul24_fa8_2_xor1;
  wire [0:0] h_u_arrmul24_fa8_2_or0;
  wire [0:0] h_u_arrmul24_and9_2;
  wire [0:0] h_u_arrmul24_fa9_2_xor1;
  wire [0:0] h_u_arrmul24_fa9_2_or0;
  wire [0:0] h_u_arrmul24_and10_2;
  wire [0:0] h_u_arrmul24_fa10_2_xor1;
  wire [0:0] h_u_arrmul24_fa10_2_or0;
  wire [0:0] h_u_arrmul24_and11_2;
  wire [0:0] h_u_arrmul24_fa11_2_xor1;
  wire [0:0] h_u_arrmul24_fa11_2_or0;
  wire [0:0] h_u_arrmul24_and12_2;
  wire [0:0] h_u_arrmul24_fa12_2_xor1;
  wire [0:0] h_u_arrmul24_fa12_2_or0;
  wire [0:0] h_u_arrmul24_and13_2;
  wire [0:0] h_u_arrmul24_fa13_2_xor1;
  wire [0:0] h_u_arrmul24_fa13_2_or0;
  wire [0:0] h_u_arrmul24_and14_2;
  wire [0:0] h_u_arrmul24_fa14_2_xor1;
  wire [0:0] h_u_arrmul24_fa14_2_or0;
  wire [0:0] h_u_arrmul24_and15_2;
  wire [0:0] h_u_arrmul24_fa15_2_xor1;
  wire [0:0] h_u_arrmul24_fa15_2_or0;
  wire [0:0] h_u_arrmul24_and16_2;
  wire [0:0] h_u_arrmul24_fa16_2_xor1;
  wire [0:0] h_u_arrmul24_fa16_2_or0;
  wire [0:0] h_u_arrmul24_and17_2;
  wire [0:0] h_u_arrmul24_fa17_2_xor1;
  wire [0:0] h_u_arrmul24_fa17_2_or0;
  wire [0:0] h_u_arrmul24_and18_2;
  wire [0:0] h_u_arrmul24_fa18_2_xor1;
  wire [0:0] h_u_arrmul24_fa18_2_or0;
  wire [0:0] h_u_arrmul24_and19_2;
  wire [0:0] h_u_arrmul24_fa19_2_xor1;
  wire [0:0] h_u_arrmul24_fa19_2_or0;
  wire [0:0] h_u_arrmul24_and20_2;
  wire [0:0] h_u_arrmul24_fa20_2_xor1;
  wire [0:0] h_u_arrmul24_fa20_2_or0;
  wire [0:0] h_u_arrmul24_and21_2;
  wire [0:0] h_u_arrmul24_fa21_2_xor1;
  wire [0:0] h_u_arrmul24_fa21_2_or0;
  wire [0:0] h_u_arrmul24_and22_2;
  wire [0:0] h_u_arrmul24_fa22_2_xor1;
  wire [0:0] h_u_arrmul24_fa22_2_or0;
  wire [0:0] h_u_arrmul24_and23_2;
  wire [0:0] h_u_arrmul24_fa23_2_xor1;
  wire [0:0] h_u_arrmul24_fa23_2_or0;
  wire [0:0] h_u_arrmul24_and0_3;
  wire [0:0] h_u_arrmul24_ha0_3_xor0;
  wire [0:0] h_u_arrmul24_ha0_3_and0;
  wire [0:0] h_u_arrmul24_and1_3;
  wire [0:0] h_u_arrmul24_fa1_3_xor1;
  wire [0:0] h_u_arrmul24_fa1_3_or0;
  wire [0:0] h_u_arrmul24_and2_3;
  wire [0:0] h_u_arrmul24_fa2_3_xor1;
  wire [0:0] h_u_arrmul24_fa2_3_or0;
  wire [0:0] h_u_arrmul24_and3_3;
  wire [0:0] h_u_arrmul24_fa3_3_xor1;
  wire [0:0] h_u_arrmul24_fa3_3_or0;
  wire [0:0] h_u_arrmul24_and4_3;
  wire [0:0] h_u_arrmul24_fa4_3_xor1;
  wire [0:0] h_u_arrmul24_fa4_3_or0;
  wire [0:0] h_u_arrmul24_and5_3;
  wire [0:0] h_u_arrmul24_fa5_3_xor1;
  wire [0:0] h_u_arrmul24_fa5_3_or0;
  wire [0:0] h_u_arrmul24_and6_3;
  wire [0:0] h_u_arrmul24_fa6_3_xor1;
  wire [0:0] h_u_arrmul24_fa6_3_or0;
  wire [0:0] h_u_arrmul24_and7_3;
  wire [0:0] h_u_arrmul24_fa7_3_xor1;
  wire [0:0] h_u_arrmul24_fa7_3_or0;
  wire [0:0] h_u_arrmul24_and8_3;
  wire [0:0] h_u_arrmul24_fa8_3_xor1;
  wire [0:0] h_u_arrmul24_fa8_3_or0;
  wire [0:0] h_u_arrmul24_and9_3;
  wire [0:0] h_u_arrmul24_fa9_3_xor1;
  wire [0:0] h_u_arrmul24_fa9_3_or0;
  wire [0:0] h_u_arrmul24_and10_3;
  wire [0:0] h_u_arrmul24_fa10_3_xor1;
  wire [0:0] h_u_arrmul24_fa10_3_or0;
  wire [0:0] h_u_arrmul24_and11_3;
  wire [0:0] h_u_arrmul24_fa11_3_xor1;
  wire [0:0] h_u_arrmul24_fa11_3_or0;
  wire [0:0] h_u_arrmul24_and12_3;
  wire [0:0] h_u_arrmul24_fa12_3_xor1;
  wire [0:0] h_u_arrmul24_fa12_3_or0;
  wire [0:0] h_u_arrmul24_and13_3;
  wire [0:0] h_u_arrmul24_fa13_3_xor1;
  wire [0:0] h_u_arrmul24_fa13_3_or0;
  wire [0:0] h_u_arrmul24_and14_3;
  wire [0:0] h_u_arrmul24_fa14_3_xor1;
  wire [0:0] h_u_arrmul24_fa14_3_or0;
  wire [0:0] h_u_arrmul24_and15_3;
  wire [0:0] h_u_arrmul24_fa15_3_xor1;
  wire [0:0] h_u_arrmul24_fa15_3_or0;
  wire [0:0] h_u_arrmul24_and16_3;
  wire [0:0] h_u_arrmul24_fa16_3_xor1;
  wire [0:0] h_u_arrmul24_fa16_3_or0;
  wire [0:0] h_u_arrmul24_and17_3;
  wire [0:0] h_u_arrmul24_fa17_3_xor1;
  wire [0:0] h_u_arrmul24_fa17_3_or0;
  wire [0:0] h_u_arrmul24_and18_3;
  wire [0:0] h_u_arrmul24_fa18_3_xor1;
  wire [0:0] h_u_arrmul24_fa18_3_or0;
  wire [0:0] h_u_arrmul24_and19_3;
  wire [0:0] h_u_arrmul24_fa19_3_xor1;
  wire [0:0] h_u_arrmul24_fa19_3_or0;
  wire [0:0] h_u_arrmul24_and20_3;
  wire [0:0] h_u_arrmul24_fa20_3_xor1;
  wire [0:0] h_u_arrmul24_fa20_3_or0;
  wire [0:0] h_u_arrmul24_and21_3;
  wire [0:0] h_u_arrmul24_fa21_3_xor1;
  wire [0:0] h_u_arrmul24_fa21_3_or0;
  wire [0:0] h_u_arrmul24_and22_3;
  wire [0:0] h_u_arrmul24_fa22_3_xor1;
  wire [0:0] h_u_arrmul24_fa22_3_or0;
  wire [0:0] h_u_arrmul24_and23_3;
  wire [0:0] h_u_arrmul24_fa23_3_xor1;
  wire [0:0] h_u_arrmul24_fa23_3_or0;
  wire [0:0] h_u_arrmul24_and0_4;
  wire [0:0] h_u_arrmul24_ha0_4_xor0;
  wire [0:0] h_u_arrmul24_ha0_4_and0;
  wire [0:0] h_u_arrmul24_and1_4;
  wire [0:0] h_u_arrmul24_fa1_4_xor1;
  wire [0:0] h_u_arrmul24_fa1_4_or0;
  wire [0:0] h_u_arrmul24_and2_4;
  wire [0:0] h_u_arrmul24_fa2_4_xor1;
  wire [0:0] h_u_arrmul24_fa2_4_or0;
  wire [0:0] h_u_arrmul24_and3_4;
  wire [0:0] h_u_arrmul24_fa3_4_xor1;
  wire [0:0] h_u_arrmul24_fa3_4_or0;
  wire [0:0] h_u_arrmul24_and4_4;
  wire [0:0] h_u_arrmul24_fa4_4_xor1;
  wire [0:0] h_u_arrmul24_fa4_4_or0;
  wire [0:0] h_u_arrmul24_and5_4;
  wire [0:0] h_u_arrmul24_fa5_4_xor1;
  wire [0:0] h_u_arrmul24_fa5_4_or0;
  wire [0:0] h_u_arrmul24_and6_4;
  wire [0:0] h_u_arrmul24_fa6_4_xor1;
  wire [0:0] h_u_arrmul24_fa6_4_or0;
  wire [0:0] h_u_arrmul24_and7_4;
  wire [0:0] h_u_arrmul24_fa7_4_xor1;
  wire [0:0] h_u_arrmul24_fa7_4_or0;
  wire [0:0] h_u_arrmul24_and8_4;
  wire [0:0] h_u_arrmul24_fa8_4_xor1;
  wire [0:0] h_u_arrmul24_fa8_4_or0;
  wire [0:0] h_u_arrmul24_and9_4;
  wire [0:0] h_u_arrmul24_fa9_4_xor1;
  wire [0:0] h_u_arrmul24_fa9_4_or0;
  wire [0:0] h_u_arrmul24_and10_4;
  wire [0:0] h_u_arrmul24_fa10_4_xor1;
  wire [0:0] h_u_arrmul24_fa10_4_or0;
  wire [0:0] h_u_arrmul24_and11_4;
  wire [0:0] h_u_arrmul24_fa11_4_xor1;
  wire [0:0] h_u_arrmul24_fa11_4_or0;
  wire [0:0] h_u_arrmul24_and12_4;
  wire [0:0] h_u_arrmul24_fa12_4_xor1;
  wire [0:0] h_u_arrmul24_fa12_4_or0;
  wire [0:0] h_u_arrmul24_and13_4;
  wire [0:0] h_u_arrmul24_fa13_4_xor1;
  wire [0:0] h_u_arrmul24_fa13_4_or0;
  wire [0:0] h_u_arrmul24_and14_4;
  wire [0:0] h_u_arrmul24_fa14_4_xor1;
  wire [0:0] h_u_arrmul24_fa14_4_or0;
  wire [0:0] h_u_arrmul24_and15_4;
  wire [0:0] h_u_arrmul24_fa15_4_xor1;
  wire [0:0] h_u_arrmul24_fa15_4_or0;
  wire [0:0] h_u_arrmul24_and16_4;
  wire [0:0] h_u_arrmul24_fa16_4_xor1;
  wire [0:0] h_u_arrmul24_fa16_4_or0;
  wire [0:0] h_u_arrmul24_and17_4;
  wire [0:0] h_u_arrmul24_fa17_4_xor1;
  wire [0:0] h_u_arrmul24_fa17_4_or0;
  wire [0:0] h_u_arrmul24_and18_4;
  wire [0:0] h_u_arrmul24_fa18_4_xor1;
  wire [0:0] h_u_arrmul24_fa18_4_or0;
  wire [0:0] h_u_arrmul24_and19_4;
  wire [0:0] h_u_arrmul24_fa19_4_xor1;
  wire [0:0] h_u_arrmul24_fa19_4_or0;
  wire [0:0] h_u_arrmul24_and20_4;
  wire [0:0] h_u_arrmul24_fa20_4_xor1;
  wire [0:0] h_u_arrmul24_fa20_4_or0;
  wire [0:0] h_u_arrmul24_and21_4;
  wire [0:0] h_u_arrmul24_fa21_4_xor1;
  wire [0:0] h_u_arrmul24_fa21_4_or0;
  wire [0:0] h_u_arrmul24_and22_4;
  wire [0:0] h_u_arrmul24_fa22_4_xor1;
  wire [0:0] h_u_arrmul24_fa22_4_or0;
  wire [0:0] h_u_arrmul24_and23_4;
  wire [0:0] h_u_arrmul24_fa23_4_xor1;
  wire [0:0] h_u_arrmul24_fa23_4_or0;
  wire [0:0] h_u_arrmul24_and0_5;
  wire [0:0] h_u_arrmul24_ha0_5_xor0;
  wire [0:0] h_u_arrmul24_ha0_5_and0;
  wire [0:0] h_u_arrmul24_and1_5;
  wire [0:0] h_u_arrmul24_fa1_5_xor1;
  wire [0:0] h_u_arrmul24_fa1_5_or0;
  wire [0:0] h_u_arrmul24_and2_5;
  wire [0:0] h_u_arrmul24_fa2_5_xor1;
  wire [0:0] h_u_arrmul24_fa2_5_or0;
  wire [0:0] h_u_arrmul24_and3_5;
  wire [0:0] h_u_arrmul24_fa3_5_xor1;
  wire [0:0] h_u_arrmul24_fa3_5_or0;
  wire [0:0] h_u_arrmul24_and4_5;
  wire [0:0] h_u_arrmul24_fa4_5_xor1;
  wire [0:0] h_u_arrmul24_fa4_5_or0;
  wire [0:0] h_u_arrmul24_and5_5;
  wire [0:0] h_u_arrmul24_fa5_5_xor1;
  wire [0:0] h_u_arrmul24_fa5_5_or0;
  wire [0:0] h_u_arrmul24_and6_5;
  wire [0:0] h_u_arrmul24_fa6_5_xor1;
  wire [0:0] h_u_arrmul24_fa6_5_or0;
  wire [0:0] h_u_arrmul24_and7_5;
  wire [0:0] h_u_arrmul24_fa7_5_xor1;
  wire [0:0] h_u_arrmul24_fa7_5_or0;
  wire [0:0] h_u_arrmul24_and8_5;
  wire [0:0] h_u_arrmul24_fa8_5_xor1;
  wire [0:0] h_u_arrmul24_fa8_5_or0;
  wire [0:0] h_u_arrmul24_and9_5;
  wire [0:0] h_u_arrmul24_fa9_5_xor1;
  wire [0:0] h_u_arrmul24_fa9_5_or0;
  wire [0:0] h_u_arrmul24_and10_5;
  wire [0:0] h_u_arrmul24_fa10_5_xor1;
  wire [0:0] h_u_arrmul24_fa10_5_or0;
  wire [0:0] h_u_arrmul24_and11_5;
  wire [0:0] h_u_arrmul24_fa11_5_xor1;
  wire [0:0] h_u_arrmul24_fa11_5_or0;
  wire [0:0] h_u_arrmul24_and12_5;
  wire [0:0] h_u_arrmul24_fa12_5_xor1;
  wire [0:0] h_u_arrmul24_fa12_5_or0;
  wire [0:0] h_u_arrmul24_and13_5;
  wire [0:0] h_u_arrmul24_fa13_5_xor1;
  wire [0:0] h_u_arrmul24_fa13_5_or0;
  wire [0:0] h_u_arrmul24_and14_5;
  wire [0:0] h_u_arrmul24_fa14_5_xor1;
  wire [0:0] h_u_arrmul24_fa14_5_or0;
  wire [0:0] h_u_arrmul24_and15_5;
  wire [0:0] h_u_arrmul24_fa15_5_xor1;
  wire [0:0] h_u_arrmul24_fa15_5_or0;
  wire [0:0] h_u_arrmul24_and16_5;
  wire [0:0] h_u_arrmul24_fa16_5_xor1;
  wire [0:0] h_u_arrmul24_fa16_5_or0;
  wire [0:0] h_u_arrmul24_and17_5;
  wire [0:0] h_u_arrmul24_fa17_5_xor1;
  wire [0:0] h_u_arrmul24_fa17_5_or0;
  wire [0:0] h_u_arrmul24_and18_5;
  wire [0:0] h_u_arrmul24_fa18_5_xor1;
  wire [0:0] h_u_arrmul24_fa18_5_or0;
  wire [0:0] h_u_arrmul24_and19_5;
  wire [0:0] h_u_arrmul24_fa19_5_xor1;
  wire [0:0] h_u_arrmul24_fa19_5_or0;
  wire [0:0] h_u_arrmul24_and20_5;
  wire [0:0] h_u_arrmul24_fa20_5_xor1;
  wire [0:0] h_u_arrmul24_fa20_5_or0;
  wire [0:0] h_u_arrmul24_and21_5;
  wire [0:0] h_u_arrmul24_fa21_5_xor1;
  wire [0:0] h_u_arrmul24_fa21_5_or0;
  wire [0:0] h_u_arrmul24_and22_5;
  wire [0:0] h_u_arrmul24_fa22_5_xor1;
  wire [0:0] h_u_arrmul24_fa22_5_or0;
  wire [0:0] h_u_arrmul24_and23_5;
  wire [0:0] h_u_arrmul24_fa23_5_xor1;
  wire [0:0] h_u_arrmul24_fa23_5_or0;
  wire [0:0] h_u_arrmul24_and0_6;
  wire [0:0] h_u_arrmul24_ha0_6_xor0;
  wire [0:0] h_u_arrmul24_ha0_6_and0;
  wire [0:0] h_u_arrmul24_and1_6;
  wire [0:0] h_u_arrmul24_fa1_6_xor1;
  wire [0:0] h_u_arrmul24_fa1_6_or0;
  wire [0:0] h_u_arrmul24_and2_6;
  wire [0:0] h_u_arrmul24_fa2_6_xor1;
  wire [0:0] h_u_arrmul24_fa2_6_or0;
  wire [0:0] h_u_arrmul24_and3_6;
  wire [0:0] h_u_arrmul24_fa3_6_xor1;
  wire [0:0] h_u_arrmul24_fa3_6_or0;
  wire [0:0] h_u_arrmul24_and4_6;
  wire [0:0] h_u_arrmul24_fa4_6_xor1;
  wire [0:0] h_u_arrmul24_fa4_6_or0;
  wire [0:0] h_u_arrmul24_and5_6;
  wire [0:0] h_u_arrmul24_fa5_6_xor1;
  wire [0:0] h_u_arrmul24_fa5_6_or0;
  wire [0:0] h_u_arrmul24_and6_6;
  wire [0:0] h_u_arrmul24_fa6_6_xor1;
  wire [0:0] h_u_arrmul24_fa6_6_or0;
  wire [0:0] h_u_arrmul24_and7_6;
  wire [0:0] h_u_arrmul24_fa7_6_xor1;
  wire [0:0] h_u_arrmul24_fa7_6_or0;
  wire [0:0] h_u_arrmul24_and8_6;
  wire [0:0] h_u_arrmul24_fa8_6_xor1;
  wire [0:0] h_u_arrmul24_fa8_6_or0;
  wire [0:0] h_u_arrmul24_and9_6;
  wire [0:0] h_u_arrmul24_fa9_6_xor1;
  wire [0:0] h_u_arrmul24_fa9_6_or0;
  wire [0:0] h_u_arrmul24_and10_6;
  wire [0:0] h_u_arrmul24_fa10_6_xor1;
  wire [0:0] h_u_arrmul24_fa10_6_or0;
  wire [0:0] h_u_arrmul24_and11_6;
  wire [0:0] h_u_arrmul24_fa11_6_xor1;
  wire [0:0] h_u_arrmul24_fa11_6_or0;
  wire [0:0] h_u_arrmul24_and12_6;
  wire [0:0] h_u_arrmul24_fa12_6_xor1;
  wire [0:0] h_u_arrmul24_fa12_6_or0;
  wire [0:0] h_u_arrmul24_and13_6;
  wire [0:0] h_u_arrmul24_fa13_6_xor1;
  wire [0:0] h_u_arrmul24_fa13_6_or0;
  wire [0:0] h_u_arrmul24_and14_6;
  wire [0:0] h_u_arrmul24_fa14_6_xor1;
  wire [0:0] h_u_arrmul24_fa14_6_or0;
  wire [0:0] h_u_arrmul24_and15_6;
  wire [0:0] h_u_arrmul24_fa15_6_xor1;
  wire [0:0] h_u_arrmul24_fa15_6_or0;
  wire [0:0] h_u_arrmul24_and16_6;
  wire [0:0] h_u_arrmul24_fa16_6_xor1;
  wire [0:0] h_u_arrmul24_fa16_6_or0;
  wire [0:0] h_u_arrmul24_and17_6;
  wire [0:0] h_u_arrmul24_fa17_6_xor1;
  wire [0:0] h_u_arrmul24_fa17_6_or0;
  wire [0:0] h_u_arrmul24_and18_6;
  wire [0:0] h_u_arrmul24_fa18_6_xor1;
  wire [0:0] h_u_arrmul24_fa18_6_or0;
  wire [0:0] h_u_arrmul24_and19_6;
  wire [0:0] h_u_arrmul24_fa19_6_xor1;
  wire [0:0] h_u_arrmul24_fa19_6_or0;
  wire [0:0] h_u_arrmul24_and20_6;
  wire [0:0] h_u_arrmul24_fa20_6_xor1;
  wire [0:0] h_u_arrmul24_fa20_6_or0;
  wire [0:0] h_u_arrmul24_and21_6;
  wire [0:0] h_u_arrmul24_fa21_6_xor1;
  wire [0:0] h_u_arrmul24_fa21_6_or0;
  wire [0:0] h_u_arrmul24_and22_6;
  wire [0:0] h_u_arrmul24_fa22_6_xor1;
  wire [0:0] h_u_arrmul24_fa22_6_or0;
  wire [0:0] h_u_arrmul24_and23_6;
  wire [0:0] h_u_arrmul24_fa23_6_xor1;
  wire [0:0] h_u_arrmul24_fa23_6_or0;
  wire [0:0] h_u_arrmul24_and0_7;
  wire [0:0] h_u_arrmul24_ha0_7_xor0;
  wire [0:0] h_u_arrmul24_ha0_7_and0;
  wire [0:0] h_u_arrmul24_and1_7;
  wire [0:0] h_u_arrmul24_fa1_7_xor1;
  wire [0:0] h_u_arrmul24_fa1_7_or0;
  wire [0:0] h_u_arrmul24_and2_7;
  wire [0:0] h_u_arrmul24_fa2_7_xor1;
  wire [0:0] h_u_arrmul24_fa2_7_or0;
  wire [0:0] h_u_arrmul24_and3_7;
  wire [0:0] h_u_arrmul24_fa3_7_xor1;
  wire [0:0] h_u_arrmul24_fa3_7_or0;
  wire [0:0] h_u_arrmul24_and4_7;
  wire [0:0] h_u_arrmul24_fa4_7_xor1;
  wire [0:0] h_u_arrmul24_fa4_7_or0;
  wire [0:0] h_u_arrmul24_and5_7;
  wire [0:0] h_u_arrmul24_fa5_7_xor1;
  wire [0:0] h_u_arrmul24_fa5_7_or0;
  wire [0:0] h_u_arrmul24_and6_7;
  wire [0:0] h_u_arrmul24_fa6_7_xor1;
  wire [0:0] h_u_arrmul24_fa6_7_or0;
  wire [0:0] h_u_arrmul24_and7_7;
  wire [0:0] h_u_arrmul24_fa7_7_xor1;
  wire [0:0] h_u_arrmul24_fa7_7_or0;
  wire [0:0] h_u_arrmul24_and8_7;
  wire [0:0] h_u_arrmul24_fa8_7_xor1;
  wire [0:0] h_u_arrmul24_fa8_7_or0;
  wire [0:0] h_u_arrmul24_and9_7;
  wire [0:0] h_u_arrmul24_fa9_7_xor1;
  wire [0:0] h_u_arrmul24_fa9_7_or0;
  wire [0:0] h_u_arrmul24_and10_7;
  wire [0:0] h_u_arrmul24_fa10_7_xor1;
  wire [0:0] h_u_arrmul24_fa10_7_or0;
  wire [0:0] h_u_arrmul24_and11_7;
  wire [0:0] h_u_arrmul24_fa11_7_xor1;
  wire [0:0] h_u_arrmul24_fa11_7_or0;
  wire [0:0] h_u_arrmul24_and12_7;
  wire [0:0] h_u_arrmul24_fa12_7_xor1;
  wire [0:0] h_u_arrmul24_fa12_7_or0;
  wire [0:0] h_u_arrmul24_and13_7;
  wire [0:0] h_u_arrmul24_fa13_7_xor1;
  wire [0:0] h_u_arrmul24_fa13_7_or0;
  wire [0:0] h_u_arrmul24_and14_7;
  wire [0:0] h_u_arrmul24_fa14_7_xor1;
  wire [0:0] h_u_arrmul24_fa14_7_or0;
  wire [0:0] h_u_arrmul24_and15_7;
  wire [0:0] h_u_arrmul24_fa15_7_xor1;
  wire [0:0] h_u_arrmul24_fa15_7_or0;
  wire [0:0] h_u_arrmul24_and16_7;
  wire [0:0] h_u_arrmul24_fa16_7_xor1;
  wire [0:0] h_u_arrmul24_fa16_7_or0;
  wire [0:0] h_u_arrmul24_and17_7;
  wire [0:0] h_u_arrmul24_fa17_7_xor1;
  wire [0:0] h_u_arrmul24_fa17_7_or0;
  wire [0:0] h_u_arrmul24_and18_7;
  wire [0:0] h_u_arrmul24_fa18_7_xor1;
  wire [0:0] h_u_arrmul24_fa18_7_or0;
  wire [0:0] h_u_arrmul24_and19_7;
  wire [0:0] h_u_arrmul24_fa19_7_xor1;
  wire [0:0] h_u_arrmul24_fa19_7_or0;
  wire [0:0] h_u_arrmul24_and20_7;
  wire [0:0] h_u_arrmul24_fa20_7_xor1;
  wire [0:0] h_u_arrmul24_fa20_7_or0;
  wire [0:0] h_u_arrmul24_and21_7;
  wire [0:0] h_u_arrmul24_fa21_7_xor1;
  wire [0:0] h_u_arrmul24_fa21_7_or0;
  wire [0:0] h_u_arrmul24_and22_7;
  wire [0:0] h_u_arrmul24_fa22_7_xor1;
  wire [0:0] h_u_arrmul24_fa22_7_or0;
  wire [0:0] h_u_arrmul24_and23_7;
  wire [0:0] h_u_arrmul24_fa23_7_xor1;
  wire [0:0] h_u_arrmul24_fa23_7_or0;
  wire [0:0] h_u_arrmul24_and0_8;
  wire [0:0] h_u_arrmul24_ha0_8_xor0;
  wire [0:0] h_u_arrmul24_ha0_8_and0;
  wire [0:0] h_u_arrmul24_and1_8;
  wire [0:0] h_u_arrmul24_fa1_8_xor1;
  wire [0:0] h_u_arrmul24_fa1_8_or0;
  wire [0:0] h_u_arrmul24_and2_8;
  wire [0:0] h_u_arrmul24_fa2_8_xor1;
  wire [0:0] h_u_arrmul24_fa2_8_or0;
  wire [0:0] h_u_arrmul24_and3_8;
  wire [0:0] h_u_arrmul24_fa3_8_xor1;
  wire [0:0] h_u_arrmul24_fa3_8_or0;
  wire [0:0] h_u_arrmul24_and4_8;
  wire [0:0] h_u_arrmul24_fa4_8_xor1;
  wire [0:0] h_u_arrmul24_fa4_8_or0;
  wire [0:0] h_u_arrmul24_and5_8;
  wire [0:0] h_u_arrmul24_fa5_8_xor1;
  wire [0:0] h_u_arrmul24_fa5_8_or0;
  wire [0:0] h_u_arrmul24_and6_8;
  wire [0:0] h_u_arrmul24_fa6_8_xor1;
  wire [0:0] h_u_arrmul24_fa6_8_or0;
  wire [0:0] h_u_arrmul24_and7_8;
  wire [0:0] h_u_arrmul24_fa7_8_xor1;
  wire [0:0] h_u_arrmul24_fa7_8_or0;
  wire [0:0] h_u_arrmul24_and8_8;
  wire [0:0] h_u_arrmul24_fa8_8_xor1;
  wire [0:0] h_u_arrmul24_fa8_8_or0;
  wire [0:0] h_u_arrmul24_and9_8;
  wire [0:0] h_u_arrmul24_fa9_8_xor1;
  wire [0:0] h_u_arrmul24_fa9_8_or0;
  wire [0:0] h_u_arrmul24_and10_8;
  wire [0:0] h_u_arrmul24_fa10_8_xor1;
  wire [0:0] h_u_arrmul24_fa10_8_or0;
  wire [0:0] h_u_arrmul24_and11_8;
  wire [0:0] h_u_arrmul24_fa11_8_xor1;
  wire [0:0] h_u_arrmul24_fa11_8_or0;
  wire [0:0] h_u_arrmul24_and12_8;
  wire [0:0] h_u_arrmul24_fa12_8_xor1;
  wire [0:0] h_u_arrmul24_fa12_8_or0;
  wire [0:0] h_u_arrmul24_and13_8;
  wire [0:0] h_u_arrmul24_fa13_8_xor1;
  wire [0:0] h_u_arrmul24_fa13_8_or0;
  wire [0:0] h_u_arrmul24_and14_8;
  wire [0:0] h_u_arrmul24_fa14_8_xor1;
  wire [0:0] h_u_arrmul24_fa14_8_or0;
  wire [0:0] h_u_arrmul24_and15_8;
  wire [0:0] h_u_arrmul24_fa15_8_xor1;
  wire [0:0] h_u_arrmul24_fa15_8_or0;
  wire [0:0] h_u_arrmul24_and16_8;
  wire [0:0] h_u_arrmul24_fa16_8_xor1;
  wire [0:0] h_u_arrmul24_fa16_8_or0;
  wire [0:0] h_u_arrmul24_and17_8;
  wire [0:0] h_u_arrmul24_fa17_8_xor1;
  wire [0:0] h_u_arrmul24_fa17_8_or0;
  wire [0:0] h_u_arrmul24_and18_8;
  wire [0:0] h_u_arrmul24_fa18_8_xor1;
  wire [0:0] h_u_arrmul24_fa18_8_or0;
  wire [0:0] h_u_arrmul24_and19_8;
  wire [0:0] h_u_arrmul24_fa19_8_xor1;
  wire [0:0] h_u_arrmul24_fa19_8_or0;
  wire [0:0] h_u_arrmul24_and20_8;
  wire [0:0] h_u_arrmul24_fa20_8_xor1;
  wire [0:0] h_u_arrmul24_fa20_8_or0;
  wire [0:0] h_u_arrmul24_and21_8;
  wire [0:0] h_u_arrmul24_fa21_8_xor1;
  wire [0:0] h_u_arrmul24_fa21_8_or0;
  wire [0:0] h_u_arrmul24_and22_8;
  wire [0:0] h_u_arrmul24_fa22_8_xor1;
  wire [0:0] h_u_arrmul24_fa22_8_or0;
  wire [0:0] h_u_arrmul24_and23_8;
  wire [0:0] h_u_arrmul24_fa23_8_xor1;
  wire [0:0] h_u_arrmul24_fa23_8_or0;
  wire [0:0] h_u_arrmul24_and0_9;
  wire [0:0] h_u_arrmul24_ha0_9_xor0;
  wire [0:0] h_u_arrmul24_ha0_9_and0;
  wire [0:0] h_u_arrmul24_and1_9;
  wire [0:0] h_u_arrmul24_fa1_9_xor1;
  wire [0:0] h_u_arrmul24_fa1_9_or0;
  wire [0:0] h_u_arrmul24_and2_9;
  wire [0:0] h_u_arrmul24_fa2_9_xor1;
  wire [0:0] h_u_arrmul24_fa2_9_or0;
  wire [0:0] h_u_arrmul24_and3_9;
  wire [0:0] h_u_arrmul24_fa3_9_xor1;
  wire [0:0] h_u_arrmul24_fa3_9_or0;
  wire [0:0] h_u_arrmul24_and4_9;
  wire [0:0] h_u_arrmul24_fa4_9_xor1;
  wire [0:0] h_u_arrmul24_fa4_9_or0;
  wire [0:0] h_u_arrmul24_and5_9;
  wire [0:0] h_u_arrmul24_fa5_9_xor1;
  wire [0:0] h_u_arrmul24_fa5_9_or0;
  wire [0:0] h_u_arrmul24_and6_9;
  wire [0:0] h_u_arrmul24_fa6_9_xor1;
  wire [0:0] h_u_arrmul24_fa6_9_or0;
  wire [0:0] h_u_arrmul24_and7_9;
  wire [0:0] h_u_arrmul24_fa7_9_xor1;
  wire [0:0] h_u_arrmul24_fa7_9_or0;
  wire [0:0] h_u_arrmul24_and8_9;
  wire [0:0] h_u_arrmul24_fa8_9_xor1;
  wire [0:0] h_u_arrmul24_fa8_9_or0;
  wire [0:0] h_u_arrmul24_and9_9;
  wire [0:0] h_u_arrmul24_fa9_9_xor1;
  wire [0:0] h_u_arrmul24_fa9_9_or0;
  wire [0:0] h_u_arrmul24_and10_9;
  wire [0:0] h_u_arrmul24_fa10_9_xor1;
  wire [0:0] h_u_arrmul24_fa10_9_or0;
  wire [0:0] h_u_arrmul24_and11_9;
  wire [0:0] h_u_arrmul24_fa11_9_xor1;
  wire [0:0] h_u_arrmul24_fa11_9_or0;
  wire [0:0] h_u_arrmul24_and12_9;
  wire [0:0] h_u_arrmul24_fa12_9_xor1;
  wire [0:0] h_u_arrmul24_fa12_9_or0;
  wire [0:0] h_u_arrmul24_and13_9;
  wire [0:0] h_u_arrmul24_fa13_9_xor1;
  wire [0:0] h_u_arrmul24_fa13_9_or0;
  wire [0:0] h_u_arrmul24_and14_9;
  wire [0:0] h_u_arrmul24_fa14_9_xor1;
  wire [0:0] h_u_arrmul24_fa14_9_or0;
  wire [0:0] h_u_arrmul24_and15_9;
  wire [0:0] h_u_arrmul24_fa15_9_xor1;
  wire [0:0] h_u_arrmul24_fa15_9_or0;
  wire [0:0] h_u_arrmul24_and16_9;
  wire [0:0] h_u_arrmul24_fa16_9_xor1;
  wire [0:0] h_u_arrmul24_fa16_9_or0;
  wire [0:0] h_u_arrmul24_and17_9;
  wire [0:0] h_u_arrmul24_fa17_9_xor1;
  wire [0:0] h_u_arrmul24_fa17_9_or0;
  wire [0:0] h_u_arrmul24_and18_9;
  wire [0:0] h_u_arrmul24_fa18_9_xor1;
  wire [0:0] h_u_arrmul24_fa18_9_or0;
  wire [0:0] h_u_arrmul24_and19_9;
  wire [0:0] h_u_arrmul24_fa19_9_xor1;
  wire [0:0] h_u_arrmul24_fa19_9_or0;
  wire [0:0] h_u_arrmul24_and20_9;
  wire [0:0] h_u_arrmul24_fa20_9_xor1;
  wire [0:0] h_u_arrmul24_fa20_9_or0;
  wire [0:0] h_u_arrmul24_and21_9;
  wire [0:0] h_u_arrmul24_fa21_9_xor1;
  wire [0:0] h_u_arrmul24_fa21_9_or0;
  wire [0:0] h_u_arrmul24_and22_9;
  wire [0:0] h_u_arrmul24_fa22_9_xor1;
  wire [0:0] h_u_arrmul24_fa22_9_or0;
  wire [0:0] h_u_arrmul24_and23_9;
  wire [0:0] h_u_arrmul24_fa23_9_xor1;
  wire [0:0] h_u_arrmul24_fa23_9_or0;
  wire [0:0] h_u_arrmul24_and0_10;
  wire [0:0] h_u_arrmul24_ha0_10_xor0;
  wire [0:0] h_u_arrmul24_ha0_10_and0;
  wire [0:0] h_u_arrmul24_and1_10;
  wire [0:0] h_u_arrmul24_fa1_10_xor1;
  wire [0:0] h_u_arrmul24_fa1_10_or0;
  wire [0:0] h_u_arrmul24_and2_10;
  wire [0:0] h_u_arrmul24_fa2_10_xor1;
  wire [0:0] h_u_arrmul24_fa2_10_or0;
  wire [0:0] h_u_arrmul24_and3_10;
  wire [0:0] h_u_arrmul24_fa3_10_xor1;
  wire [0:0] h_u_arrmul24_fa3_10_or0;
  wire [0:0] h_u_arrmul24_and4_10;
  wire [0:0] h_u_arrmul24_fa4_10_xor1;
  wire [0:0] h_u_arrmul24_fa4_10_or0;
  wire [0:0] h_u_arrmul24_and5_10;
  wire [0:0] h_u_arrmul24_fa5_10_xor1;
  wire [0:0] h_u_arrmul24_fa5_10_or0;
  wire [0:0] h_u_arrmul24_and6_10;
  wire [0:0] h_u_arrmul24_fa6_10_xor1;
  wire [0:0] h_u_arrmul24_fa6_10_or0;
  wire [0:0] h_u_arrmul24_and7_10;
  wire [0:0] h_u_arrmul24_fa7_10_xor1;
  wire [0:0] h_u_arrmul24_fa7_10_or0;
  wire [0:0] h_u_arrmul24_and8_10;
  wire [0:0] h_u_arrmul24_fa8_10_xor1;
  wire [0:0] h_u_arrmul24_fa8_10_or0;
  wire [0:0] h_u_arrmul24_and9_10;
  wire [0:0] h_u_arrmul24_fa9_10_xor1;
  wire [0:0] h_u_arrmul24_fa9_10_or0;
  wire [0:0] h_u_arrmul24_and10_10;
  wire [0:0] h_u_arrmul24_fa10_10_xor1;
  wire [0:0] h_u_arrmul24_fa10_10_or0;
  wire [0:0] h_u_arrmul24_and11_10;
  wire [0:0] h_u_arrmul24_fa11_10_xor1;
  wire [0:0] h_u_arrmul24_fa11_10_or0;
  wire [0:0] h_u_arrmul24_and12_10;
  wire [0:0] h_u_arrmul24_fa12_10_xor1;
  wire [0:0] h_u_arrmul24_fa12_10_or0;
  wire [0:0] h_u_arrmul24_and13_10;
  wire [0:0] h_u_arrmul24_fa13_10_xor1;
  wire [0:0] h_u_arrmul24_fa13_10_or0;
  wire [0:0] h_u_arrmul24_and14_10;
  wire [0:0] h_u_arrmul24_fa14_10_xor1;
  wire [0:0] h_u_arrmul24_fa14_10_or0;
  wire [0:0] h_u_arrmul24_and15_10;
  wire [0:0] h_u_arrmul24_fa15_10_xor1;
  wire [0:0] h_u_arrmul24_fa15_10_or0;
  wire [0:0] h_u_arrmul24_and16_10;
  wire [0:0] h_u_arrmul24_fa16_10_xor1;
  wire [0:0] h_u_arrmul24_fa16_10_or0;
  wire [0:0] h_u_arrmul24_and17_10;
  wire [0:0] h_u_arrmul24_fa17_10_xor1;
  wire [0:0] h_u_arrmul24_fa17_10_or0;
  wire [0:0] h_u_arrmul24_and18_10;
  wire [0:0] h_u_arrmul24_fa18_10_xor1;
  wire [0:0] h_u_arrmul24_fa18_10_or0;
  wire [0:0] h_u_arrmul24_and19_10;
  wire [0:0] h_u_arrmul24_fa19_10_xor1;
  wire [0:0] h_u_arrmul24_fa19_10_or0;
  wire [0:0] h_u_arrmul24_and20_10;
  wire [0:0] h_u_arrmul24_fa20_10_xor1;
  wire [0:0] h_u_arrmul24_fa20_10_or0;
  wire [0:0] h_u_arrmul24_and21_10;
  wire [0:0] h_u_arrmul24_fa21_10_xor1;
  wire [0:0] h_u_arrmul24_fa21_10_or0;
  wire [0:0] h_u_arrmul24_and22_10;
  wire [0:0] h_u_arrmul24_fa22_10_xor1;
  wire [0:0] h_u_arrmul24_fa22_10_or0;
  wire [0:0] h_u_arrmul24_and23_10;
  wire [0:0] h_u_arrmul24_fa23_10_xor1;
  wire [0:0] h_u_arrmul24_fa23_10_or0;
  wire [0:0] h_u_arrmul24_and0_11;
  wire [0:0] h_u_arrmul24_ha0_11_xor0;
  wire [0:0] h_u_arrmul24_ha0_11_and0;
  wire [0:0] h_u_arrmul24_and1_11;
  wire [0:0] h_u_arrmul24_fa1_11_xor1;
  wire [0:0] h_u_arrmul24_fa1_11_or0;
  wire [0:0] h_u_arrmul24_and2_11;
  wire [0:0] h_u_arrmul24_fa2_11_xor1;
  wire [0:0] h_u_arrmul24_fa2_11_or0;
  wire [0:0] h_u_arrmul24_and3_11;
  wire [0:0] h_u_arrmul24_fa3_11_xor1;
  wire [0:0] h_u_arrmul24_fa3_11_or0;
  wire [0:0] h_u_arrmul24_and4_11;
  wire [0:0] h_u_arrmul24_fa4_11_xor1;
  wire [0:0] h_u_arrmul24_fa4_11_or0;
  wire [0:0] h_u_arrmul24_and5_11;
  wire [0:0] h_u_arrmul24_fa5_11_xor1;
  wire [0:0] h_u_arrmul24_fa5_11_or0;
  wire [0:0] h_u_arrmul24_and6_11;
  wire [0:0] h_u_arrmul24_fa6_11_xor1;
  wire [0:0] h_u_arrmul24_fa6_11_or0;
  wire [0:0] h_u_arrmul24_and7_11;
  wire [0:0] h_u_arrmul24_fa7_11_xor1;
  wire [0:0] h_u_arrmul24_fa7_11_or0;
  wire [0:0] h_u_arrmul24_and8_11;
  wire [0:0] h_u_arrmul24_fa8_11_xor1;
  wire [0:0] h_u_arrmul24_fa8_11_or0;
  wire [0:0] h_u_arrmul24_and9_11;
  wire [0:0] h_u_arrmul24_fa9_11_xor1;
  wire [0:0] h_u_arrmul24_fa9_11_or0;
  wire [0:0] h_u_arrmul24_and10_11;
  wire [0:0] h_u_arrmul24_fa10_11_xor1;
  wire [0:0] h_u_arrmul24_fa10_11_or0;
  wire [0:0] h_u_arrmul24_and11_11;
  wire [0:0] h_u_arrmul24_fa11_11_xor1;
  wire [0:0] h_u_arrmul24_fa11_11_or0;
  wire [0:0] h_u_arrmul24_and12_11;
  wire [0:0] h_u_arrmul24_fa12_11_xor1;
  wire [0:0] h_u_arrmul24_fa12_11_or0;
  wire [0:0] h_u_arrmul24_and13_11;
  wire [0:0] h_u_arrmul24_fa13_11_xor1;
  wire [0:0] h_u_arrmul24_fa13_11_or0;
  wire [0:0] h_u_arrmul24_and14_11;
  wire [0:0] h_u_arrmul24_fa14_11_xor1;
  wire [0:0] h_u_arrmul24_fa14_11_or0;
  wire [0:0] h_u_arrmul24_and15_11;
  wire [0:0] h_u_arrmul24_fa15_11_xor1;
  wire [0:0] h_u_arrmul24_fa15_11_or0;
  wire [0:0] h_u_arrmul24_and16_11;
  wire [0:0] h_u_arrmul24_fa16_11_xor1;
  wire [0:0] h_u_arrmul24_fa16_11_or0;
  wire [0:0] h_u_arrmul24_and17_11;
  wire [0:0] h_u_arrmul24_fa17_11_xor1;
  wire [0:0] h_u_arrmul24_fa17_11_or0;
  wire [0:0] h_u_arrmul24_and18_11;
  wire [0:0] h_u_arrmul24_fa18_11_xor1;
  wire [0:0] h_u_arrmul24_fa18_11_or0;
  wire [0:0] h_u_arrmul24_and19_11;
  wire [0:0] h_u_arrmul24_fa19_11_xor1;
  wire [0:0] h_u_arrmul24_fa19_11_or0;
  wire [0:0] h_u_arrmul24_and20_11;
  wire [0:0] h_u_arrmul24_fa20_11_xor1;
  wire [0:0] h_u_arrmul24_fa20_11_or0;
  wire [0:0] h_u_arrmul24_and21_11;
  wire [0:0] h_u_arrmul24_fa21_11_xor1;
  wire [0:0] h_u_arrmul24_fa21_11_or0;
  wire [0:0] h_u_arrmul24_and22_11;
  wire [0:0] h_u_arrmul24_fa22_11_xor1;
  wire [0:0] h_u_arrmul24_fa22_11_or0;
  wire [0:0] h_u_arrmul24_and23_11;
  wire [0:0] h_u_arrmul24_fa23_11_xor1;
  wire [0:0] h_u_arrmul24_fa23_11_or0;
  wire [0:0] h_u_arrmul24_and0_12;
  wire [0:0] h_u_arrmul24_ha0_12_xor0;
  wire [0:0] h_u_arrmul24_ha0_12_and0;
  wire [0:0] h_u_arrmul24_and1_12;
  wire [0:0] h_u_arrmul24_fa1_12_xor1;
  wire [0:0] h_u_arrmul24_fa1_12_or0;
  wire [0:0] h_u_arrmul24_and2_12;
  wire [0:0] h_u_arrmul24_fa2_12_xor1;
  wire [0:0] h_u_arrmul24_fa2_12_or0;
  wire [0:0] h_u_arrmul24_and3_12;
  wire [0:0] h_u_arrmul24_fa3_12_xor1;
  wire [0:0] h_u_arrmul24_fa3_12_or0;
  wire [0:0] h_u_arrmul24_and4_12;
  wire [0:0] h_u_arrmul24_fa4_12_xor1;
  wire [0:0] h_u_arrmul24_fa4_12_or0;
  wire [0:0] h_u_arrmul24_and5_12;
  wire [0:0] h_u_arrmul24_fa5_12_xor1;
  wire [0:0] h_u_arrmul24_fa5_12_or0;
  wire [0:0] h_u_arrmul24_and6_12;
  wire [0:0] h_u_arrmul24_fa6_12_xor1;
  wire [0:0] h_u_arrmul24_fa6_12_or0;
  wire [0:0] h_u_arrmul24_and7_12;
  wire [0:0] h_u_arrmul24_fa7_12_xor1;
  wire [0:0] h_u_arrmul24_fa7_12_or0;
  wire [0:0] h_u_arrmul24_and8_12;
  wire [0:0] h_u_arrmul24_fa8_12_xor1;
  wire [0:0] h_u_arrmul24_fa8_12_or0;
  wire [0:0] h_u_arrmul24_and9_12;
  wire [0:0] h_u_arrmul24_fa9_12_xor1;
  wire [0:0] h_u_arrmul24_fa9_12_or0;
  wire [0:0] h_u_arrmul24_and10_12;
  wire [0:0] h_u_arrmul24_fa10_12_xor1;
  wire [0:0] h_u_arrmul24_fa10_12_or0;
  wire [0:0] h_u_arrmul24_and11_12;
  wire [0:0] h_u_arrmul24_fa11_12_xor1;
  wire [0:0] h_u_arrmul24_fa11_12_or0;
  wire [0:0] h_u_arrmul24_and12_12;
  wire [0:0] h_u_arrmul24_fa12_12_xor1;
  wire [0:0] h_u_arrmul24_fa12_12_or0;
  wire [0:0] h_u_arrmul24_and13_12;
  wire [0:0] h_u_arrmul24_fa13_12_xor1;
  wire [0:0] h_u_arrmul24_fa13_12_or0;
  wire [0:0] h_u_arrmul24_and14_12;
  wire [0:0] h_u_arrmul24_fa14_12_xor1;
  wire [0:0] h_u_arrmul24_fa14_12_or0;
  wire [0:0] h_u_arrmul24_and15_12;
  wire [0:0] h_u_arrmul24_fa15_12_xor1;
  wire [0:0] h_u_arrmul24_fa15_12_or0;
  wire [0:0] h_u_arrmul24_and16_12;
  wire [0:0] h_u_arrmul24_fa16_12_xor1;
  wire [0:0] h_u_arrmul24_fa16_12_or0;
  wire [0:0] h_u_arrmul24_and17_12;
  wire [0:0] h_u_arrmul24_fa17_12_xor1;
  wire [0:0] h_u_arrmul24_fa17_12_or0;
  wire [0:0] h_u_arrmul24_and18_12;
  wire [0:0] h_u_arrmul24_fa18_12_xor1;
  wire [0:0] h_u_arrmul24_fa18_12_or0;
  wire [0:0] h_u_arrmul24_and19_12;
  wire [0:0] h_u_arrmul24_fa19_12_xor1;
  wire [0:0] h_u_arrmul24_fa19_12_or0;
  wire [0:0] h_u_arrmul24_and20_12;
  wire [0:0] h_u_arrmul24_fa20_12_xor1;
  wire [0:0] h_u_arrmul24_fa20_12_or0;
  wire [0:0] h_u_arrmul24_and21_12;
  wire [0:0] h_u_arrmul24_fa21_12_xor1;
  wire [0:0] h_u_arrmul24_fa21_12_or0;
  wire [0:0] h_u_arrmul24_and22_12;
  wire [0:0] h_u_arrmul24_fa22_12_xor1;
  wire [0:0] h_u_arrmul24_fa22_12_or0;
  wire [0:0] h_u_arrmul24_and23_12;
  wire [0:0] h_u_arrmul24_fa23_12_xor1;
  wire [0:0] h_u_arrmul24_fa23_12_or0;
  wire [0:0] h_u_arrmul24_and0_13;
  wire [0:0] h_u_arrmul24_ha0_13_xor0;
  wire [0:0] h_u_arrmul24_ha0_13_and0;
  wire [0:0] h_u_arrmul24_and1_13;
  wire [0:0] h_u_arrmul24_fa1_13_xor1;
  wire [0:0] h_u_arrmul24_fa1_13_or0;
  wire [0:0] h_u_arrmul24_and2_13;
  wire [0:0] h_u_arrmul24_fa2_13_xor1;
  wire [0:0] h_u_arrmul24_fa2_13_or0;
  wire [0:0] h_u_arrmul24_and3_13;
  wire [0:0] h_u_arrmul24_fa3_13_xor1;
  wire [0:0] h_u_arrmul24_fa3_13_or0;
  wire [0:0] h_u_arrmul24_and4_13;
  wire [0:0] h_u_arrmul24_fa4_13_xor1;
  wire [0:0] h_u_arrmul24_fa4_13_or0;
  wire [0:0] h_u_arrmul24_and5_13;
  wire [0:0] h_u_arrmul24_fa5_13_xor1;
  wire [0:0] h_u_arrmul24_fa5_13_or0;
  wire [0:0] h_u_arrmul24_and6_13;
  wire [0:0] h_u_arrmul24_fa6_13_xor1;
  wire [0:0] h_u_arrmul24_fa6_13_or0;
  wire [0:0] h_u_arrmul24_and7_13;
  wire [0:0] h_u_arrmul24_fa7_13_xor1;
  wire [0:0] h_u_arrmul24_fa7_13_or0;
  wire [0:0] h_u_arrmul24_and8_13;
  wire [0:0] h_u_arrmul24_fa8_13_xor1;
  wire [0:0] h_u_arrmul24_fa8_13_or0;
  wire [0:0] h_u_arrmul24_and9_13;
  wire [0:0] h_u_arrmul24_fa9_13_xor1;
  wire [0:0] h_u_arrmul24_fa9_13_or0;
  wire [0:0] h_u_arrmul24_and10_13;
  wire [0:0] h_u_arrmul24_fa10_13_xor1;
  wire [0:0] h_u_arrmul24_fa10_13_or0;
  wire [0:0] h_u_arrmul24_and11_13;
  wire [0:0] h_u_arrmul24_fa11_13_xor1;
  wire [0:0] h_u_arrmul24_fa11_13_or0;
  wire [0:0] h_u_arrmul24_and12_13;
  wire [0:0] h_u_arrmul24_fa12_13_xor1;
  wire [0:0] h_u_arrmul24_fa12_13_or0;
  wire [0:0] h_u_arrmul24_and13_13;
  wire [0:0] h_u_arrmul24_fa13_13_xor1;
  wire [0:0] h_u_arrmul24_fa13_13_or0;
  wire [0:0] h_u_arrmul24_and14_13;
  wire [0:0] h_u_arrmul24_fa14_13_xor1;
  wire [0:0] h_u_arrmul24_fa14_13_or0;
  wire [0:0] h_u_arrmul24_and15_13;
  wire [0:0] h_u_arrmul24_fa15_13_xor1;
  wire [0:0] h_u_arrmul24_fa15_13_or0;
  wire [0:0] h_u_arrmul24_and16_13;
  wire [0:0] h_u_arrmul24_fa16_13_xor1;
  wire [0:0] h_u_arrmul24_fa16_13_or0;
  wire [0:0] h_u_arrmul24_and17_13;
  wire [0:0] h_u_arrmul24_fa17_13_xor1;
  wire [0:0] h_u_arrmul24_fa17_13_or0;
  wire [0:0] h_u_arrmul24_and18_13;
  wire [0:0] h_u_arrmul24_fa18_13_xor1;
  wire [0:0] h_u_arrmul24_fa18_13_or0;
  wire [0:0] h_u_arrmul24_and19_13;
  wire [0:0] h_u_arrmul24_fa19_13_xor1;
  wire [0:0] h_u_arrmul24_fa19_13_or0;
  wire [0:0] h_u_arrmul24_and20_13;
  wire [0:0] h_u_arrmul24_fa20_13_xor1;
  wire [0:0] h_u_arrmul24_fa20_13_or0;
  wire [0:0] h_u_arrmul24_and21_13;
  wire [0:0] h_u_arrmul24_fa21_13_xor1;
  wire [0:0] h_u_arrmul24_fa21_13_or0;
  wire [0:0] h_u_arrmul24_and22_13;
  wire [0:0] h_u_arrmul24_fa22_13_xor1;
  wire [0:0] h_u_arrmul24_fa22_13_or0;
  wire [0:0] h_u_arrmul24_and23_13;
  wire [0:0] h_u_arrmul24_fa23_13_xor1;
  wire [0:0] h_u_arrmul24_fa23_13_or0;
  wire [0:0] h_u_arrmul24_and0_14;
  wire [0:0] h_u_arrmul24_ha0_14_xor0;
  wire [0:0] h_u_arrmul24_ha0_14_and0;
  wire [0:0] h_u_arrmul24_and1_14;
  wire [0:0] h_u_arrmul24_fa1_14_xor1;
  wire [0:0] h_u_arrmul24_fa1_14_or0;
  wire [0:0] h_u_arrmul24_and2_14;
  wire [0:0] h_u_arrmul24_fa2_14_xor1;
  wire [0:0] h_u_arrmul24_fa2_14_or0;
  wire [0:0] h_u_arrmul24_and3_14;
  wire [0:0] h_u_arrmul24_fa3_14_xor1;
  wire [0:0] h_u_arrmul24_fa3_14_or0;
  wire [0:0] h_u_arrmul24_and4_14;
  wire [0:0] h_u_arrmul24_fa4_14_xor1;
  wire [0:0] h_u_arrmul24_fa4_14_or0;
  wire [0:0] h_u_arrmul24_and5_14;
  wire [0:0] h_u_arrmul24_fa5_14_xor1;
  wire [0:0] h_u_arrmul24_fa5_14_or0;
  wire [0:0] h_u_arrmul24_and6_14;
  wire [0:0] h_u_arrmul24_fa6_14_xor1;
  wire [0:0] h_u_arrmul24_fa6_14_or0;
  wire [0:0] h_u_arrmul24_and7_14;
  wire [0:0] h_u_arrmul24_fa7_14_xor1;
  wire [0:0] h_u_arrmul24_fa7_14_or0;
  wire [0:0] h_u_arrmul24_and8_14;
  wire [0:0] h_u_arrmul24_fa8_14_xor1;
  wire [0:0] h_u_arrmul24_fa8_14_or0;
  wire [0:0] h_u_arrmul24_and9_14;
  wire [0:0] h_u_arrmul24_fa9_14_xor1;
  wire [0:0] h_u_arrmul24_fa9_14_or0;
  wire [0:0] h_u_arrmul24_and10_14;
  wire [0:0] h_u_arrmul24_fa10_14_xor1;
  wire [0:0] h_u_arrmul24_fa10_14_or0;
  wire [0:0] h_u_arrmul24_and11_14;
  wire [0:0] h_u_arrmul24_fa11_14_xor1;
  wire [0:0] h_u_arrmul24_fa11_14_or0;
  wire [0:0] h_u_arrmul24_and12_14;
  wire [0:0] h_u_arrmul24_fa12_14_xor1;
  wire [0:0] h_u_arrmul24_fa12_14_or0;
  wire [0:0] h_u_arrmul24_and13_14;
  wire [0:0] h_u_arrmul24_fa13_14_xor1;
  wire [0:0] h_u_arrmul24_fa13_14_or0;
  wire [0:0] h_u_arrmul24_and14_14;
  wire [0:0] h_u_arrmul24_fa14_14_xor1;
  wire [0:0] h_u_arrmul24_fa14_14_or0;
  wire [0:0] h_u_arrmul24_and15_14;
  wire [0:0] h_u_arrmul24_fa15_14_xor1;
  wire [0:0] h_u_arrmul24_fa15_14_or0;
  wire [0:0] h_u_arrmul24_and16_14;
  wire [0:0] h_u_arrmul24_fa16_14_xor1;
  wire [0:0] h_u_arrmul24_fa16_14_or0;
  wire [0:0] h_u_arrmul24_and17_14;
  wire [0:0] h_u_arrmul24_fa17_14_xor1;
  wire [0:0] h_u_arrmul24_fa17_14_or0;
  wire [0:0] h_u_arrmul24_and18_14;
  wire [0:0] h_u_arrmul24_fa18_14_xor1;
  wire [0:0] h_u_arrmul24_fa18_14_or0;
  wire [0:0] h_u_arrmul24_and19_14;
  wire [0:0] h_u_arrmul24_fa19_14_xor1;
  wire [0:0] h_u_arrmul24_fa19_14_or0;
  wire [0:0] h_u_arrmul24_and20_14;
  wire [0:0] h_u_arrmul24_fa20_14_xor1;
  wire [0:0] h_u_arrmul24_fa20_14_or0;
  wire [0:0] h_u_arrmul24_and21_14;
  wire [0:0] h_u_arrmul24_fa21_14_xor1;
  wire [0:0] h_u_arrmul24_fa21_14_or0;
  wire [0:0] h_u_arrmul24_and22_14;
  wire [0:0] h_u_arrmul24_fa22_14_xor1;
  wire [0:0] h_u_arrmul24_fa22_14_or0;
  wire [0:0] h_u_arrmul24_and23_14;
  wire [0:0] h_u_arrmul24_fa23_14_xor1;
  wire [0:0] h_u_arrmul24_fa23_14_or0;
  wire [0:0] h_u_arrmul24_and0_15;
  wire [0:0] h_u_arrmul24_ha0_15_xor0;
  wire [0:0] h_u_arrmul24_ha0_15_and0;
  wire [0:0] h_u_arrmul24_and1_15;
  wire [0:0] h_u_arrmul24_fa1_15_xor1;
  wire [0:0] h_u_arrmul24_fa1_15_or0;
  wire [0:0] h_u_arrmul24_and2_15;
  wire [0:0] h_u_arrmul24_fa2_15_xor1;
  wire [0:0] h_u_arrmul24_fa2_15_or0;
  wire [0:0] h_u_arrmul24_and3_15;
  wire [0:0] h_u_arrmul24_fa3_15_xor1;
  wire [0:0] h_u_arrmul24_fa3_15_or0;
  wire [0:0] h_u_arrmul24_and4_15;
  wire [0:0] h_u_arrmul24_fa4_15_xor1;
  wire [0:0] h_u_arrmul24_fa4_15_or0;
  wire [0:0] h_u_arrmul24_and5_15;
  wire [0:0] h_u_arrmul24_fa5_15_xor1;
  wire [0:0] h_u_arrmul24_fa5_15_or0;
  wire [0:0] h_u_arrmul24_and6_15;
  wire [0:0] h_u_arrmul24_fa6_15_xor1;
  wire [0:0] h_u_arrmul24_fa6_15_or0;
  wire [0:0] h_u_arrmul24_and7_15;
  wire [0:0] h_u_arrmul24_fa7_15_xor1;
  wire [0:0] h_u_arrmul24_fa7_15_or0;
  wire [0:0] h_u_arrmul24_and8_15;
  wire [0:0] h_u_arrmul24_fa8_15_xor1;
  wire [0:0] h_u_arrmul24_fa8_15_or0;
  wire [0:0] h_u_arrmul24_and9_15;
  wire [0:0] h_u_arrmul24_fa9_15_xor1;
  wire [0:0] h_u_arrmul24_fa9_15_or0;
  wire [0:0] h_u_arrmul24_and10_15;
  wire [0:0] h_u_arrmul24_fa10_15_xor1;
  wire [0:0] h_u_arrmul24_fa10_15_or0;
  wire [0:0] h_u_arrmul24_and11_15;
  wire [0:0] h_u_arrmul24_fa11_15_xor1;
  wire [0:0] h_u_arrmul24_fa11_15_or0;
  wire [0:0] h_u_arrmul24_and12_15;
  wire [0:0] h_u_arrmul24_fa12_15_xor1;
  wire [0:0] h_u_arrmul24_fa12_15_or0;
  wire [0:0] h_u_arrmul24_and13_15;
  wire [0:0] h_u_arrmul24_fa13_15_xor1;
  wire [0:0] h_u_arrmul24_fa13_15_or0;
  wire [0:0] h_u_arrmul24_and14_15;
  wire [0:0] h_u_arrmul24_fa14_15_xor1;
  wire [0:0] h_u_arrmul24_fa14_15_or0;
  wire [0:0] h_u_arrmul24_and15_15;
  wire [0:0] h_u_arrmul24_fa15_15_xor1;
  wire [0:0] h_u_arrmul24_fa15_15_or0;
  wire [0:0] h_u_arrmul24_and16_15;
  wire [0:0] h_u_arrmul24_fa16_15_xor1;
  wire [0:0] h_u_arrmul24_fa16_15_or0;
  wire [0:0] h_u_arrmul24_and17_15;
  wire [0:0] h_u_arrmul24_fa17_15_xor1;
  wire [0:0] h_u_arrmul24_fa17_15_or0;
  wire [0:0] h_u_arrmul24_and18_15;
  wire [0:0] h_u_arrmul24_fa18_15_xor1;
  wire [0:0] h_u_arrmul24_fa18_15_or0;
  wire [0:0] h_u_arrmul24_and19_15;
  wire [0:0] h_u_arrmul24_fa19_15_xor1;
  wire [0:0] h_u_arrmul24_fa19_15_or0;
  wire [0:0] h_u_arrmul24_and20_15;
  wire [0:0] h_u_arrmul24_fa20_15_xor1;
  wire [0:0] h_u_arrmul24_fa20_15_or0;
  wire [0:0] h_u_arrmul24_and21_15;
  wire [0:0] h_u_arrmul24_fa21_15_xor1;
  wire [0:0] h_u_arrmul24_fa21_15_or0;
  wire [0:0] h_u_arrmul24_and22_15;
  wire [0:0] h_u_arrmul24_fa22_15_xor1;
  wire [0:0] h_u_arrmul24_fa22_15_or0;
  wire [0:0] h_u_arrmul24_and23_15;
  wire [0:0] h_u_arrmul24_fa23_15_xor1;
  wire [0:0] h_u_arrmul24_fa23_15_or0;
  wire [0:0] h_u_arrmul24_and0_16;
  wire [0:0] h_u_arrmul24_ha0_16_xor0;
  wire [0:0] h_u_arrmul24_ha0_16_and0;
  wire [0:0] h_u_arrmul24_and1_16;
  wire [0:0] h_u_arrmul24_fa1_16_xor1;
  wire [0:0] h_u_arrmul24_fa1_16_or0;
  wire [0:0] h_u_arrmul24_and2_16;
  wire [0:0] h_u_arrmul24_fa2_16_xor1;
  wire [0:0] h_u_arrmul24_fa2_16_or0;
  wire [0:0] h_u_arrmul24_and3_16;
  wire [0:0] h_u_arrmul24_fa3_16_xor1;
  wire [0:0] h_u_arrmul24_fa3_16_or0;
  wire [0:0] h_u_arrmul24_and4_16;
  wire [0:0] h_u_arrmul24_fa4_16_xor1;
  wire [0:0] h_u_arrmul24_fa4_16_or0;
  wire [0:0] h_u_arrmul24_and5_16;
  wire [0:0] h_u_arrmul24_fa5_16_xor1;
  wire [0:0] h_u_arrmul24_fa5_16_or0;
  wire [0:0] h_u_arrmul24_and6_16;
  wire [0:0] h_u_arrmul24_fa6_16_xor1;
  wire [0:0] h_u_arrmul24_fa6_16_or0;
  wire [0:0] h_u_arrmul24_and7_16;
  wire [0:0] h_u_arrmul24_fa7_16_xor1;
  wire [0:0] h_u_arrmul24_fa7_16_or0;
  wire [0:0] h_u_arrmul24_and8_16;
  wire [0:0] h_u_arrmul24_fa8_16_xor1;
  wire [0:0] h_u_arrmul24_fa8_16_or0;
  wire [0:0] h_u_arrmul24_and9_16;
  wire [0:0] h_u_arrmul24_fa9_16_xor1;
  wire [0:0] h_u_arrmul24_fa9_16_or0;
  wire [0:0] h_u_arrmul24_and10_16;
  wire [0:0] h_u_arrmul24_fa10_16_xor1;
  wire [0:0] h_u_arrmul24_fa10_16_or0;
  wire [0:0] h_u_arrmul24_and11_16;
  wire [0:0] h_u_arrmul24_fa11_16_xor1;
  wire [0:0] h_u_arrmul24_fa11_16_or0;
  wire [0:0] h_u_arrmul24_and12_16;
  wire [0:0] h_u_arrmul24_fa12_16_xor1;
  wire [0:0] h_u_arrmul24_fa12_16_or0;
  wire [0:0] h_u_arrmul24_and13_16;
  wire [0:0] h_u_arrmul24_fa13_16_xor1;
  wire [0:0] h_u_arrmul24_fa13_16_or0;
  wire [0:0] h_u_arrmul24_and14_16;
  wire [0:0] h_u_arrmul24_fa14_16_xor1;
  wire [0:0] h_u_arrmul24_fa14_16_or0;
  wire [0:0] h_u_arrmul24_and15_16;
  wire [0:0] h_u_arrmul24_fa15_16_xor1;
  wire [0:0] h_u_arrmul24_fa15_16_or0;
  wire [0:0] h_u_arrmul24_and16_16;
  wire [0:0] h_u_arrmul24_fa16_16_xor1;
  wire [0:0] h_u_arrmul24_fa16_16_or0;
  wire [0:0] h_u_arrmul24_and17_16;
  wire [0:0] h_u_arrmul24_fa17_16_xor1;
  wire [0:0] h_u_arrmul24_fa17_16_or0;
  wire [0:0] h_u_arrmul24_and18_16;
  wire [0:0] h_u_arrmul24_fa18_16_xor1;
  wire [0:0] h_u_arrmul24_fa18_16_or0;
  wire [0:0] h_u_arrmul24_and19_16;
  wire [0:0] h_u_arrmul24_fa19_16_xor1;
  wire [0:0] h_u_arrmul24_fa19_16_or0;
  wire [0:0] h_u_arrmul24_and20_16;
  wire [0:0] h_u_arrmul24_fa20_16_xor1;
  wire [0:0] h_u_arrmul24_fa20_16_or0;
  wire [0:0] h_u_arrmul24_and21_16;
  wire [0:0] h_u_arrmul24_fa21_16_xor1;
  wire [0:0] h_u_arrmul24_fa21_16_or0;
  wire [0:0] h_u_arrmul24_and22_16;
  wire [0:0] h_u_arrmul24_fa22_16_xor1;
  wire [0:0] h_u_arrmul24_fa22_16_or0;
  wire [0:0] h_u_arrmul24_and23_16;
  wire [0:0] h_u_arrmul24_fa23_16_xor1;
  wire [0:0] h_u_arrmul24_fa23_16_or0;
  wire [0:0] h_u_arrmul24_and0_17;
  wire [0:0] h_u_arrmul24_ha0_17_xor0;
  wire [0:0] h_u_arrmul24_ha0_17_and0;
  wire [0:0] h_u_arrmul24_and1_17;
  wire [0:0] h_u_arrmul24_fa1_17_xor1;
  wire [0:0] h_u_arrmul24_fa1_17_or0;
  wire [0:0] h_u_arrmul24_and2_17;
  wire [0:0] h_u_arrmul24_fa2_17_xor1;
  wire [0:0] h_u_arrmul24_fa2_17_or0;
  wire [0:0] h_u_arrmul24_and3_17;
  wire [0:0] h_u_arrmul24_fa3_17_xor1;
  wire [0:0] h_u_arrmul24_fa3_17_or0;
  wire [0:0] h_u_arrmul24_and4_17;
  wire [0:0] h_u_arrmul24_fa4_17_xor1;
  wire [0:0] h_u_arrmul24_fa4_17_or0;
  wire [0:0] h_u_arrmul24_and5_17;
  wire [0:0] h_u_arrmul24_fa5_17_xor1;
  wire [0:0] h_u_arrmul24_fa5_17_or0;
  wire [0:0] h_u_arrmul24_and6_17;
  wire [0:0] h_u_arrmul24_fa6_17_xor1;
  wire [0:0] h_u_arrmul24_fa6_17_or0;
  wire [0:0] h_u_arrmul24_and7_17;
  wire [0:0] h_u_arrmul24_fa7_17_xor1;
  wire [0:0] h_u_arrmul24_fa7_17_or0;
  wire [0:0] h_u_arrmul24_and8_17;
  wire [0:0] h_u_arrmul24_fa8_17_xor1;
  wire [0:0] h_u_arrmul24_fa8_17_or0;
  wire [0:0] h_u_arrmul24_and9_17;
  wire [0:0] h_u_arrmul24_fa9_17_xor1;
  wire [0:0] h_u_arrmul24_fa9_17_or0;
  wire [0:0] h_u_arrmul24_and10_17;
  wire [0:0] h_u_arrmul24_fa10_17_xor1;
  wire [0:0] h_u_arrmul24_fa10_17_or0;
  wire [0:0] h_u_arrmul24_and11_17;
  wire [0:0] h_u_arrmul24_fa11_17_xor1;
  wire [0:0] h_u_arrmul24_fa11_17_or0;
  wire [0:0] h_u_arrmul24_and12_17;
  wire [0:0] h_u_arrmul24_fa12_17_xor1;
  wire [0:0] h_u_arrmul24_fa12_17_or0;
  wire [0:0] h_u_arrmul24_and13_17;
  wire [0:0] h_u_arrmul24_fa13_17_xor1;
  wire [0:0] h_u_arrmul24_fa13_17_or0;
  wire [0:0] h_u_arrmul24_and14_17;
  wire [0:0] h_u_arrmul24_fa14_17_xor1;
  wire [0:0] h_u_arrmul24_fa14_17_or0;
  wire [0:0] h_u_arrmul24_and15_17;
  wire [0:0] h_u_arrmul24_fa15_17_xor1;
  wire [0:0] h_u_arrmul24_fa15_17_or0;
  wire [0:0] h_u_arrmul24_and16_17;
  wire [0:0] h_u_arrmul24_fa16_17_xor1;
  wire [0:0] h_u_arrmul24_fa16_17_or0;
  wire [0:0] h_u_arrmul24_and17_17;
  wire [0:0] h_u_arrmul24_fa17_17_xor1;
  wire [0:0] h_u_arrmul24_fa17_17_or0;
  wire [0:0] h_u_arrmul24_and18_17;
  wire [0:0] h_u_arrmul24_fa18_17_xor1;
  wire [0:0] h_u_arrmul24_fa18_17_or0;
  wire [0:0] h_u_arrmul24_and19_17;
  wire [0:0] h_u_arrmul24_fa19_17_xor1;
  wire [0:0] h_u_arrmul24_fa19_17_or0;
  wire [0:0] h_u_arrmul24_and20_17;
  wire [0:0] h_u_arrmul24_fa20_17_xor1;
  wire [0:0] h_u_arrmul24_fa20_17_or0;
  wire [0:0] h_u_arrmul24_and21_17;
  wire [0:0] h_u_arrmul24_fa21_17_xor1;
  wire [0:0] h_u_arrmul24_fa21_17_or0;
  wire [0:0] h_u_arrmul24_and22_17;
  wire [0:0] h_u_arrmul24_fa22_17_xor1;
  wire [0:0] h_u_arrmul24_fa22_17_or0;
  wire [0:0] h_u_arrmul24_and23_17;
  wire [0:0] h_u_arrmul24_fa23_17_xor1;
  wire [0:0] h_u_arrmul24_fa23_17_or0;
  wire [0:0] h_u_arrmul24_and0_18;
  wire [0:0] h_u_arrmul24_ha0_18_xor0;
  wire [0:0] h_u_arrmul24_ha0_18_and0;
  wire [0:0] h_u_arrmul24_and1_18;
  wire [0:0] h_u_arrmul24_fa1_18_xor1;
  wire [0:0] h_u_arrmul24_fa1_18_or0;
  wire [0:0] h_u_arrmul24_and2_18;
  wire [0:0] h_u_arrmul24_fa2_18_xor1;
  wire [0:0] h_u_arrmul24_fa2_18_or0;
  wire [0:0] h_u_arrmul24_and3_18;
  wire [0:0] h_u_arrmul24_fa3_18_xor1;
  wire [0:0] h_u_arrmul24_fa3_18_or0;
  wire [0:0] h_u_arrmul24_and4_18;
  wire [0:0] h_u_arrmul24_fa4_18_xor1;
  wire [0:0] h_u_arrmul24_fa4_18_or0;
  wire [0:0] h_u_arrmul24_and5_18;
  wire [0:0] h_u_arrmul24_fa5_18_xor1;
  wire [0:0] h_u_arrmul24_fa5_18_or0;
  wire [0:0] h_u_arrmul24_and6_18;
  wire [0:0] h_u_arrmul24_fa6_18_xor1;
  wire [0:0] h_u_arrmul24_fa6_18_or0;
  wire [0:0] h_u_arrmul24_and7_18;
  wire [0:0] h_u_arrmul24_fa7_18_xor1;
  wire [0:0] h_u_arrmul24_fa7_18_or0;
  wire [0:0] h_u_arrmul24_and8_18;
  wire [0:0] h_u_arrmul24_fa8_18_xor1;
  wire [0:0] h_u_arrmul24_fa8_18_or0;
  wire [0:0] h_u_arrmul24_and9_18;
  wire [0:0] h_u_arrmul24_fa9_18_xor1;
  wire [0:0] h_u_arrmul24_fa9_18_or0;
  wire [0:0] h_u_arrmul24_and10_18;
  wire [0:0] h_u_arrmul24_fa10_18_xor1;
  wire [0:0] h_u_arrmul24_fa10_18_or0;
  wire [0:0] h_u_arrmul24_and11_18;
  wire [0:0] h_u_arrmul24_fa11_18_xor1;
  wire [0:0] h_u_arrmul24_fa11_18_or0;
  wire [0:0] h_u_arrmul24_and12_18;
  wire [0:0] h_u_arrmul24_fa12_18_xor1;
  wire [0:0] h_u_arrmul24_fa12_18_or0;
  wire [0:0] h_u_arrmul24_and13_18;
  wire [0:0] h_u_arrmul24_fa13_18_xor1;
  wire [0:0] h_u_arrmul24_fa13_18_or0;
  wire [0:0] h_u_arrmul24_and14_18;
  wire [0:0] h_u_arrmul24_fa14_18_xor1;
  wire [0:0] h_u_arrmul24_fa14_18_or0;
  wire [0:0] h_u_arrmul24_and15_18;
  wire [0:0] h_u_arrmul24_fa15_18_xor1;
  wire [0:0] h_u_arrmul24_fa15_18_or0;
  wire [0:0] h_u_arrmul24_and16_18;
  wire [0:0] h_u_arrmul24_fa16_18_xor1;
  wire [0:0] h_u_arrmul24_fa16_18_or0;
  wire [0:0] h_u_arrmul24_and17_18;
  wire [0:0] h_u_arrmul24_fa17_18_xor1;
  wire [0:0] h_u_arrmul24_fa17_18_or0;
  wire [0:0] h_u_arrmul24_and18_18;
  wire [0:0] h_u_arrmul24_fa18_18_xor1;
  wire [0:0] h_u_arrmul24_fa18_18_or0;
  wire [0:0] h_u_arrmul24_and19_18;
  wire [0:0] h_u_arrmul24_fa19_18_xor1;
  wire [0:0] h_u_arrmul24_fa19_18_or0;
  wire [0:0] h_u_arrmul24_and20_18;
  wire [0:0] h_u_arrmul24_fa20_18_xor1;
  wire [0:0] h_u_arrmul24_fa20_18_or0;
  wire [0:0] h_u_arrmul24_and21_18;
  wire [0:0] h_u_arrmul24_fa21_18_xor1;
  wire [0:0] h_u_arrmul24_fa21_18_or0;
  wire [0:0] h_u_arrmul24_and22_18;
  wire [0:0] h_u_arrmul24_fa22_18_xor1;
  wire [0:0] h_u_arrmul24_fa22_18_or0;
  wire [0:0] h_u_arrmul24_and23_18;
  wire [0:0] h_u_arrmul24_fa23_18_xor1;
  wire [0:0] h_u_arrmul24_fa23_18_or0;
  wire [0:0] h_u_arrmul24_and0_19;
  wire [0:0] h_u_arrmul24_ha0_19_xor0;
  wire [0:0] h_u_arrmul24_ha0_19_and0;
  wire [0:0] h_u_arrmul24_and1_19;
  wire [0:0] h_u_arrmul24_fa1_19_xor1;
  wire [0:0] h_u_arrmul24_fa1_19_or0;
  wire [0:0] h_u_arrmul24_and2_19;
  wire [0:0] h_u_arrmul24_fa2_19_xor1;
  wire [0:0] h_u_arrmul24_fa2_19_or0;
  wire [0:0] h_u_arrmul24_and3_19;
  wire [0:0] h_u_arrmul24_fa3_19_xor1;
  wire [0:0] h_u_arrmul24_fa3_19_or0;
  wire [0:0] h_u_arrmul24_and4_19;
  wire [0:0] h_u_arrmul24_fa4_19_xor1;
  wire [0:0] h_u_arrmul24_fa4_19_or0;
  wire [0:0] h_u_arrmul24_and5_19;
  wire [0:0] h_u_arrmul24_fa5_19_xor1;
  wire [0:0] h_u_arrmul24_fa5_19_or0;
  wire [0:0] h_u_arrmul24_and6_19;
  wire [0:0] h_u_arrmul24_fa6_19_xor1;
  wire [0:0] h_u_arrmul24_fa6_19_or0;
  wire [0:0] h_u_arrmul24_and7_19;
  wire [0:0] h_u_arrmul24_fa7_19_xor1;
  wire [0:0] h_u_arrmul24_fa7_19_or0;
  wire [0:0] h_u_arrmul24_and8_19;
  wire [0:0] h_u_arrmul24_fa8_19_xor1;
  wire [0:0] h_u_arrmul24_fa8_19_or0;
  wire [0:0] h_u_arrmul24_and9_19;
  wire [0:0] h_u_arrmul24_fa9_19_xor1;
  wire [0:0] h_u_arrmul24_fa9_19_or0;
  wire [0:0] h_u_arrmul24_and10_19;
  wire [0:0] h_u_arrmul24_fa10_19_xor1;
  wire [0:0] h_u_arrmul24_fa10_19_or0;
  wire [0:0] h_u_arrmul24_and11_19;
  wire [0:0] h_u_arrmul24_fa11_19_xor1;
  wire [0:0] h_u_arrmul24_fa11_19_or0;
  wire [0:0] h_u_arrmul24_and12_19;
  wire [0:0] h_u_arrmul24_fa12_19_xor1;
  wire [0:0] h_u_arrmul24_fa12_19_or0;
  wire [0:0] h_u_arrmul24_and13_19;
  wire [0:0] h_u_arrmul24_fa13_19_xor1;
  wire [0:0] h_u_arrmul24_fa13_19_or0;
  wire [0:0] h_u_arrmul24_and14_19;
  wire [0:0] h_u_arrmul24_fa14_19_xor1;
  wire [0:0] h_u_arrmul24_fa14_19_or0;
  wire [0:0] h_u_arrmul24_and15_19;
  wire [0:0] h_u_arrmul24_fa15_19_xor1;
  wire [0:0] h_u_arrmul24_fa15_19_or0;
  wire [0:0] h_u_arrmul24_and16_19;
  wire [0:0] h_u_arrmul24_fa16_19_xor1;
  wire [0:0] h_u_arrmul24_fa16_19_or0;
  wire [0:0] h_u_arrmul24_and17_19;
  wire [0:0] h_u_arrmul24_fa17_19_xor1;
  wire [0:0] h_u_arrmul24_fa17_19_or0;
  wire [0:0] h_u_arrmul24_and18_19;
  wire [0:0] h_u_arrmul24_fa18_19_xor1;
  wire [0:0] h_u_arrmul24_fa18_19_or0;
  wire [0:0] h_u_arrmul24_and19_19;
  wire [0:0] h_u_arrmul24_fa19_19_xor1;
  wire [0:0] h_u_arrmul24_fa19_19_or0;
  wire [0:0] h_u_arrmul24_and20_19;
  wire [0:0] h_u_arrmul24_fa20_19_xor1;
  wire [0:0] h_u_arrmul24_fa20_19_or0;
  wire [0:0] h_u_arrmul24_and21_19;
  wire [0:0] h_u_arrmul24_fa21_19_xor1;
  wire [0:0] h_u_arrmul24_fa21_19_or0;
  wire [0:0] h_u_arrmul24_and22_19;
  wire [0:0] h_u_arrmul24_fa22_19_xor1;
  wire [0:0] h_u_arrmul24_fa22_19_or0;
  wire [0:0] h_u_arrmul24_and23_19;
  wire [0:0] h_u_arrmul24_fa23_19_xor1;
  wire [0:0] h_u_arrmul24_fa23_19_or0;
  wire [0:0] h_u_arrmul24_and0_20;
  wire [0:0] h_u_arrmul24_ha0_20_xor0;
  wire [0:0] h_u_arrmul24_ha0_20_and0;
  wire [0:0] h_u_arrmul24_and1_20;
  wire [0:0] h_u_arrmul24_fa1_20_xor1;
  wire [0:0] h_u_arrmul24_fa1_20_or0;
  wire [0:0] h_u_arrmul24_and2_20;
  wire [0:0] h_u_arrmul24_fa2_20_xor1;
  wire [0:0] h_u_arrmul24_fa2_20_or0;
  wire [0:0] h_u_arrmul24_and3_20;
  wire [0:0] h_u_arrmul24_fa3_20_xor1;
  wire [0:0] h_u_arrmul24_fa3_20_or0;
  wire [0:0] h_u_arrmul24_and4_20;
  wire [0:0] h_u_arrmul24_fa4_20_xor1;
  wire [0:0] h_u_arrmul24_fa4_20_or0;
  wire [0:0] h_u_arrmul24_and5_20;
  wire [0:0] h_u_arrmul24_fa5_20_xor1;
  wire [0:0] h_u_arrmul24_fa5_20_or0;
  wire [0:0] h_u_arrmul24_and6_20;
  wire [0:0] h_u_arrmul24_fa6_20_xor1;
  wire [0:0] h_u_arrmul24_fa6_20_or0;
  wire [0:0] h_u_arrmul24_and7_20;
  wire [0:0] h_u_arrmul24_fa7_20_xor1;
  wire [0:0] h_u_arrmul24_fa7_20_or0;
  wire [0:0] h_u_arrmul24_and8_20;
  wire [0:0] h_u_arrmul24_fa8_20_xor1;
  wire [0:0] h_u_arrmul24_fa8_20_or0;
  wire [0:0] h_u_arrmul24_and9_20;
  wire [0:0] h_u_arrmul24_fa9_20_xor1;
  wire [0:0] h_u_arrmul24_fa9_20_or0;
  wire [0:0] h_u_arrmul24_and10_20;
  wire [0:0] h_u_arrmul24_fa10_20_xor1;
  wire [0:0] h_u_arrmul24_fa10_20_or0;
  wire [0:0] h_u_arrmul24_and11_20;
  wire [0:0] h_u_arrmul24_fa11_20_xor1;
  wire [0:0] h_u_arrmul24_fa11_20_or0;
  wire [0:0] h_u_arrmul24_and12_20;
  wire [0:0] h_u_arrmul24_fa12_20_xor1;
  wire [0:0] h_u_arrmul24_fa12_20_or0;
  wire [0:0] h_u_arrmul24_and13_20;
  wire [0:0] h_u_arrmul24_fa13_20_xor1;
  wire [0:0] h_u_arrmul24_fa13_20_or0;
  wire [0:0] h_u_arrmul24_and14_20;
  wire [0:0] h_u_arrmul24_fa14_20_xor1;
  wire [0:0] h_u_arrmul24_fa14_20_or0;
  wire [0:0] h_u_arrmul24_and15_20;
  wire [0:0] h_u_arrmul24_fa15_20_xor1;
  wire [0:0] h_u_arrmul24_fa15_20_or0;
  wire [0:0] h_u_arrmul24_and16_20;
  wire [0:0] h_u_arrmul24_fa16_20_xor1;
  wire [0:0] h_u_arrmul24_fa16_20_or0;
  wire [0:0] h_u_arrmul24_and17_20;
  wire [0:0] h_u_arrmul24_fa17_20_xor1;
  wire [0:0] h_u_arrmul24_fa17_20_or0;
  wire [0:0] h_u_arrmul24_and18_20;
  wire [0:0] h_u_arrmul24_fa18_20_xor1;
  wire [0:0] h_u_arrmul24_fa18_20_or0;
  wire [0:0] h_u_arrmul24_and19_20;
  wire [0:0] h_u_arrmul24_fa19_20_xor1;
  wire [0:0] h_u_arrmul24_fa19_20_or0;
  wire [0:0] h_u_arrmul24_and20_20;
  wire [0:0] h_u_arrmul24_fa20_20_xor1;
  wire [0:0] h_u_arrmul24_fa20_20_or0;
  wire [0:0] h_u_arrmul24_and21_20;
  wire [0:0] h_u_arrmul24_fa21_20_xor1;
  wire [0:0] h_u_arrmul24_fa21_20_or0;
  wire [0:0] h_u_arrmul24_and22_20;
  wire [0:0] h_u_arrmul24_fa22_20_xor1;
  wire [0:0] h_u_arrmul24_fa22_20_or0;
  wire [0:0] h_u_arrmul24_and23_20;
  wire [0:0] h_u_arrmul24_fa23_20_xor1;
  wire [0:0] h_u_arrmul24_fa23_20_or0;
  wire [0:0] h_u_arrmul24_and0_21;
  wire [0:0] h_u_arrmul24_ha0_21_xor0;
  wire [0:0] h_u_arrmul24_ha0_21_and0;
  wire [0:0] h_u_arrmul24_and1_21;
  wire [0:0] h_u_arrmul24_fa1_21_xor1;
  wire [0:0] h_u_arrmul24_fa1_21_or0;
  wire [0:0] h_u_arrmul24_and2_21;
  wire [0:0] h_u_arrmul24_fa2_21_xor1;
  wire [0:0] h_u_arrmul24_fa2_21_or0;
  wire [0:0] h_u_arrmul24_and3_21;
  wire [0:0] h_u_arrmul24_fa3_21_xor1;
  wire [0:0] h_u_arrmul24_fa3_21_or0;
  wire [0:0] h_u_arrmul24_and4_21;
  wire [0:0] h_u_arrmul24_fa4_21_xor1;
  wire [0:0] h_u_arrmul24_fa4_21_or0;
  wire [0:0] h_u_arrmul24_and5_21;
  wire [0:0] h_u_arrmul24_fa5_21_xor1;
  wire [0:0] h_u_arrmul24_fa5_21_or0;
  wire [0:0] h_u_arrmul24_and6_21;
  wire [0:0] h_u_arrmul24_fa6_21_xor1;
  wire [0:0] h_u_arrmul24_fa6_21_or0;
  wire [0:0] h_u_arrmul24_and7_21;
  wire [0:0] h_u_arrmul24_fa7_21_xor1;
  wire [0:0] h_u_arrmul24_fa7_21_or0;
  wire [0:0] h_u_arrmul24_and8_21;
  wire [0:0] h_u_arrmul24_fa8_21_xor1;
  wire [0:0] h_u_arrmul24_fa8_21_or0;
  wire [0:0] h_u_arrmul24_and9_21;
  wire [0:0] h_u_arrmul24_fa9_21_xor1;
  wire [0:0] h_u_arrmul24_fa9_21_or0;
  wire [0:0] h_u_arrmul24_and10_21;
  wire [0:0] h_u_arrmul24_fa10_21_xor1;
  wire [0:0] h_u_arrmul24_fa10_21_or0;
  wire [0:0] h_u_arrmul24_and11_21;
  wire [0:0] h_u_arrmul24_fa11_21_xor1;
  wire [0:0] h_u_arrmul24_fa11_21_or0;
  wire [0:0] h_u_arrmul24_and12_21;
  wire [0:0] h_u_arrmul24_fa12_21_xor1;
  wire [0:0] h_u_arrmul24_fa12_21_or0;
  wire [0:0] h_u_arrmul24_and13_21;
  wire [0:0] h_u_arrmul24_fa13_21_xor1;
  wire [0:0] h_u_arrmul24_fa13_21_or0;
  wire [0:0] h_u_arrmul24_and14_21;
  wire [0:0] h_u_arrmul24_fa14_21_xor1;
  wire [0:0] h_u_arrmul24_fa14_21_or0;
  wire [0:0] h_u_arrmul24_and15_21;
  wire [0:0] h_u_arrmul24_fa15_21_xor1;
  wire [0:0] h_u_arrmul24_fa15_21_or0;
  wire [0:0] h_u_arrmul24_and16_21;
  wire [0:0] h_u_arrmul24_fa16_21_xor1;
  wire [0:0] h_u_arrmul24_fa16_21_or0;
  wire [0:0] h_u_arrmul24_and17_21;
  wire [0:0] h_u_arrmul24_fa17_21_xor1;
  wire [0:0] h_u_arrmul24_fa17_21_or0;
  wire [0:0] h_u_arrmul24_and18_21;
  wire [0:0] h_u_arrmul24_fa18_21_xor1;
  wire [0:0] h_u_arrmul24_fa18_21_or0;
  wire [0:0] h_u_arrmul24_and19_21;
  wire [0:0] h_u_arrmul24_fa19_21_xor1;
  wire [0:0] h_u_arrmul24_fa19_21_or0;
  wire [0:0] h_u_arrmul24_and20_21;
  wire [0:0] h_u_arrmul24_fa20_21_xor1;
  wire [0:0] h_u_arrmul24_fa20_21_or0;
  wire [0:0] h_u_arrmul24_and21_21;
  wire [0:0] h_u_arrmul24_fa21_21_xor1;
  wire [0:0] h_u_arrmul24_fa21_21_or0;
  wire [0:0] h_u_arrmul24_and22_21;
  wire [0:0] h_u_arrmul24_fa22_21_xor1;
  wire [0:0] h_u_arrmul24_fa22_21_or0;
  wire [0:0] h_u_arrmul24_and23_21;
  wire [0:0] h_u_arrmul24_fa23_21_xor1;
  wire [0:0] h_u_arrmul24_fa23_21_or0;
  wire [0:0] h_u_arrmul24_and0_22;
  wire [0:0] h_u_arrmul24_ha0_22_xor0;
  wire [0:0] h_u_arrmul24_ha0_22_and0;
  wire [0:0] h_u_arrmul24_and1_22;
  wire [0:0] h_u_arrmul24_fa1_22_xor1;
  wire [0:0] h_u_arrmul24_fa1_22_or0;
  wire [0:0] h_u_arrmul24_and2_22;
  wire [0:0] h_u_arrmul24_fa2_22_xor1;
  wire [0:0] h_u_arrmul24_fa2_22_or0;
  wire [0:0] h_u_arrmul24_and3_22;
  wire [0:0] h_u_arrmul24_fa3_22_xor1;
  wire [0:0] h_u_arrmul24_fa3_22_or0;
  wire [0:0] h_u_arrmul24_and4_22;
  wire [0:0] h_u_arrmul24_fa4_22_xor1;
  wire [0:0] h_u_arrmul24_fa4_22_or0;
  wire [0:0] h_u_arrmul24_and5_22;
  wire [0:0] h_u_arrmul24_fa5_22_xor1;
  wire [0:0] h_u_arrmul24_fa5_22_or0;
  wire [0:0] h_u_arrmul24_and6_22;
  wire [0:0] h_u_arrmul24_fa6_22_xor1;
  wire [0:0] h_u_arrmul24_fa6_22_or0;
  wire [0:0] h_u_arrmul24_and7_22;
  wire [0:0] h_u_arrmul24_fa7_22_xor1;
  wire [0:0] h_u_arrmul24_fa7_22_or0;
  wire [0:0] h_u_arrmul24_and8_22;
  wire [0:0] h_u_arrmul24_fa8_22_xor1;
  wire [0:0] h_u_arrmul24_fa8_22_or0;
  wire [0:0] h_u_arrmul24_and9_22;
  wire [0:0] h_u_arrmul24_fa9_22_xor1;
  wire [0:0] h_u_arrmul24_fa9_22_or0;
  wire [0:0] h_u_arrmul24_and10_22;
  wire [0:0] h_u_arrmul24_fa10_22_xor1;
  wire [0:0] h_u_arrmul24_fa10_22_or0;
  wire [0:0] h_u_arrmul24_and11_22;
  wire [0:0] h_u_arrmul24_fa11_22_xor1;
  wire [0:0] h_u_arrmul24_fa11_22_or0;
  wire [0:0] h_u_arrmul24_and12_22;
  wire [0:0] h_u_arrmul24_fa12_22_xor1;
  wire [0:0] h_u_arrmul24_fa12_22_or0;
  wire [0:0] h_u_arrmul24_and13_22;
  wire [0:0] h_u_arrmul24_fa13_22_xor1;
  wire [0:0] h_u_arrmul24_fa13_22_or0;
  wire [0:0] h_u_arrmul24_and14_22;
  wire [0:0] h_u_arrmul24_fa14_22_xor1;
  wire [0:0] h_u_arrmul24_fa14_22_or0;
  wire [0:0] h_u_arrmul24_and15_22;
  wire [0:0] h_u_arrmul24_fa15_22_xor1;
  wire [0:0] h_u_arrmul24_fa15_22_or0;
  wire [0:0] h_u_arrmul24_and16_22;
  wire [0:0] h_u_arrmul24_fa16_22_xor1;
  wire [0:0] h_u_arrmul24_fa16_22_or0;
  wire [0:0] h_u_arrmul24_and17_22;
  wire [0:0] h_u_arrmul24_fa17_22_xor1;
  wire [0:0] h_u_arrmul24_fa17_22_or0;
  wire [0:0] h_u_arrmul24_and18_22;
  wire [0:0] h_u_arrmul24_fa18_22_xor1;
  wire [0:0] h_u_arrmul24_fa18_22_or0;
  wire [0:0] h_u_arrmul24_and19_22;
  wire [0:0] h_u_arrmul24_fa19_22_xor1;
  wire [0:0] h_u_arrmul24_fa19_22_or0;
  wire [0:0] h_u_arrmul24_and20_22;
  wire [0:0] h_u_arrmul24_fa20_22_xor1;
  wire [0:0] h_u_arrmul24_fa20_22_or0;
  wire [0:0] h_u_arrmul24_and21_22;
  wire [0:0] h_u_arrmul24_fa21_22_xor1;
  wire [0:0] h_u_arrmul24_fa21_22_or0;
  wire [0:0] h_u_arrmul24_and22_22;
  wire [0:0] h_u_arrmul24_fa22_22_xor1;
  wire [0:0] h_u_arrmul24_fa22_22_or0;
  wire [0:0] h_u_arrmul24_and23_22;
  wire [0:0] h_u_arrmul24_fa23_22_xor1;
  wire [0:0] h_u_arrmul24_fa23_22_or0;
  wire [0:0] h_u_arrmul24_and0_23;
  wire [0:0] h_u_arrmul24_ha0_23_xor0;
  wire [0:0] h_u_arrmul24_ha0_23_and0;
  wire [0:0] h_u_arrmul24_and1_23;
  wire [0:0] h_u_arrmul24_fa1_23_xor1;
  wire [0:0] h_u_arrmul24_fa1_23_or0;
  wire [0:0] h_u_arrmul24_and2_23;
  wire [0:0] h_u_arrmul24_fa2_23_xor1;
  wire [0:0] h_u_arrmul24_fa2_23_or0;
  wire [0:0] h_u_arrmul24_and3_23;
  wire [0:0] h_u_arrmul24_fa3_23_xor1;
  wire [0:0] h_u_arrmul24_fa3_23_or0;
  wire [0:0] h_u_arrmul24_and4_23;
  wire [0:0] h_u_arrmul24_fa4_23_xor1;
  wire [0:0] h_u_arrmul24_fa4_23_or0;
  wire [0:0] h_u_arrmul24_and5_23;
  wire [0:0] h_u_arrmul24_fa5_23_xor1;
  wire [0:0] h_u_arrmul24_fa5_23_or0;
  wire [0:0] h_u_arrmul24_and6_23;
  wire [0:0] h_u_arrmul24_fa6_23_xor1;
  wire [0:0] h_u_arrmul24_fa6_23_or0;
  wire [0:0] h_u_arrmul24_and7_23;
  wire [0:0] h_u_arrmul24_fa7_23_xor1;
  wire [0:0] h_u_arrmul24_fa7_23_or0;
  wire [0:0] h_u_arrmul24_and8_23;
  wire [0:0] h_u_arrmul24_fa8_23_xor1;
  wire [0:0] h_u_arrmul24_fa8_23_or0;
  wire [0:0] h_u_arrmul24_and9_23;
  wire [0:0] h_u_arrmul24_fa9_23_xor1;
  wire [0:0] h_u_arrmul24_fa9_23_or0;
  wire [0:0] h_u_arrmul24_and10_23;
  wire [0:0] h_u_arrmul24_fa10_23_xor1;
  wire [0:0] h_u_arrmul24_fa10_23_or0;
  wire [0:0] h_u_arrmul24_and11_23;
  wire [0:0] h_u_arrmul24_fa11_23_xor1;
  wire [0:0] h_u_arrmul24_fa11_23_or0;
  wire [0:0] h_u_arrmul24_and12_23;
  wire [0:0] h_u_arrmul24_fa12_23_xor1;
  wire [0:0] h_u_arrmul24_fa12_23_or0;
  wire [0:0] h_u_arrmul24_and13_23;
  wire [0:0] h_u_arrmul24_fa13_23_xor1;
  wire [0:0] h_u_arrmul24_fa13_23_or0;
  wire [0:0] h_u_arrmul24_and14_23;
  wire [0:0] h_u_arrmul24_fa14_23_xor1;
  wire [0:0] h_u_arrmul24_fa14_23_or0;
  wire [0:0] h_u_arrmul24_and15_23;
  wire [0:0] h_u_arrmul24_fa15_23_xor1;
  wire [0:0] h_u_arrmul24_fa15_23_or0;
  wire [0:0] h_u_arrmul24_and16_23;
  wire [0:0] h_u_arrmul24_fa16_23_xor1;
  wire [0:0] h_u_arrmul24_fa16_23_or0;
  wire [0:0] h_u_arrmul24_and17_23;
  wire [0:0] h_u_arrmul24_fa17_23_xor1;
  wire [0:0] h_u_arrmul24_fa17_23_or0;
  wire [0:0] h_u_arrmul24_and18_23;
  wire [0:0] h_u_arrmul24_fa18_23_xor1;
  wire [0:0] h_u_arrmul24_fa18_23_or0;
  wire [0:0] h_u_arrmul24_and19_23;
  wire [0:0] h_u_arrmul24_fa19_23_xor1;
  wire [0:0] h_u_arrmul24_fa19_23_or0;
  wire [0:0] h_u_arrmul24_and20_23;
  wire [0:0] h_u_arrmul24_fa20_23_xor1;
  wire [0:0] h_u_arrmul24_fa20_23_or0;
  wire [0:0] h_u_arrmul24_and21_23;
  wire [0:0] h_u_arrmul24_fa21_23_xor1;
  wire [0:0] h_u_arrmul24_fa21_23_or0;
  wire [0:0] h_u_arrmul24_and22_23;
  wire [0:0] h_u_arrmul24_fa22_23_xor1;
  wire [0:0] h_u_arrmul24_fa22_23_or0;
  wire [0:0] h_u_arrmul24_and23_23;
  wire [0:0] h_u_arrmul24_fa23_23_xor1;
  wire [0:0] h_u_arrmul24_fa23_23_or0;

  and_gate and_gate_h_u_arrmul24_and0_0(a[0], b[0], h_u_arrmul24_and0_0);
  and_gate and_gate_h_u_arrmul24_and1_0(a[1], b[0], h_u_arrmul24_and1_0);
  and_gate and_gate_h_u_arrmul24_and2_0(a[2], b[0], h_u_arrmul24_and2_0);
  and_gate and_gate_h_u_arrmul24_and3_0(a[3], b[0], h_u_arrmul24_and3_0);
  and_gate and_gate_h_u_arrmul24_and4_0(a[4], b[0], h_u_arrmul24_and4_0);
  and_gate and_gate_h_u_arrmul24_and5_0(a[5], b[0], h_u_arrmul24_and5_0);
  and_gate and_gate_h_u_arrmul24_and6_0(a[6], b[0], h_u_arrmul24_and6_0);
  and_gate and_gate_h_u_arrmul24_and7_0(a[7], b[0], h_u_arrmul24_and7_0);
  and_gate and_gate_h_u_arrmul24_and8_0(a[8], b[0], h_u_arrmul24_and8_0);
  and_gate and_gate_h_u_arrmul24_and9_0(a[9], b[0], h_u_arrmul24_and9_0);
  and_gate and_gate_h_u_arrmul24_and10_0(a[10], b[0], h_u_arrmul24_and10_0);
  and_gate and_gate_h_u_arrmul24_and11_0(a[11], b[0], h_u_arrmul24_and11_0);
  and_gate and_gate_h_u_arrmul24_and12_0(a[12], b[0], h_u_arrmul24_and12_0);
  and_gate and_gate_h_u_arrmul24_and13_0(a[13], b[0], h_u_arrmul24_and13_0);
  and_gate and_gate_h_u_arrmul24_and14_0(a[14], b[0], h_u_arrmul24_and14_0);
  and_gate and_gate_h_u_arrmul24_and15_0(a[15], b[0], h_u_arrmul24_and15_0);
  and_gate and_gate_h_u_arrmul24_and16_0(a[16], b[0], h_u_arrmul24_and16_0);
  and_gate and_gate_h_u_arrmul24_and17_0(a[17], b[0], h_u_arrmul24_and17_0);
  and_gate and_gate_h_u_arrmul24_and18_0(a[18], b[0], h_u_arrmul24_and18_0);
  and_gate and_gate_h_u_arrmul24_and19_0(a[19], b[0], h_u_arrmul24_and19_0);
  and_gate and_gate_h_u_arrmul24_and20_0(a[20], b[0], h_u_arrmul24_and20_0);
  and_gate and_gate_h_u_arrmul24_and21_0(a[21], b[0], h_u_arrmul24_and21_0);
  and_gate and_gate_h_u_arrmul24_and22_0(a[22], b[0], h_u_arrmul24_and22_0);
  and_gate and_gate_h_u_arrmul24_and23_0(a[23], b[0], h_u_arrmul24_and23_0);
  and_gate and_gate_h_u_arrmul24_and0_1(a[0], b[1], h_u_arrmul24_and0_1);
  ha ha_h_u_arrmul24_ha0_1_out(h_u_arrmul24_and0_1[0], h_u_arrmul24_and1_0[0], h_u_arrmul24_ha0_1_xor0, h_u_arrmul24_ha0_1_and0);
  and_gate and_gate_h_u_arrmul24_and1_1(a[1], b[1], h_u_arrmul24_and1_1);
  fa fa_h_u_arrmul24_fa1_1_out(h_u_arrmul24_and1_1[0], h_u_arrmul24_and2_0[0], h_u_arrmul24_ha0_1_and0[0], h_u_arrmul24_fa1_1_xor1, h_u_arrmul24_fa1_1_or0);
  and_gate and_gate_h_u_arrmul24_and2_1(a[2], b[1], h_u_arrmul24_and2_1);
  fa fa_h_u_arrmul24_fa2_1_out(h_u_arrmul24_and2_1[0], h_u_arrmul24_and3_0[0], h_u_arrmul24_fa1_1_or0[0], h_u_arrmul24_fa2_1_xor1, h_u_arrmul24_fa2_1_or0);
  and_gate and_gate_h_u_arrmul24_and3_1(a[3], b[1], h_u_arrmul24_and3_1);
  fa fa_h_u_arrmul24_fa3_1_out(h_u_arrmul24_and3_1[0], h_u_arrmul24_and4_0[0], h_u_arrmul24_fa2_1_or0[0], h_u_arrmul24_fa3_1_xor1, h_u_arrmul24_fa3_1_or0);
  and_gate and_gate_h_u_arrmul24_and4_1(a[4], b[1], h_u_arrmul24_and4_1);
  fa fa_h_u_arrmul24_fa4_1_out(h_u_arrmul24_and4_1[0], h_u_arrmul24_and5_0[0], h_u_arrmul24_fa3_1_or0[0], h_u_arrmul24_fa4_1_xor1, h_u_arrmul24_fa4_1_or0);
  and_gate and_gate_h_u_arrmul24_and5_1(a[5], b[1], h_u_arrmul24_and5_1);
  fa fa_h_u_arrmul24_fa5_1_out(h_u_arrmul24_and5_1[0], h_u_arrmul24_and6_0[0], h_u_arrmul24_fa4_1_or0[0], h_u_arrmul24_fa5_1_xor1, h_u_arrmul24_fa5_1_or0);
  and_gate and_gate_h_u_arrmul24_and6_1(a[6], b[1], h_u_arrmul24_and6_1);
  fa fa_h_u_arrmul24_fa6_1_out(h_u_arrmul24_and6_1[0], h_u_arrmul24_and7_0[0], h_u_arrmul24_fa5_1_or0[0], h_u_arrmul24_fa6_1_xor1, h_u_arrmul24_fa6_1_or0);
  and_gate and_gate_h_u_arrmul24_and7_1(a[7], b[1], h_u_arrmul24_and7_1);
  fa fa_h_u_arrmul24_fa7_1_out(h_u_arrmul24_and7_1[0], h_u_arrmul24_and8_0[0], h_u_arrmul24_fa6_1_or0[0], h_u_arrmul24_fa7_1_xor1, h_u_arrmul24_fa7_1_or0);
  and_gate and_gate_h_u_arrmul24_and8_1(a[8], b[1], h_u_arrmul24_and8_1);
  fa fa_h_u_arrmul24_fa8_1_out(h_u_arrmul24_and8_1[0], h_u_arrmul24_and9_0[0], h_u_arrmul24_fa7_1_or0[0], h_u_arrmul24_fa8_1_xor1, h_u_arrmul24_fa8_1_or0);
  and_gate and_gate_h_u_arrmul24_and9_1(a[9], b[1], h_u_arrmul24_and9_1);
  fa fa_h_u_arrmul24_fa9_1_out(h_u_arrmul24_and9_1[0], h_u_arrmul24_and10_0[0], h_u_arrmul24_fa8_1_or0[0], h_u_arrmul24_fa9_1_xor1, h_u_arrmul24_fa9_1_or0);
  and_gate and_gate_h_u_arrmul24_and10_1(a[10], b[1], h_u_arrmul24_and10_1);
  fa fa_h_u_arrmul24_fa10_1_out(h_u_arrmul24_and10_1[0], h_u_arrmul24_and11_0[0], h_u_arrmul24_fa9_1_or0[0], h_u_arrmul24_fa10_1_xor1, h_u_arrmul24_fa10_1_or0);
  and_gate and_gate_h_u_arrmul24_and11_1(a[11], b[1], h_u_arrmul24_and11_1);
  fa fa_h_u_arrmul24_fa11_1_out(h_u_arrmul24_and11_1[0], h_u_arrmul24_and12_0[0], h_u_arrmul24_fa10_1_or0[0], h_u_arrmul24_fa11_1_xor1, h_u_arrmul24_fa11_1_or0);
  and_gate and_gate_h_u_arrmul24_and12_1(a[12], b[1], h_u_arrmul24_and12_1);
  fa fa_h_u_arrmul24_fa12_1_out(h_u_arrmul24_and12_1[0], h_u_arrmul24_and13_0[0], h_u_arrmul24_fa11_1_or0[0], h_u_arrmul24_fa12_1_xor1, h_u_arrmul24_fa12_1_or0);
  and_gate and_gate_h_u_arrmul24_and13_1(a[13], b[1], h_u_arrmul24_and13_1);
  fa fa_h_u_arrmul24_fa13_1_out(h_u_arrmul24_and13_1[0], h_u_arrmul24_and14_0[0], h_u_arrmul24_fa12_1_or0[0], h_u_arrmul24_fa13_1_xor1, h_u_arrmul24_fa13_1_or0);
  and_gate and_gate_h_u_arrmul24_and14_1(a[14], b[1], h_u_arrmul24_and14_1);
  fa fa_h_u_arrmul24_fa14_1_out(h_u_arrmul24_and14_1[0], h_u_arrmul24_and15_0[0], h_u_arrmul24_fa13_1_or0[0], h_u_arrmul24_fa14_1_xor1, h_u_arrmul24_fa14_1_or0);
  and_gate and_gate_h_u_arrmul24_and15_1(a[15], b[1], h_u_arrmul24_and15_1);
  fa fa_h_u_arrmul24_fa15_1_out(h_u_arrmul24_and15_1[0], h_u_arrmul24_and16_0[0], h_u_arrmul24_fa14_1_or0[0], h_u_arrmul24_fa15_1_xor1, h_u_arrmul24_fa15_1_or0);
  and_gate and_gate_h_u_arrmul24_and16_1(a[16], b[1], h_u_arrmul24_and16_1);
  fa fa_h_u_arrmul24_fa16_1_out(h_u_arrmul24_and16_1[0], h_u_arrmul24_and17_0[0], h_u_arrmul24_fa15_1_or0[0], h_u_arrmul24_fa16_1_xor1, h_u_arrmul24_fa16_1_or0);
  and_gate and_gate_h_u_arrmul24_and17_1(a[17], b[1], h_u_arrmul24_and17_1);
  fa fa_h_u_arrmul24_fa17_1_out(h_u_arrmul24_and17_1[0], h_u_arrmul24_and18_0[0], h_u_arrmul24_fa16_1_or0[0], h_u_arrmul24_fa17_1_xor1, h_u_arrmul24_fa17_1_or0);
  and_gate and_gate_h_u_arrmul24_and18_1(a[18], b[1], h_u_arrmul24_and18_1);
  fa fa_h_u_arrmul24_fa18_1_out(h_u_arrmul24_and18_1[0], h_u_arrmul24_and19_0[0], h_u_arrmul24_fa17_1_or0[0], h_u_arrmul24_fa18_1_xor1, h_u_arrmul24_fa18_1_or0);
  and_gate and_gate_h_u_arrmul24_and19_1(a[19], b[1], h_u_arrmul24_and19_1);
  fa fa_h_u_arrmul24_fa19_1_out(h_u_arrmul24_and19_1[0], h_u_arrmul24_and20_0[0], h_u_arrmul24_fa18_1_or0[0], h_u_arrmul24_fa19_1_xor1, h_u_arrmul24_fa19_1_or0);
  and_gate and_gate_h_u_arrmul24_and20_1(a[20], b[1], h_u_arrmul24_and20_1);
  fa fa_h_u_arrmul24_fa20_1_out(h_u_arrmul24_and20_1[0], h_u_arrmul24_and21_0[0], h_u_arrmul24_fa19_1_or0[0], h_u_arrmul24_fa20_1_xor1, h_u_arrmul24_fa20_1_or0);
  and_gate and_gate_h_u_arrmul24_and21_1(a[21], b[1], h_u_arrmul24_and21_1);
  fa fa_h_u_arrmul24_fa21_1_out(h_u_arrmul24_and21_1[0], h_u_arrmul24_and22_0[0], h_u_arrmul24_fa20_1_or0[0], h_u_arrmul24_fa21_1_xor1, h_u_arrmul24_fa21_1_or0);
  and_gate and_gate_h_u_arrmul24_and22_1(a[22], b[1], h_u_arrmul24_and22_1);
  fa fa_h_u_arrmul24_fa22_1_out(h_u_arrmul24_and22_1[0], h_u_arrmul24_and23_0[0], h_u_arrmul24_fa21_1_or0[0], h_u_arrmul24_fa22_1_xor1, h_u_arrmul24_fa22_1_or0);
  and_gate and_gate_h_u_arrmul24_and23_1(a[23], b[1], h_u_arrmul24_and23_1);
  ha ha_h_u_arrmul24_ha23_1_out(h_u_arrmul24_and23_1[0], h_u_arrmul24_fa22_1_or0[0], h_u_arrmul24_ha23_1_xor0, h_u_arrmul24_ha23_1_and0);
  and_gate and_gate_h_u_arrmul24_and0_2(a[0], b[2], h_u_arrmul24_and0_2);
  ha ha_h_u_arrmul24_ha0_2_out(h_u_arrmul24_and0_2[0], h_u_arrmul24_fa1_1_xor1[0], h_u_arrmul24_ha0_2_xor0, h_u_arrmul24_ha0_2_and0);
  and_gate and_gate_h_u_arrmul24_and1_2(a[1], b[2], h_u_arrmul24_and1_2);
  fa fa_h_u_arrmul24_fa1_2_out(h_u_arrmul24_and1_2[0], h_u_arrmul24_fa2_1_xor1[0], h_u_arrmul24_ha0_2_and0[0], h_u_arrmul24_fa1_2_xor1, h_u_arrmul24_fa1_2_or0);
  and_gate and_gate_h_u_arrmul24_and2_2(a[2], b[2], h_u_arrmul24_and2_2);
  fa fa_h_u_arrmul24_fa2_2_out(h_u_arrmul24_and2_2[0], h_u_arrmul24_fa3_1_xor1[0], h_u_arrmul24_fa1_2_or0[0], h_u_arrmul24_fa2_2_xor1, h_u_arrmul24_fa2_2_or0);
  and_gate and_gate_h_u_arrmul24_and3_2(a[3], b[2], h_u_arrmul24_and3_2);
  fa fa_h_u_arrmul24_fa3_2_out(h_u_arrmul24_and3_2[0], h_u_arrmul24_fa4_1_xor1[0], h_u_arrmul24_fa2_2_or0[0], h_u_arrmul24_fa3_2_xor1, h_u_arrmul24_fa3_2_or0);
  and_gate and_gate_h_u_arrmul24_and4_2(a[4], b[2], h_u_arrmul24_and4_2);
  fa fa_h_u_arrmul24_fa4_2_out(h_u_arrmul24_and4_2[0], h_u_arrmul24_fa5_1_xor1[0], h_u_arrmul24_fa3_2_or0[0], h_u_arrmul24_fa4_2_xor1, h_u_arrmul24_fa4_2_or0);
  and_gate and_gate_h_u_arrmul24_and5_2(a[5], b[2], h_u_arrmul24_and5_2);
  fa fa_h_u_arrmul24_fa5_2_out(h_u_arrmul24_and5_2[0], h_u_arrmul24_fa6_1_xor1[0], h_u_arrmul24_fa4_2_or0[0], h_u_arrmul24_fa5_2_xor1, h_u_arrmul24_fa5_2_or0);
  and_gate and_gate_h_u_arrmul24_and6_2(a[6], b[2], h_u_arrmul24_and6_2);
  fa fa_h_u_arrmul24_fa6_2_out(h_u_arrmul24_and6_2[0], h_u_arrmul24_fa7_1_xor1[0], h_u_arrmul24_fa5_2_or0[0], h_u_arrmul24_fa6_2_xor1, h_u_arrmul24_fa6_2_or0);
  and_gate and_gate_h_u_arrmul24_and7_2(a[7], b[2], h_u_arrmul24_and7_2);
  fa fa_h_u_arrmul24_fa7_2_out(h_u_arrmul24_and7_2[0], h_u_arrmul24_fa8_1_xor1[0], h_u_arrmul24_fa6_2_or0[0], h_u_arrmul24_fa7_2_xor1, h_u_arrmul24_fa7_2_or0);
  and_gate and_gate_h_u_arrmul24_and8_2(a[8], b[2], h_u_arrmul24_and8_2);
  fa fa_h_u_arrmul24_fa8_2_out(h_u_arrmul24_and8_2[0], h_u_arrmul24_fa9_1_xor1[0], h_u_arrmul24_fa7_2_or0[0], h_u_arrmul24_fa8_2_xor1, h_u_arrmul24_fa8_2_or0);
  and_gate and_gate_h_u_arrmul24_and9_2(a[9], b[2], h_u_arrmul24_and9_2);
  fa fa_h_u_arrmul24_fa9_2_out(h_u_arrmul24_and9_2[0], h_u_arrmul24_fa10_1_xor1[0], h_u_arrmul24_fa8_2_or0[0], h_u_arrmul24_fa9_2_xor1, h_u_arrmul24_fa9_2_or0);
  and_gate and_gate_h_u_arrmul24_and10_2(a[10], b[2], h_u_arrmul24_and10_2);
  fa fa_h_u_arrmul24_fa10_2_out(h_u_arrmul24_and10_2[0], h_u_arrmul24_fa11_1_xor1[0], h_u_arrmul24_fa9_2_or0[0], h_u_arrmul24_fa10_2_xor1, h_u_arrmul24_fa10_2_or0);
  and_gate and_gate_h_u_arrmul24_and11_2(a[11], b[2], h_u_arrmul24_and11_2);
  fa fa_h_u_arrmul24_fa11_2_out(h_u_arrmul24_and11_2[0], h_u_arrmul24_fa12_1_xor1[0], h_u_arrmul24_fa10_2_or0[0], h_u_arrmul24_fa11_2_xor1, h_u_arrmul24_fa11_2_or0);
  and_gate and_gate_h_u_arrmul24_and12_2(a[12], b[2], h_u_arrmul24_and12_2);
  fa fa_h_u_arrmul24_fa12_2_out(h_u_arrmul24_and12_2[0], h_u_arrmul24_fa13_1_xor1[0], h_u_arrmul24_fa11_2_or0[0], h_u_arrmul24_fa12_2_xor1, h_u_arrmul24_fa12_2_or0);
  and_gate and_gate_h_u_arrmul24_and13_2(a[13], b[2], h_u_arrmul24_and13_2);
  fa fa_h_u_arrmul24_fa13_2_out(h_u_arrmul24_and13_2[0], h_u_arrmul24_fa14_1_xor1[0], h_u_arrmul24_fa12_2_or0[0], h_u_arrmul24_fa13_2_xor1, h_u_arrmul24_fa13_2_or0);
  and_gate and_gate_h_u_arrmul24_and14_2(a[14], b[2], h_u_arrmul24_and14_2);
  fa fa_h_u_arrmul24_fa14_2_out(h_u_arrmul24_and14_2[0], h_u_arrmul24_fa15_1_xor1[0], h_u_arrmul24_fa13_2_or0[0], h_u_arrmul24_fa14_2_xor1, h_u_arrmul24_fa14_2_or0);
  and_gate and_gate_h_u_arrmul24_and15_2(a[15], b[2], h_u_arrmul24_and15_2);
  fa fa_h_u_arrmul24_fa15_2_out(h_u_arrmul24_and15_2[0], h_u_arrmul24_fa16_1_xor1[0], h_u_arrmul24_fa14_2_or0[0], h_u_arrmul24_fa15_2_xor1, h_u_arrmul24_fa15_2_or0);
  and_gate and_gate_h_u_arrmul24_and16_2(a[16], b[2], h_u_arrmul24_and16_2);
  fa fa_h_u_arrmul24_fa16_2_out(h_u_arrmul24_and16_2[0], h_u_arrmul24_fa17_1_xor1[0], h_u_arrmul24_fa15_2_or0[0], h_u_arrmul24_fa16_2_xor1, h_u_arrmul24_fa16_2_or0);
  and_gate and_gate_h_u_arrmul24_and17_2(a[17], b[2], h_u_arrmul24_and17_2);
  fa fa_h_u_arrmul24_fa17_2_out(h_u_arrmul24_and17_2[0], h_u_arrmul24_fa18_1_xor1[0], h_u_arrmul24_fa16_2_or0[0], h_u_arrmul24_fa17_2_xor1, h_u_arrmul24_fa17_2_or0);
  and_gate and_gate_h_u_arrmul24_and18_2(a[18], b[2], h_u_arrmul24_and18_2);
  fa fa_h_u_arrmul24_fa18_2_out(h_u_arrmul24_and18_2[0], h_u_arrmul24_fa19_1_xor1[0], h_u_arrmul24_fa17_2_or0[0], h_u_arrmul24_fa18_2_xor1, h_u_arrmul24_fa18_2_or0);
  and_gate and_gate_h_u_arrmul24_and19_2(a[19], b[2], h_u_arrmul24_and19_2);
  fa fa_h_u_arrmul24_fa19_2_out(h_u_arrmul24_and19_2[0], h_u_arrmul24_fa20_1_xor1[0], h_u_arrmul24_fa18_2_or0[0], h_u_arrmul24_fa19_2_xor1, h_u_arrmul24_fa19_2_or0);
  and_gate and_gate_h_u_arrmul24_and20_2(a[20], b[2], h_u_arrmul24_and20_2);
  fa fa_h_u_arrmul24_fa20_2_out(h_u_arrmul24_and20_2[0], h_u_arrmul24_fa21_1_xor1[0], h_u_arrmul24_fa19_2_or0[0], h_u_arrmul24_fa20_2_xor1, h_u_arrmul24_fa20_2_or0);
  and_gate and_gate_h_u_arrmul24_and21_2(a[21], b[2], h_u_arrmul24_and21_2);
  fa fa_h_u_arrmul24_fa21_2_out(h_u_arrmul24_and21_2[0], h_u_arrmul24_fa22_1_xor1[0], h_u_arrmul24_fa20_2_or0[0], h_u_arrmul24_fa21_2_xor1, h_u_arrmul24_fa21_2_or0);
  and_gate and_gate_h_u_arrmul24_and22_2(a[22], b[2], h_u_arrmul24_and22_2);
  fa fa_h_u_arrmul24_fa22_2_out(h_u_arrmul24_and22_2[0], h_u_arrmul24_ha23_1_xor0[0], h_u_arrmul24_fa21_2_or0[0], h_u_arrmul24_fa22_2_xor1, h_u_arrmul24_fa22_2_or0);
  and_gate and_gate_h_u_arrmul24_and23_2(a[23], b[2], h_u_arrmul24_and23_2);
  fa fa_h_u_arrmul24_fa23_2_out(h_u_arrmul24_and23_2[0], h_u_arrmul24_ha23_1_and0[0], h_u_arrmul24_fa22_2_or0[0], h_u_arrmul24_fa23_2_xor1, h_u_arrmul24_fa23_2_or0);
  and_gate and_gate_h_u_arrmul24_and0_3(a[0], b[3], h_u_arrmul24_and0_3);
  ha ha_h_u_arrmul24_ha0_3_out(h_u_arrmul24_and0_3[0], h_u_arrmul24_fa1_2_xor1[0], h_u_arrmul24_ha0_3_xor0, h_u_arrmul24_ha0_3_and0);
  and_gate and_gate_h_u_arrmul24_and1_3(a[1], b[3], h_u_arrmul24_and1_3);
  fa fa_h_u_arrmul24_fa1_3_out(h_u_arrmul24_and1_3[0], h_u_arrmul24_fa2_2_xor1[0], h_u_arrmul24_ha0_3_and0[0], h_u_arrmul24_fa1_3_xor1, h_u_arrmul24_fa1_3_or0);
  and_gate and_gate_h_u_arrmul24_and2_3(a[2], b[3], h_u_arrmul24_and2_3);
  fa fa_h_u_arrmul24_fa2_3_out(h_u_arrmul24_and2_3[0], h_u_arrmul24_fa3_2_xor1[0], h_u_arrmul24_fa1_3_or0[0], h_u_arrmul24_fa2_3_xor1, h_u_arrmul24_fa2_3_or0);
  and_gate and_gate_h_u_arrmul24_and3_3(a[3], b[3], h_u_arrmul24_and3_3);
  fa fa_h_u_arrmul24_fa3_3_out(h_u_arrmul24_and3_3[0], h_u_arrmul24_fa4_2_xor1[0], h_u_arrmul24_fa2_3_or0[0], h_u_arrmul24_fa3_3_xor1, h_u_arrmul24_fa3_3_or0);
  and_gate and_gate_h_u_arrmul24_and4_3(a[4], b[3], h_u_arrmul24_and4_3);
  fa fa_h_u_arrmul24_fa4_3_out(h_u_arrmul24_and4_3[0], h_u_arrmul24_fa5_2_xor1[0], h_u_arrmul24_fa3_3_or0[0], h_u_arrmul24_fa4_3_xor1, h_u_arrmul24_fa4_3_or0);
  and_gate and_gate_h_u_arrmul24_and5_3(a[5], b[3], h_u_arrmul24_and5_3);
  fa fa_h_u_arrmul24_fa5_3_out(h_u_arrmul24_and5_3[0], h_u_arrmul24_fa6_2_xor1[0], h_u_arrmul24_fa4_3_or0[0], h_u_arrmul24_fa5_3_xor1, h_u_arrmul24_fa5_3_or0);
  and_gate and_gate_h_u_arrmul24_and6_3(a[6], b[3], h_u_arrmul24_and6_3);
  fa fa_h_u_arrmul24_fa6_3_out(h_u_arrmul24_and6_3[0], h_u_arrmul24_fa7_2_xor1[0], h_u_arrmul24_fa5_3_or0[0], h_u_arrmul24_fa6_3_xor1, h_u_arrmul24_fa6_3_or0);
  and_gate and_gate_h_u_arrmul24_and7_3(a[7], b[3], h_u_arrmul24_and7_3);
  fa fa_h_u_arrmul24_fa7_3_out(h_u_arrmul24_and7_3[0], h_u_arrmul24_fa8_2_xor1[0], h_u_arrmul24_fa6_3_or0[0], h_u_arrmul24_fa7_3_xor1, h_u_arrmul24_fa7_3_or0);
  and_gate and_gate_h_u_arrmul24_and8_3(a[8], b[3], h_u_arrmul24_and8_3);
  fa fa_h_u_arrmul24_fa8_3_out(h_u_arrmul24_and8_3[0], h_u_arrmul24_fa9_2_xor1[0], h_u_arrmul24_fa7_3_or0[0], h_u_arrmul24_fa8_3_xor1, h_u_arrmul24_fa8_3_or0);
  and_gate and_gate_h_u_arrmul24_and9_3(a[9], b[3], h_u_arrmul24_and9_3);
  fa fa_h_u_arrmul24_fa9_3_out(h_u_arrmul24_and9_3[0], h_u_arrmul24_fa10_2_xor1[0], h_u_arrmul24_fa8_3_or0[0], h_u_arrmul24_fa9_3_xor1, h_u_arrmul24_fa9_3_or0);
  and_gate and_gate_h_u_arrmul24_and10_3(a[10], b[3], h_u_arrmul24_and10_3);
  fa fa_h_u_arrmul24_fa10_3_out(h_u_arrmul24_and10_3[0], h_u_arrmul24_fa11_2_xor1[0], h_u_arrmul24_fa9_3_or0[0], h_u_arrmul24_fa10_3_xor1, h_u_arrmul24_fa10_3_or0);
  and_gate and_gate_h_u_arrmul24_and11_3(a[11], b[3], h_u_arrmul24_and11_3);
  fa fa_h_u_arrmul24_fa11_3_out(h_u_arrmul24_and11_3[0], h_u_arrmul24_fa12_2_xor1[0], h_u_arrmul24_fa10_3_or0[0], h_u_arrmul24_fa11_3_xor1, h_u_arrmul24_fa11_3_or0);
  and_gate and_gate_h_u_arrmul24_and12_3(a[12], b[3], h_u_arrmul24_and12_3);
  fa fa_h_u_arrmul24_fa12_3_out(h_u_arrmul24_and12_3[0], h_u_arrmul24_fa13_2_xor1[0], h_u_arrmul24_fa11_3_or0[0], h_u_arrmul24_fa12_3_xor1, h_u_arrmul24_fa12_3_or0);
  and_gate and_gate_h_u_arrmul24_and13_3(a[13], b[3], h_u_arrmul24_and13_3);
  fa fa_h_u_arrmul24_fa13_3_out(h_u_arrmul24_and13_3[0], h_u_arrmul24_fa14_2_xor1[0], h_u_arrmul24_fa12_3_or0[0], h_u_arrmul24_fa13_3_xor1, h_u_arrmul24_fa13_3_or0);
  and_gate and_gate_h_u_arrmul24_and14_3(a[14], b[3], h_u_arrmul24_and14_3);
  fa fa_h_u_arrmul24_fa14_3_out(h_u_arrmul24_and14_3[0], h_u_arrmul24_fa15_2_xor1[0], h_u_arrmul24_fa13_3_or0[0], h_u_arrmul24_fa14_3_xor1, h_u_arrmul24_fa14_3_or0);
  and_gate and_gate_h_u_arrmul24_and15_3(a[15], b[3], h_u_arrmul24_and15_3);
  fa fa_h_u_arrmul24_fa15_3_out(h_u_arrmul24_and15_3[0], h_u_arrmul24_fa16_2_xor1[0], h_u_arrmul24_fa14_3_or0[0], h_u_arrmul24_fa15_3_xor1, h_u_arrmul24_fa15_3_or0);
  and_gate and_gate_h_u_arrmul24_and16_3(a[16], b[3], h_u_arrmul24_and16_3);
  fa fa_h_u_arrmul24_fa16_3_out(h_u_arrmul24_and16_3[0], h_u_arrmul24_fa17_2_xor1[0], h_u_arrmul24_fa15_3_or0[0], h_u_arrmul24_fa16_3_xor1, h_u_arrmul24_fa16_3_or0);
  and_gate and_gate_h_u_arrmul24_and17_3(a[17], b[3], h_u_arrmul24_and17_3);
  fa fa_h_u_arrmul24_fa17_3_out(h_u_arrmul24_and17_3[0], h_u_arrmul24_fa18_2_xor1[0], h_u_arrmul24_fa16_3_or0[0], h_u_arrmul24_fa17_3_xor1, h_u_arrmul24_fa17_3_or0);
  and_gate and_gate_h_u_arrmul24_and18_3(a[18], b[3], h_u_arrmul24_and18_3);
  fa fa_h_u_arrmul24_fa18_3_out(h_u_arrmul24_and18_3[0], h_u_arrmul24_fa19_2_xor1[0], h_u_arrmul24_fa17_3_or0[0], h_u_arrmul24_fa18_3_xor1, h_u_arrmul24_fa18_3_or0);
  and_gate and_gate_h_u_arrmul24_and19_3(a[19], b[3], h_u_arrmul24_and19_3);
  fa fa_h_u_arrmul24_fa19_3_out(h_u_arrmul24_and19_3[0], h_u_arrmul24_fa20_2_xor1[0], h_u_arrmul24_fa18_3_or0[0], h_u_arrmul24_fa19_3_xor1, h_u_arrmul24_fa19_3_or0);
  and_gate and_gate_h_u_arrmul24_and20_3(a[20], b[3], h_u_arrmul24_and20_3);
  fa fa_h_u_arrmul24_fa20_3_out(h_u_arrmul24_and20_3[0], h_u_arrmul24_fa21_2_xor1[0], h_u_arrmul24_fa19_3_or0[0], h_u_arrmul24_fa20_3_xor1, h_u_arrmul24_fa20_3_or0);
  and_gate and_gate_h_u_arrmul24_and21_3(a[21], b[3], h_u_arrmul24_and21_3);
  fa fa_h_u_arrmul24_fa21_3_out(h_u_arrmul24_and21_3[0], h_u_arrmul24_fa22_2_xor1[0], h_u_arrmul24_fa20_3_or0[0], h_u_arrmul24_fa21_3_xor1, h_u_arrmul24_fa21_3_or0);
  and_gate and_gate_h_u_arrmul24_and22_3(a[22], b[3], h_u_arrmul24_and22_3);
  fa fa_h_u_arrmul24_fa22_3_out(h_u_arrmul24_and22_3[0], h_u_arrmul24_fa23_2_xor1[0], h_u_arrmul24_fa21_3_or0[0], h_u_arrmul24_fa22_3_xor1, h_u_arrmul24_fa22_3_or0);
  and_gate and_gate_h_u_arrmul24_and23_3(a[23], b[3], h_u_arrmul24_and23_3);
  fa fa_h_u_arrmul24_fa23_3_out(h_u_arrmul24_and23_3[0], h_u_arrmul24_fa23_2_or0[0], h_u_arrmul24_fa22_3_or0[0], h_u_arrmul24_fa23_3_xor1, h_u_arrmul24_fa23_3_or0);
  and_gate and_gate_h_u_arrmul24_and0_4(a[0], b[4], h_u_arrmul24_and0_4);
  ha ha_h_u_arrmul24_ha0_4_out(h_u_arrmul24_and0_4[0], h_u_arrmul24_fa1_3_xor1[0], h_u_arrmul24_ha0_4_xor0, h_u_arrmul24_ha0_4_and0);
  and_gate and_gate_h_u_arrmul24_and1_4(a[1], b[4], h_u_arrmul24_and1_4);
  fa fa_h_u_arrmul24_fa1_4_out(h_u_arrmul24_and1_4[0], h_u_arrmul24_fa2_3_xor1[0], h_u_arrmul24_ha0_4_and0[0], h_u_arrmul24_fa1_4_xor1, h_u_arrmul24_fa1_4_or0);
  and_gate and_gate_h_u_arrmul24_and2_4(a[2], b[4], h_u_arrmul24_and2_4);
  fa fa_h_u_arrmul24_fa2_4_out(h_u_arrmul24_and2_4[0], h_u_arrmul24_fa3_3_xor1[0], h_u_arrmul24_fa1_4_or0[0], h_u_arrmul24_fa2_4_xor1, h_u_arrmul24_fa2_4_or0);
  and_gate and_gate_h_u_arrmul24_and3_4(a[3], b[4], h_u_arrmul24_and3_4);
  fa fa_h_u_arrmul24_fa3_4_out(h_u_arrmul24_and3_4[0], h_u_arrmul24_fa4_3_xor1[0], h_u_arrmul24_fa2_4_or0[0], h_u_arrmul24_fa3_4_xor1, h_u_arrmul24_fa3_4_or0);
  and_gate and_gate_h_u_arrmul24_and4_4(a[4], b[4], h_u_arrmul24_and4_4);
  fa fa_h_u_arrmul24_fa4_4_out(h_u_arrmul24_and4_4[0], h_u_arrmul24_fa5_3_xor1[0], h_u_arrmul24_fa3_4_or0[0], h_u_arrmul24_fa4_4_xor1, h_u_arrmul24_fa4_4_or0);
  and_gate and_gate_h_u_arrmul24_and5_4(a[5], b[4], h_u_arrmul24_and5_4);
  fa fa_h_u_arrmul24_fa5_4_out(h_u_arrmul24_and5_4[0], h_u_arrmul24_fa6_3_xor1[0], h_u_arrmul24_fa4_4_or0[0], h_u_arrmul24_fa5_4_xor1, h_u_arrmul24_fa5_4_or0);
  and_gate and_gate_h_u_arrmul24_and6_4(a[6], b[4], h_u_arrmul24_and6_4);
  fa fa_h_u_arrmul24_fa6_4_out(h_u_arrmul24_and6_4[0], h_u_arrmul24_fa7_3_xor1[0], h_u_arrmul24_fa5_4_or0[0], h_u_arrmul24_fa6_4_xor1, h_u_arrmul24_fa6_4_or0);
  and_gate and_gate_h_u_arrmul24_and7_4(a[7], b[4], h_u_arrmul24_and7_4);
  fa fa_h_u_arrmul24_fa7_4_out(h_u_arrmul24_and7_4[0], h_u_arrmul24_fa8_3_xor1[0], h_u_arrmul24_fa6_4_or0[0], h_u_arrmul24_fa7_4_xor1, h_u_arrmul24_fa7_4_or0);
  and_gate and_gate_h_u_arrmul24_and8_4(a[8], b[4], h_u_arrmul24_and8_4);
  fa fa_h_u_arrmul24_fa8_4_out(h_u_arrmul24_and8_4[0], h_u_arrmul24_fa9_3_xor1[0], h_u_arrmul24_fa7_4_or0[0], h_u_arrmul24_fa8_4_xor1, h_u_arrmul24_fa8_4_or0);
  and_gate and_gate_h_u_arrmul24_and9_4(a[9], b[4], h_u_arrmul24_and9_4);
  fa fa_h_u_arrmul24_fa9_4_out(h_u_arrmul24_and9_4[0], h_u_arrmul24_fa10_3_xor1[0], h_u_arrmul24_fa8_4_or0[0], h_u_arrmul24_fa9_4_xor1, h_u_arrmul24_fa9_4_or0);
  and_gate and_gate_h_u_arrmul24_and10_4(a[10], b[4], h_u_arrmul24_and10_4);
  fa fa_h_u_arrmul24_fa10_4_out(h_u_arrmul24_and10_4[0], h_u_arrmul24_fa11_3_xor1[0], h_u_arrmul24_fa9_4_or0[0], h_u_arrmul24_fa10_4_xor1, h_u_arrmul24_fa10_4_or0);
  and_gate and_gate_h_u_arrmul24_and11_4(a[11], b[4], h_u_arrmul24_and11_4);
  fa fa_h_u_arrmul24_fa11_4_out(h_u_arrmul24_and11_4[0], h_u_arrmul24_fa12_3_xor1[0], h_u_arrmul24_fa10_4_or0[0], h_u_arrmul24_fa11_4_xor1, h_u_arrmul24_fa11_4_or0);
  and_gate and_gate_h_u_arrmul24_and12_4(a[12], b[4], h_u_arrmul24_and12_4);
  fa fa_h_u_arrmul24_fa12_4_out(h_u_arrmul24_and12_4[0], h_u_arrmul24_fa13_3_xor1[0], h_u_arrmul24_fa11_4_or0[0], h_u_arrmul24_fa12_4_xor1, h_u_arrmul24_fa12_4_or0);
  and_gate and_gate_h_u_arrmul24_and13_4(a[13], b[4], h_u_arrmul24_and13_4);
  fa fa_h_u_arrmul24_fa13_4_out(h_u_arrmul24_and13_4[0], h_u_arrmul24_fa14_3_xor1[0], h_u_arrmul24_fa12_4_or0[0], h_u_arrmul24_fa13_4_xor1, h_u_arrmul24_fa13_4_or0);
  and_gate and_gate_h_u_arrmul24_and14_4(a[14], b[4], h_u_arrmul24_and14_4);
  fa fa_h_u_arrmul24_fa14_4_out(h_u_arrmul24_and14_4[0], h_u_arrmul24_fa15_3_xor1[0], h_u_arrmul24_fa13_4_or0[0], h_u_arrmul24_fa14_4_xor1, h_u_arrmul24_fa14_4_or0);
  and_gate and_gate_h_u_arrmul24_and15_4(a[15], b[4], h_u_arrmul24_and15_4);
  fa fa_h_u_arrmul24_fa15_4_out(h_u_arrmul24_and15_4[0], h_u_arrmul24_fa16_3_xor1[0], h_u_arrmul24_fa14_4_or0[0], h_u_arrmul24_fa15_4_xor1, h_u_arrmul24_fa15_4_or0);
  and_gate and_gate_h_u_arrmul24_and16_4(a[16], b[4], h_u_arrmul24_and16_4);
  fa fa_h_u_arrmul24_fa16_4_out(h_u_arrmul24_and16_4[0], h_u_arrmul24_fa17_3_xor1[0], h_u_arrmul24_fa15_4_or0[0], h_u_arrmul24_fa16_4_xor1, h_u_arrmul24_fa16_4_or0);
  and_gate and_gate_h_u_arrmul24_and17_4(a[17], b[4], h_u_arrmul24_and17_4);
  fa fa_h_u_arrmul24_fa17_4_out(h_u_arrmul24_and17_4[0], h_u_arrmul24_fa18_3_xor1[0], h_u_arrmul24_fa16_4_or0[0], h_u_arrmul24_fa17_4_xor1, h_u_arrmul24_fa17_4_or0);
  and_gate and_gate_h_u_arrmul24_and18_4(a[18], b[4], h_u_arrmul24_and18_4);
  fa fa_h_u_arrmul24_fa18_4_out(h_u_arrmul24_and18_4[0], h_u_arrmul24_fa19_3_xor1[0], h_u_arrmul24_fa17_4_or0[0], h_u_arrmul24_fa18_4_xor1, h_u_arrmul24_fa18_4_or0);
  and_gate and_gate_h_u_arrmul24_and19_4(a[19], b[4], h_u_arrmul24_and19_4);
  fa fa_h_u_arrmul24_fa19_4_out(h_u_arrmul24_and19_4[0], h_u_arrmul24_fa20_3_xor1[0], h_u_arrmul24_fa18_4_or0[0], h_u_arrmul24_fa19_4_xor1, h_u_arrmul24_fa19_4_or0);
  and_gate and_gate_h_u_arrmul24_and20_4(a[20], b[4], h_u_arrmul24_and20_4);
  fa fa_h_u_arrmul24_fa20_4_out(h_u_arrmul24_and20_4[0], h_u_arrmul24_fa21_3_xor1[0], h_u_arrmul24_fa19_4_or0[0], h_u_arrmul24_fa20_4_xor1, h_u_arrmul24_fa20_4_or0);
  and_gate and_gate_h_u_arrmul24_and21_4(a[21], b[4], h_u_arrmul24_and21_4);
  fa fa_h_u_arrmul24_fa21_4_out(h_u_arrmul24_and21_4[0], h_u_arrmul24_fa22_3_xor1[0], h_u_arrmul24_fa20_4_or0[0], h_u_arrmul24_fa21_4_xor1, h_u_arrmul24_fa21_4_or0);
  and_gate and_gate_h_u_arrmul24_and22_4(a[22], b[4], h_u_arrmul24_and22_4);
  fa fa_h_u_arrmul24_fa22_4_out(h_u_arrmul24_and22_4[0], h_u_arrmul24_fa23_3_xor1[0], h_u_arrmul24_fa21_4_or0[0], h_u_arrmul24_fa22_4_xor1, h_u_arrmul24_fa22_4_or0);
  and_gate and_gate_h_u_arrmul24_and23_4(a[23], b[4], h_u_arrmul24_and23_4);
  fa fa_h_u_arrmul24_fa23_4_out(h_u_arrmul24_and23_4[0], h_u_arrmul24_fa23_3_or0[0], h_u_arrmul24_fa22_4_or0[0], h_u_arrmul24_fa23_4_xor1, h_u_arrmul24_fa23_4_or0);
  and_gate and_gate_h_u_arrmul24_and0_5(a[0], b[5], h_u_arrmul24_and0_5);
  ha ha_h_u_arrmul24_ha0_5_out(h_u_arrmul24_and0_5[0], h_u_arrmul24_fa1_4_xor1[0], h_u_arrmul24_ha0_5_xor0, h_u_arrmul24_ha0_5_and0);
  and_gate and_gate_h_u_arrmul24_and1_5(a[1], b[5], h_u_arrmul24_and1_5);
  fa fa_h_u_arrmul24_fa1_5_out(h_u_arrmul24_and1_5[0], h_u_arrmul24_fa2_4_xor1[0], h_u_arrmul24_ha0_5_and0[0], h_u_arrmul24_fa1_5_xor1, h_u_arrmul24_fa1_5_or0);
  and_gate and_gate_h_u_arrmul24_and2_5(a[2], b[5], h_u_arrmul24_and2_5);
  fa fa_h_u_arrmul24_fa2_5_out(h_u_arrmul24_and2_5[0], h_u_arrmul24_fa3_4_xor1[0], h_u_arrmul24_fa1_5_or0[0], h_u_arrmul24_fa2_5_xor1, h_u_arrmul24_fa2_5_or0);
  and_gate and_gate_h_u_arrmul24_and3_5(a[3], b[5], h_u_arrmul24_and3_5);
  fa fa_h_u_arrmul24_fa3_5_out(h_u_arrmul24_and3_5[0], h_u_arrmul24_fa4_4_xor1[0], h_u_arrmul24_fa2_5_or0[0], h_u_arrmul24_fa3_5_xor1, h_u_arrmul24_fa3_5_or0);
  and_gate and_gate_h_u_arrmul24_and4_5(a[4], b[5], h_u_arrmul24_and4_5);
  fa fa_h_u_arrmul24_fa4_5_out(h_u_arrmul24_and4_5[0], h_u_arrmul24_fa5_4_xor1[0], h_u_arrmul24_fa3_5_or0[0], h_u_arrmul24_fa4_5_xor1, h_u_arrmul24_fa4_5_or0);
  and_gate and_gate_h_u_arrmul24_and5_5(a[5], b[5], h_u_arrmul24_and5_5);
  fa fa_h_u_arrmul24_fa5_5_out(h_u_arrmul24_and5_5[0], h_u_arrmul24_fa6_4_xor1[0], h_u_arrmul24_fa4_5_or0[0], h_u_arrmul24_fa5_5_xor1, h_u_arrmul24_fa5_5_or0);
  and_gate and_gate_h_u_arrmul24_and6_5(a[6], b[5], h_u_arrmul24_and6_5);
  fa fa_h_u_arrmul24_fa6_5_out(h_u_arrmul24_and6_5[0], h_u_arrmul24_fa7_4_xor1[0], h_u_arrmul24_fa5_5_or0[0], h_u_arrmul24_fa6_5_xor1, h_u_arrmul24_fa6_5_or0);
  and_gate and_gate_h_u_arrmul24_and7_5(a[7], b[5], h_u_arrmul24_and7_5);
  fa fa_h_u_arrmul24_fa7_5_out(h_u_arrmul24_and7_5[0], h_u_arrmul24_fa8_4_xor1[0], h_u_arrmul24_fa6_5_or0[0], h_u_arrmul24_fa7_5_xor1, h_u_arrmul24_fa7_5_or0);
  and_gate and_gate_h_u_arrmul24_and8_5(a[8], b[5], h_u_arrmul24_and8_5);
  fa fa_h_u_arrmul24_fa8_5_out(h_u_arrmul24_and8_5[0], h_u_arrmul24_fa9_4_xor1[0], h_u_arrmul24_fa7_5_or0[0], h_u_arrmul24_fa8_5_xor1, h_u_arrmul24_fa8_5_or0);
  and_gate and_gate_h_u_arrmul24_and9_5(a[9], b[5], h_u_arrmul24_and9_5);
  fa fa_h_u_arrmul24_fa9_5_out(h_u_arrmul24_and9_5[0], h_u_arrmul24_fa10_4_xor1[0], h_u_arrmul24_fa8_5_or0[0], h_u_arrmul24_fa9_5_xor1, h_u_arrmul24_fa9_5_or0);
  and_gate and_gate_h_u_arrmul24_and10_5(a[10], b[5], h_u_arrmul24_and10_5);
  fa fa_h_u_arrmul24_fa10_5_out(h_u_arrmul24_and10_5[0], h_u_arrmul24_fa11_4_xor1[0], h_u_arrmul24_fa9_5_or0[0], h_u_arrmul24_fa10_5_xor1, h_u_arrmul24_fa10_5_or0);
  and_gate and_gate_h_u_arrmul24_and11_5(a[11], b[5], h_u_arrmul24_and11_5);
  fa fa_h_u_arrmul24_fa11_5_out(h_u_arrmul24_and11_5[0], h_u_arrmul24_fa12_4_xor1[0], h_u_arrmul24_fa10_5_or0[0], h_u_arrmul24_fa11_5_xor1, h_u_arrmul24_fa11_5_or0);
  and_gate and_gate_h_u_arrmul24_and12_5(a[12], b[5], h_u_arrmul24_and12_5);
  fa fa_h_u_arrmul24_fa12_5_out(h_u_arrmul24_and12_5[0], h_u_arrmul24_fa13_4_xor1[0], h_u_arrmul24_fa11_5_or0[0], h_u_arrmul24_fa12_5_xor1, h_u_arrmul24_fa12_5_or0);
  and_gate and_gate_h_u_arrmul24_and13_5(a[13], b[5], h_u_arrmul24_and13_5);
  fa fa_h_u_arrmul24_fa13_5_out(h_u_arrmul24_and13_5[0], h_u_arrmul24_fa14_4_xor1[0], h_u_arrmul24_fa12_5_or0[0], h_u_arrmul24_fa13_5_xor1, h_u_arrmul24_fa13_5_or0);
  and_gate and_gate_h_u_arrmul24_and14_5(a[14], b[5], h_u_arrmul24_and14_5);
  fa fa_h_u_arrmul24_fa14_5_out(h_u_arrmul24_and14_5[0], h_u_arrmul24_fa15_4_xor1[0], h_u_arrmul24_fa13_5_or0[0], h_u_arrmul24_fa14_5_xor1, h_u_arrmul24_fa14_5_or0);
  and_gate and_gate_h_u_arrmul24_and15_5(a[15], b[5], h_u_arrmul24_and15_5);
  fa fa_h_u_arrmul24_fa15_5_out(h_u_arrmul24_and15_5[0], h_u_arrmul24_fa16_4_xor1[0], h_u_arrmul24_fa14_5_or0[0], h_u_arrmul24_fa15_5_xor1, h_u_arrmul24_fa15_5_or0);
  and_gate and_gate_h_u_arrmul24_and16_5(a[16], b[5], h_u_arrmul24_and16_5);
  fa fa_h_u_arrmul24_fa16_5_out(h_u_arrmul24_and16_5[0], h_u_arrmul24_fa17_4_xor1[0], h_u_arrmul24_fa15_5_or0[0], h_u_arrmul24_fa16_5_xor1, h_u_arrmul24_fa16_5_or0);
  and_gate and_gate_h_u_arrmul24_and17_5(a[17], b[5], h_u_arrmul24_and17_5);
  fa fa_h_u_arrmul24_fa17_5_out(h_u_arrmul24_and17_5[0], h_u_arrmul24_fa18_4_xor1[0], h_u_arrmul24_fa16_5_or0[0], h_u_arrmul24_fa17_5_xor1, h_u_arrmul24_fa17_5_or0);
  and_gate and_gate_h_u_arrmul24_and18_5(a[18], b[5], h_u_arrmul24_and18_5);
  fa fa_h_u_arrmul24_fa18_5_out(h_u_arrmul24_and18_5[0], h_u_arrmul24_fa19_4_xor1[0], h_u_arrmul24_fa17_5_or0[0], h_u_arrmul24_fa18_5_xor1, h_u_arrmul24_fa18_5_or0);
  and_gate and_gate_h_u_arrmul24_and19_5(a[19], b[5], h_u_arrmul24_and19_5);
  fa fa_h_u_arrmul24_fa19_5_out(h_u_arrmul24_and19_5[0], h_u_arrmul24_fa20_4_xor1[0], h_u_arrmul24_fa18_5_or0[0], h_u_arrmul24_fa19_5_xor1, h_u_arrmul24_fa19_5_or0);
  and_gate and_gate_h_u_arrmul24_and20_5(a[20], b[5], h_u_arrmul24_and20_5);
  fa fa_h_u_arrmul24_fa20_5_out(h_u_arrmul24_and20_5[0], h_u_arrmul24_fa21_4_xor1[0], h_u_arrmul24_fa19_5_or0[0], h_u_arrmul24_fa20_5_xor1, h_u_arrmul24_fa20_5_or0);
  and_gate and_gate_h_u_arrmul24_and21_5(a[21], b[5], h_u_arrmul24_and21_5);
  fa fa_h_u_arrmul24_fa21_5_out(h_u_arrmul24_and21_5[0], h_u_arrmul24_fa22_4_xor1[0], h_u_arrmul24_fa20_5_or0[0], h_u_arrmul24_fa21_5_xor1, h_u_arrmul24_fa21_5_or0);
  and_gate and_gate_h_u_arrmul24_and22_5(a[22], b[5], h_u_arrmul24_and22_5);
  fa fa_h_u_arrmul24_fa22_5_out(h_u_arrmul24_and22_5[0], h_u_arrmul24_fa23_4_xor1[0], h_u_arrmul24_fa21_5_or0[0], h_u_arrmul24_fa22_5_xor1, h_u_arrmul24_fa22_5_or0);
  and_gate and_gate_h_u_arrmul24_and23_5(a[23], b[5], h_u_arrmul24_and23_5);
  fa fa_h_u_arrmul24_fa23_5_out(h_u_arrmul24_and23_5[0], h_u_arrmul24_fa23_4_or0[0], h_u_arrmul24_fa22_5_or0[0], h_u_arrmul24_fa23_5_xor1, h_u_arrmul24_fa23_5_or0);
  and_gate and_gate_h_u_arrmul24_and0_6(a[0], b[6], h_u_arrmul24_and0_6);
  ha ha_h_u_arrmul24_ha0_6_out(h_u_arrmul24_and0_6[0], h_u_arrmul24_fa1_5_xor1[0], h_u_arrmul24_ha0_6_xor0, h_u_arrmul24_ha0_6_and0);
  and_gate and_gate_h_u_arrmul24_and1_6(a[1], b[6], h_u_arrmul24_and1_6);
  fa fa_h_u_arrmul24_fa1_6_out(h_u_arrmul24_and1_6[0], h_u_arrmul24_fa2_5_xor1[0], h_u_arrmul24_ha0_6_and0[0], h_u_arrmul24_fa1_6_xor1, h_u_arrmul24_fa1_6_or0);
  and_gate and_gate_h_u_arrmul24_and2_6(a[2], b[6], h_u_arrmul24_and2_6);
  fa fa_h_u_arrmul24_fa2_6_out(h_u_arrmul24_and2_6[0], h_u_arrmul24_fa3_5_xor1[0], h_u_arrmul24_fa1_6_or0[0], h_u_arrmul24_fa2_6_xor1, h_u_arrmul24_fa2_6_or0);
  and_gate and_gate_h_u_arrmul24_and3_6(a[3], b[6], h_u_arrmul24_and3_6);
  fa fa_h_u_arrmul24_fa3_6_out(h_u_arrmul24_and3_6[0], h_u_arrmul24_fa4_5_xor1[0], h_u_arrmul24_fa2_6_or0[0], h_u_arrmul24_fa3_6_xor1, h_u_arrmul24_fa3_6_or0);
  and_gate and_gate_h_u_arrmul24_and4_6(a[4], b[6], h_u_arrmul24_and4_6);
  fa fa_h_u_arrmul24_fa4_6_out(h_u_arrmul24_and4_6[0], h_u_arrmul24_fa5_5_xor1[0], h_u_arrmul24_fa3_6_or0[0], h_u_arrmul24_fa4_6_xor1, h_u_arrmul24_fa4_6_or0);
  and_gate and_gate_h_u_arrmul24_and5_6(a[5], b[6], h_u_arrmul24_and5_6);
  fa fa_h_u_arrmul24_fa5_6_out(h_u_arrmul24_and5_6[0], h_u_arrmul24_fa6_5_xor1[0], h_u_arrmul24_fa4_6_or0[0], h_u_arrmul24_fa5_6_xor1, h_u_arrmul24_fa5_6_or0);
  and_gate and_gate_h_u_arrmul24_and6_6(a[6], b[6], h_u_arrmul24_and6_6);
  fa fa_h_u_arrmul24_fa6_6_out(h_u_arrmul24_and6_6[0], h_u_arrmul24_fa7_5_xor1[0], h_u_arrmul24_fa5_6_or0[0], h_u_arrmul24_fa6_6_xor1, h_u_arrmul24_fa6_6_or0);
  and_gate and_gate_h_u_arrmul24_and7_6(a[7], b[6], h_u_arrmul24_and7_6);
  fa fa_h_u_arrmul24_fa7_6_out(h_u_arrmul24_and7_6[0], h_u_arrmul24_fa8_5_xor1[0], h_u_arrmul24_fa6_6_or0[0], h_u_arrmul24_fa7_6_xor1, h_u_arrmul24_fa7_6_or0);
  and_gate and_gate_h_u_arrmul24_and8_6(a[8], b[6], h_u_arrmul24_and8_6);
  fa fa_h_u_arrmul24_fa8_6_out(h_u_arrmul24_and8_6[0], h_u_arrmul24_fa9_5_xor1[0], h_u_arrmul24_fa7_6_or0[0], h_u_arrmul24_fa8_6_xor1, h_u_arrmul24_fa8_6_or0);
  and_gate and_gate_h_u_arrmul24_and9_6(a[9], b[6], h_u_arrmul24_and9_6);
  fa fa_h_u_arrmul24_fa9_6_out(h_u_arrmul24_and9_6[0], h_u_arrmul24_fa10_5_xor1[0], h_u_arrmul24_fa8_6_or0[0], h_u_arrmul24_fa9_6_xor1, h_u_arrmul24_fa9_6_or0);
  and_gate and_gate_h_u_arrmul24_and10_6(a[10], b[6], h_u_arrmul24_and10_6);
  fa fa_h_u_arrmul24_fa10_6_out(h_u_arrmul24_and10_6[0], h_u_arrmul24_fa11_5_xor1[0], h_u_arrmul24_fa9_6_or0[0], h_u_arrmul24_fa10_6_xor1, h_u_arrmul24_fa10_6_or0);
  and_gate and_gate_h_u_arrmul24_and11_6(a[11], b[6], h_u_arrmul24_and11_6);
  fa fa_h_u_arrmul24_fa11_6_out(h_u_arrmul24_and11_6[0], h_u_arrmul24_fa12_5_xor1[0], h_u_arrmul24_fa10_6_or0[0], h_u_arrmul24_fa11_6_xor1, h_u_arrmul24_fa11_6_or0);
  and_gate and_gate_h_u_arrmul24_and12_6(a[12], b[6], h_u_arrmul24_and12_6);
  fa fa_h_u_arrmul24_fa12_6_out(h_u_arrmul24_and12_6[0], h_u_arrmul24_fa13_5_xor1[0], h_u_arrmul24_fa11_6_or0[0], h_u_arrmul24_fa12_6_xor1, h_u_arrmul24_fa12_6_or0);
  and_gate and_gate_h_u_arrmul24_and13_6(a[13], b[6], h_u_arrmul24_and13_6);
  fa fa_h_u_arrmul24_fa13_6_out(h_u_arrmul24_and13_6[0], h_u_arrmul24_fa14_5_xor1[0], h_u_arrmul24_fa12_6_or0[0], h_u_arrmul24_fa13_6_xor1, h_u_arrmul24_fa13_6_or0);
  and_gate and_gate_h_u_arrmul24_and14_6(a[14], b[6], h_u_arrmul24_and14_6);
  fa fa_h_u_arrmul24_fa14_6_out(h_u_arrmul24_and14_6[0], h_u_arrmul24_fa15_5_xor1[0], h_u_arrmul24_fa13_6_or0[0], h_u_arrmul24_fa14_6_xor1, h_u_arrmul24_fa14_6_or0);
  and_gate and_gate_h_u_arrmul24_and15_6(a[15], b[6], h_u_arrmul24_and15_6);
  fa fa_h_u_arrmul24_fa15_6_out(h_u_arrmul24_and15_6[0], h_u_arrmul24_fa16_5_xor1[0], h_u_arrmul24_fa14_6_or0[0], h_u_arrmul24_fa15_6_xor1, h_u_arrmul24_fa15_6_or0);
  and_gate and_gate_h_u_arrmul24_and16_6(a[16], b[6], h_u_arrmul24_and16_6);
  fa fa_h_u_arrmul24_fa16_6_out(h_u_arrmul24_and16_6[0], h_u_arrmul24_fa17_5_xor1[0], h_u_arrmul24_fa15_6_or0[0], h_u_arrmul24_fa16_6_xor1, h_u_arrmul24_fa16_6_or0);
  and_gate and_gate_h_u_arrmul24_and17_6(a[17], b[6], h_u_arrmul24_and17_6);
  fa fa_h_u_arrmul24_fa17_6_out(h_u_arrmul24_and17_6[0], h_u_arrmul24_fa18_5_xor1[0], h_u_arrmul24_fa16_6_or0[0], h_u_arrmul24_fa17_6_xor1, h_u_arrmul24_fa17_6_or0);
  and_gate and_gate_h_u_arrmul24_and18_6(a[18], b[6], h_u_arrmul24_and18_6);
  fa fa_h_u_arrmul24_fa18_6_out(h_u_arrmul24_and18_6[0], h_u_arrmul24_fa19_5_xor1[0], h_u_arrmul24_fa17_6_or0[0], h_u_arrmul24_fa18_6_xor1, h_u_arrmul24_fa18_6_or0);
  and_gate and_gate_h_u_arrmul24_and19_6(a[19], b[6], h_u_arrmul24_and19_6);
  fa fa_h_u_arrmul24_fa19_6_out(h_u_arrmul24_and19_6[0], h_u_arrmul24_fa20_5_xor1[0], h_u_arrmul24_fa18_6_or0[0], h_u_arrmul24_fa19_6_xor1, h_u_arrmul24_fa19_6_or0);
  and_gate and_gate_h_u_arrmul24_and20_6(a[20], b[6], h_u_arrmul24_and20_6);
  fa fa_h_u_arrmul24_fa20_6_out(h_u_arrmul24_and20_6[0], h_u_arrmul24_fa21_5_xor1[0], h_u_arrmul24_fa19_6_or0[0], h_u_arrmul24_fa20_6_xor1, h_u_arrmul24_fa20_6_or0);
  and_gate and_gate_h_u_arrmul24_and21_6(a[21], b[6], h_u_arrmul24_and21_6);
  fa fa_h_u_arrmul24_fa21_6_out(h_u_arrmul24_and21_6[0], h_u_arrmul24_fa22_5_xor1[0], h_u_arrmul24_fa20_6_or0[0], h_u_arrmul24_fa21_6_xor1, h_u_arrmul24_fa21_6_or0);
  and_gate and_gate_h_u_arrmul24_and22_6(a[22], b[6], h_u_arrmul24_and22_6);
  fa fa_h_u_arrmul24_fa22_6_out(h_u_arrmul24_and22_6[0], h_u_arrmul24_fa23_5_xor1[0], h_u_arrmul24_fa21_6_or0[0], h_u_arrmul24_fa22_6_xor1, h_u_arrmul24_fa22_6_or0);
  and_gate and_gate_h_u_arrmul24_and23_6(a[23], b[6], h_u_arrmul24_and23_6);
  fa fa_h_u_arrmul24_fa23_6_out(h_u_arrmul24_and23_6[0], h_u_arrmul24_fa23_5_or0[0], h_u_arrmul24_fa22_6_or0[0], h_u_arrmul24_fa23_6_xor1, h_u_arrmul24_fa23_6_or0);
  and_gate and_gate_h_u_arrmul24_and0_7(a[0], b[7], h_u_arrmul24_and0_7);
  ha ha_h_u_arrmul24_ha0_7_out(h_u_arrmul24_and0_7[0], h_u_arrmul24_fa1_6_xor1[0], h_u_arrmul24_ha0_7_xor0, h_u_arrmul24_ha0_7_and0);
  and_gate and_gate_h_u_arrmul24_and1_7(a[1], b[7], h_u_arrmul24_and1_7);
  fa fa_h_u_arrmul24_fa1_7_out(h_u_arrmul24_and1_7[0], h_u_arrmul24_fa2_6_xor1[0], h_u_arrmul24_ha0_7_and0[0], h_u_arrmul24_fa1_7_xor1, h_u_arrmul24_fa1_7_or0);
  and_gate and_gate_h_u_arrmul24_and2_7(a[2], b[7], h_u_arrmul24_and2_7);
  fa fa_h_u_arrmul24_fa2_7_out(h_u_arrmul24_and2_7[0], h_u_arrmul24_fa3_6_xor1[0], h_u_arrmul24_fa1_7_or0[0], h_u_arrmul24_fa2_7_xor1, h_u_arrmul24_fa2_7_or0);
  and_gate and_gate_h_u_arrmul24_and3_7(a[3], b[7], h_u_arrmul24_and3_7);
  fa fa_h_u_arrmul24_fa3_7_out(h_u_arrmul24_and3_7[0], h_u_arrmul24_fa4_6_xor1[0], h_u_arrmul24_fa2_7_or0[0], h_u_arrmul24_fa3_7_xor1, h_u_arrmul24_fa3_7_or0);
  and_gate and_gate_h_u_arrmul24_and4_7(a[4], b[7], h_u_arrmul24_and4_7);
  fa fa_h_u_arrmul24_fa4_7_out(h_u_arrmul24_and4_7[0], h_u_arrmul24_fa5_6_xor1[0], h_u_arrmul24_fa3_7_or0[0], h_u_arrmul24_fa4_7_xor1, h_u_arrmul24_fa4_7_or0);
  and_gate and_gate_h_u_arrmul24_and5_7(a[5], b[7], h_u_arrmul24_and5_7);
  fa fa_h_u_arrmul24_fa5_7_out(h_u_arrmul24_and5_7[0], h_u_arrmul24_fa6_6_xor1[0], h_u_arrmul24_fa4_7_or0[0], h_u_arrmul24_fa5_7_xor1, h_u_arrmul24_fa5_7_or0);
  and_gate and_gate_h_u_arrmul24_and6_7(a[6], b[7], h_u_arrmul24_and6_7);
  fa fa_h_u_arrmul24_fa6_7_out(h_u_arrmul24_and6_7[0], h_u_arrmul24_fa7_6_xor1[0], h_u_arrmul24_fa5_7_or0[0], h_u_arrmul24_fa6_7_xor1, h_u_arrmul24_fa6_7_or0);
  and_gate and_gate_h_u_arrmul24_and7_7(a[7], b[7], h_u_arrmul24_and7_7);
  fa fa_h_u_arrmul24_fa7_7_out(h_u_arrmul24_and7_7[0], h_u_arrmul24_fa8_6_xor1[0], h_u_arrmul24_fa6_7_or0[0], h_u_arrmul24_fa7_7_xor1, h_u_arrmul24_fa7_7_or0);
  and_gate and_gate_h_u_arrmul24_and8_7(a[8], b[7], h_u_arrmul24_and8_7);
  fa fa_h_u_arrmul24_fa8_7_out(h_u_arrmul24_and8_7[0], h_u_arrmul24_fa9_6_xor1[0], h_u_arrmul24_fa7_7_or0[0], h_u_arrmul24_fa8_7_xor1, h_u_arrmul24_fa8_7_or0);
  and_gate and_gate_h_u_arrmul24_and9_7(a[9], b[7], h_u_arrmul24_and9_7);
  fa fa_h_u_arrmul24_fa9_7_out(h_u_arrmul24_and9_7[0], h_u_arrmul24_fa10_6_xor1[0], h_u_arrmul24_fa8_7_or0[0], h_u_arrmul24_fa9_7_xor1, h_u_arrmul24_fa9_7_or0);
  and_gate and_gate_h_u_arrmul24_and10_7(a[10], b[7], h_u_arrmul24_and10_7);
  fa fa_h_u_arrmul24_fa10_7_out(h_u_arrmul24_and10_7[0], h_u_arrmul24_fa11_6_xor1[0], h_u_arrmul24_fa9_7_or0[0], h_u_arrmul24_fa10_7_xor1, h_u_arrmul24_fa10_7_or0);
  and_gate and_gate_h_u_arrmul24_and11_7(a[11], b[7], h_u_arrmul24_and11_7);
  fa fa_h_u_arrmul24_fa11_7_out(h_u_arrmul24_and11_7[0], h_u_arrmul24_fa12_6_xor1[0], h_u_arrmul24_fa10_7_or0[0], h_u_arrmul24_fa11_7_xor1, h_u_arrmul24_fa11_7_or0);
  and_gate and_gate_h_u_arrmul24_and12_7(a[12], b[7], h_u_arrmul24_and12_7);
  fa fa_h_u_arrmul24_fa12_7_out(h_u_arrmul24_and12_7[0], h_u_arrmul24_fa13_6_xor1[0], h_u_arrmul24_fa11_7_or0[0], h_u_arrmul24_fa12_7_xor1, h_u_arrmul24_fa12_7_or0);
  and_gate and_gate_h_u_arrmul24_and13_7(a[13], b[7], h_u_arrmul24_and13_7);
  fa fa_h_u_arrmul24_fa13_7_out(h_u_arrmul24_and13_7[0], h_u_arrmul24_fa14_6_xor1[0], h_u_arrmul24_fa12_7_or0[0], h_u_arrmul24_fa13_7_xor1, h_u_arrmul24_fa13_7_or0);
  and_gate and_gate_h_u_arrmul24_and14_7(a[14], b[7], h_u_arrmul24_and14_7);
  fa fa_h_u_arrmul24_fa14_7_out(h_u_arrmul24_and14_7[0], h_u_arrmul24_fa15_6_xor1[0], h_u_arrmul24_fa13_7_or0[0], h_u_arrmul24_fa14_7_xor1, h_u_arrmul24_fa14_7_or0);
  and_gate and_gate_h_u_arrmul24_and15_7(a[15], b[7], h_u_arrmul24_and15_7);
  fa fa_h_u_arrmul24_fa15_7_out(h_u_arrmul24_and15_7[0], h_u_arrmul24_fa16_6_xor1[0], h_u_arrmul24_fa14_7_or0[0], h_u_arrmul24_fa15_7_xor1, h_u_arrmul24_fa15_7_or0);
  and_gate and_gate_h_u_arrmul24_and16_7(a[16], b[7], h_u_arrmul24_and16_7);
  fa fa_h_u_arrmul24_fa16_7_out(h_u_arrmul24_and16_7[0], h_u_arrmul24_fa17_6_xor1[0], h_u_arrmul24_fa15_7_or0[0], h_u_arrmul24_fa16_7_xor1, h_u_arrmul24_fa16_7_or0);
  and_gate and_gate_h_u_arrmul24_and17_7(a[17], b[7], h_u_arrmul24_and17_7);
  fa fa_h_u_arrmul24_fa17_7_out(h_u_arrmul24_and17_7[0], h_u_arrmul24_fa18_6_xor1[0], h_u_arrmul24_fa16_7_or0[0], h_u_arrmul24_fa17_7_xor1, h_u_arrmul24_fa17_7_or0);
  and_gate and_gate_h_u_arrmul24_and18_7(a[18], b[7], h_u_arrmul24_and18_7);
  fa fa_h_u_arrmul24_fa18_7_out(h_u_arrmul24_and18_7[0], h_u_arrmul24_fa19_6_xor1[0], h_u_arrmul24_fa17_7_or0[0], h_u_arrmul24_fa18_7_xor1, h_u_arrmul24_fa18_7_or0);
  and_gate and_gate_h_u_arrmul24_and19_7(a[19], b[7], h_u_arrmul24_and19_7);
  fa fa_h_u_arrmul24_fa19_7_out(h_u_arrmul24_and19_7[0], h_u_arrmul24_fa20_6_xor1[0], h_u_arrmul24_fa18_7_or0[0], h_u_arrmul24_fa19_7_xor1, h_u_arrmul24_fa19_7_or0);
  and_gate and_gate_h_u_arrmul24_and20_7(a[20], b[7], h_u_arrmul24_and20_7);
  fa fa_h_u_arrmul24_fa20_7_out(h_u_arrmul24_and20_7[0], h_u_arrmul24_fa21_6_xor1[0], h_u_arrmul24_fa19_7_or0[0], h_u_arrmul24_fa20_7_xor1, h_u_arrmul24_fa20_7_or0);
  and_gate and_gate_h_u_arrmul24_and21_7(a[21], b[7], h_u_arrmul24_and21_7);
  fa fa_h_u_arrmul24_fa21_7_out(h_u_arrmul24_and21_7[0], h_u_arrmul24_fa22_6_xor1[0], h_u_arrmul24_fa20_7_or0[0], h_u_arrmul24_fa21_7_xor1, h_u_arrmul24_fa21_7_or0);
  and_gate and_gate_h_u_arrmul24_and22_7(a[22], b[7], h_u_arrmul24_and22_7);
  fa fa_h_u_arrmul24_fa22_7_out(h_u_arrmul24_and22_7[0], h_u_arrmul24_fa23_6_xor1[0], h_u_arrmul24_fa21_7_or0[0], h_u_arrmul24_fa22_7_xor1, h_u_arrmul24_fa22_7_or0);
  and_gate and_gate_h_u_arrmul24_and23_7(a[23], b[7], h_u_arrmul24_and23_7);
  fa fa_h_u_arrmul24_fa23_7_out(h_u_arrmul24_and23_7[0], h_u_arrmul24_fa23_6_or0[0], h_u_arrmul24_fa22_7_or0[0], h_u_arrmul24_fa23_7_xor1, h_u_arrmul24_fa23_7_or0);
  and_gate and_gate_h_u_arrmul24_and0_8(a[0], b[8], h_u_arrmul24_and0_8);
  ha ha_h_u_arrmul24_ha0_8_out(h_u_arrmul24_and0_8[0], h_u_arrmul24_fa1_7_xor1[0], h_u_arrmul24_ha0_8_xor0, h_u_arrmul24_ha0_8_and0);
  and_gate and_gate_h_u_arrmul24_and1_8(a[1], b[8], h_u_arrmul24_and1_8);
  fa fa_h_u_arrmul24_fa1_8_out(h_u_arrmul24_and1_8[0], h_u_arrmul24_fa2_7_xor1[0], h_u_arrmul24_ha0_8_and0[0], h_u_arrmul24_fa1_8_xor1, h_u_arrmul24_fa1_8_or0);
  and_gate and_gate_h_u_arrmul24_and2_8(a[2], b[8], h_u_arrmul24_and2_8);
  fa fa_h_u_arrmul24_fa2_8_out(h_u_arrmul24_and2_8[0], h_u_arrmul24_fa3_7_xor1[0], h_u_arrmul24_fa1_8_or0[0], h_u_arrmul24_fa2_8_xor1, h_u_arrmul24_fa2_8_or0);
  and_gate and_gate_h_u_arrmul24_and3_8(a[3], b[8], h_u_arrmul24_and3_8);
  fa fa_h_u_arrmul24_fa3_8_out(h_u_arrmul24_and3_8[0], h_u_arrmul24_fa4_7_xor1[0], h_u_arrmul24_fa2_8_or0[0], h_u_arrmul24_fa3_8_xor1, h_u_arrmul24_fa3_8_or0);
  and_gate and_gate_h_u_arrmul24_and4_8(a[4], b[8], h_u_arrmul24_and4_8);
  fa fa_h_u_arrmul24_fa4_8_out(h_u_arrmul24_and4_8[0], h_u_arrmul24_fa5_7_xor1[0], h_u_arrmul24_fa3_8_or0[0], h_u_arrmul24_fa4_8_xor1, h_u_arrmul24_fa4_8_or0);
  and_gate and_gate_h_u_arrmul24_and5_8(a[5], b[8], h_u_arrmul24_and5_8);
  fa fa_h_u_arrmul24_fa5_8_out(h_u_arrmul24_and5_8[0], h_u_arrmul24_fa6_7_xor1[0], h_u_arrmul24_fa4_8_or0[0], h_u_arrmul24_fa5_8_xor1, h_u_arrmul24_fa5_8_or0);
  and_gate and_gate_h_u_arrmul24_and6_8(a[6], b[8], h_u_arrmul24_and6_8);
  fa fa_h_u_arrmul24_fa6_8_out(h_u_arrmul24_and6_8[0], h_u_arrmul24_fa7_7_xor1[0], h_u_arrmul24_fa5_8_or0[0], h_u_arrmul24_fa6_8_xor1, h_u_arrmul24_fa6_8_or0);
  and_gate and_gate_h_u_arrmul24_and7_8(a[7], b[8], h_u_arrmul24_and7_8);
  fa fa_h_u_arrmul24_fa7_8_out(h_u_arrmul24_and7_8[0], h_u_arrmul24_fa8_7_xor1[0], h_u_arrmul24_fa6_8_or0[0], h_u_arrmul24_fa7_8_xor1, h_u_arrmul24_fa7_8_or0);
  and_gate and_gate_h_u_arrmul24_and8_8(a[8], b[8], h_u_arrmul24_and8_8);
  fa fa_h_u_arrmul24_fa8_8_out(h_u_arrmul24_and8_8[0], h_u_arrmul24_fa9_7_xor1[0], h_u_arrmul24_fa7_8_or0[0], h_u_arrmul24_fa8_8_xor1, h_u_arrmul24_fa8_8_or0);
  and_gate and_gate_h_u_arrmul24_and9_8(a[9], b[8], h_u_arrmul24_and9_8);
  fa fa_h_u_arrmul24_fa9_8_out(h_u_arrmul24_and9_8[0], h_u_arrmul24_fa10_7_xor1[0], h_u_arrmul24_fa8_8_or0[0], h_u_arrmul24_fa9_8_xor1, h_u_arrmul24_fa9_8_or0);
  and_gate and_gate_h_u_arrmul24_and10_8(a[10], b[8], h_u_arrmul24_and10_8);
  fa fa_h_u_arrmul24_fa10_8_out(h_u_arrmul24_and10_8[0], h_u_arrmul24_fa11_7_xor1[0], h_u_arrmul24_fa9_8_or0[0], h_u_arrmul24_fa10_8_xor1, h_u_arrmul24_fa10_8_or0);
  and_gate and_gate_h_u_arrmul24_and11_8(a[11], b[8], h_u_arrmul24_and11_8);
  fa fa_h_u_arrmul24_fa11_8_out(h_u_arrmul24_and11_8[0], h_u_arrmul24_fa12_7_xor1[0], h_u_arrmul24_fa10_8_or0[0], h_u_arrmul24_fa11_8_xor1, h_u_arrmul24_fa11_8_or0);
  and_gate and_gate_h_u_arrmul24_and12_8(a[12], b[8], h_u_arrmul24_and12_8);
  fa fa_h_u_arrmul24_fa12_8_out(h_u_arrmul24_and12_8[0], h_u_arrmul24_fa13_7_xor1[0], h_u_arrmul24_fa11_8_or0[0], h_u_arrmul24_fa12_8_xor1, h_u_arrmul24_fa12_8_or0);
  and_gate and_gate_h_u_arrmul24_and13_8(a[13], b[8], h_u_arrmul24_and13_8);
  fa fa_h_u_arrmul24_fa13_8_out(h_u_arrmul24_and13_8[0], h_u_arrmul24_fa14_7_xor1[0], h_u_arrmul24_fa12_8_or0[0], h_u_arrmul24_fa13_8_xor1, h_u_arrmul24_fa13_8_or0);
  and_gate and_gate_h_u_arrmul24_and14_8(a[14], b[8], h_u_arrmul24_and14_8);
  fa fa_h_u_arrmul24_fa14_8_out(h_u_arrmul24_and14_8[0], h_u_arrmul24_fa15_7_xor1[0], h_u_arrmul24_fa13_8_or0[0], h_u_arrmul24_fa14_8_xor1, h_u_arrmul24_fa14_8_or0);
  and_gate and_gate_h_u_arrmul24_and15_8(a[15], b[8], h_u_arrmul24_and15_8);
  fa fa_h_u_arrmul24_fa15_8_out(h_u_arrmul24_and15_8[0], h_u_arrmul24_fa16_7_xor1[0], h_u_arrmul24_fa14_8_or0[0], h_u_arrmul24_fa15_8_xor1, h_u_arrmul24_fa15_8_or0);
  and_gate and_gate_h_u_arrmul24_and16_8(a[16], b[8], h_u_arrmul24_and16_8);
  fa fa_h_u_arrmul24_fa16_8_out(h_u_arrmul24_and16_8[0], h_u_arrmul24_fa17_7_xor1[0], h_u_arrmul24_fa15_8_or0[0], h_u_arrmul24_fa16_8_xor1, h_u_arrmul24_fa16_8_or0);
  and_gate and_gate_h_u_arrmul24_and17_8(a[17], b[8], h_u_arrmul24_and17_8);
  fa fa_h_u_arrmul24_fa17_8_out(h_u_arrmul24_and17_8[0], h_u_arrmul24_fa18_7_xor1[0], h_u_arrmul24_fa16_8_or0[0], h_u_arrmul24_fa17_8_xor1, h_u_arrmul24_fa17_8_or0);
  and_gate and_gate_h_u_arrmul24_and18_8(a[18], b[8], h_u_arrmul24_and18_8);
  fa fa_h_u_arrmul24_fa18_8_out(h_u_arrmul24_and18_8[0], h_u_arrmul24_fa19_7_xor1[0], h_u_arrmul24_fa17_8_or0[0], h_u_arrmul24_fa18_8_xor1, h_u_arrmul24_fa18_8_or0);
  and_gate and_gate_h_u_arrmul24_and19_8(a[19], b[8], h_u_arrmul24_and19_8);
  fa fa_h_u_arrmul24_fa19_8_out(h_u_arrmul24_and19_8[0], h_u_arrmul24_fa20_7_xor1[0], h_u_arrmul24_fa18_8_or0[0], h_u_arrmul24_fa19_8_xor1, h_u_arrmul24_fa19_8_or0);
  and_gate and_gate_h_u_arrmul24_and20_8(a[20], b[8], h_u_arrmul24_and20_8);
  fa fa_h_u_arrmul24_fa20_8_out(h_u_arrmul24_and20_8[0], h_u_arrmul24_fa21_7_xor1[0], h_u_arrmul24_fa19_8_or0[0], h_u_arrmul24_fa20_8_xor1, h_u_arrmul24_fa20_8_or0);
  and_gate and_gate_h_u_arrmul24_and21_8(a[21], b[8], h_u_arrmul24_and21_8);
  fa fa_h_u_arrmul24_fa21_8_out(h_u_arrmul24_and21_8[0], h_u_arrmul24_fa22_7_xor1[0], h_u_arrmul24_fa20_8_or0[0], h_u_arrmul24_fa21_8_xor1, h_u_arrmul24_fa21_8_or0);
  and_gate and_gate_h_u_arrmul24_and22_8(a[22], b[8], h_u_arrmul24_and22_8);
  fa fa_h_u_arrmul24_fa22_8_out(h_u_arrmul24_and22_8[0], h_u_arrmul24_fa23_7_xor1[0], h_u_arrmul24_fa21_8_or0[0], h_u_arrmul24_fa22_8_xor1, h_u_arrmul24_fa22_8_or0);
  and_gate and_gate_h_u_arrmul24_and23_8(a[23], b[8], h_u_arrmul24_and23_8);
  fa fa_h_u_arrmul24_fa23_8_out(h_u_arrmul24_and23_8[0], h_u_arrmul24_fa23_7_or0[0], h_u_arrmul24_fa22_8_or0[0], h_u_arrmul24_fa23_8_xor1, h_u_arrmul24_fa23_8_or0);
  and_gate and_gate_h_u_arrmul24_and0_9(a[0], b[9], h_u_arrmul24_and0_9);
  ha ha_h_u_arrmul24_ha0_9_out(h_u_arrmul24_and0_9[0], h_u_arrmul24_fa1_8_xor1[0], h_u_arrmul24_ha0_9_xor0, h_u_arrmul24_ha0_9_and0);
  and_gate and_gate_h_u_arrmul24_and1_9(a[1], b[9], h_u_arrmul24_and1_9);
  fa fa_h_u_arrmul24_fa1_9_out(h_u_arrmul24_and1_9[0], h_u_arrmul24_fa2_8_xor1[0], h_u_arrmul24_ha0_9_and0[0], h_u_arrmul24_fa1_9_xor1, h_u_arrmul24_fa1_9_or0);
  and_gate and_gate_h_u_arrmul24_and2_9(a[2], b[9], h_u_arrmul24_and2_9);
  fa fa_h_u_arrmul24_fa2_9_out(h_u_arrmul24_and2_9[0], h_u_arrmul24_fa3_8_xor1[0], h_u_arrmul24_fa1_9_or0[0], h_u_arrmul24_fa2_9_xor1, h_u_arrmul24_fa2_9_or0);
  and_gate and_gate_h_u_arrmul24_and3_9(a[3], b[9], h_u_arrmul24_and3_9);
  fa fa_h_u_arrmul24_fa3_9_out(h_u_arrmul24_and3_9[0], h_u_arrmul24_fa4_8_xor1[0], h_u_arrmul24_fa2_9_or0[0], h_u_arrmul24_fa3_9_xor1, h_u_arrmul24_fa3_9_or0);
  and_gate and_gate_h_u_arrmul24_and4_9(a[4], b[9], h_u_arrmul24_and4_9);
  fa fa_h_u_arrmul24_fa4_9_out(h_u_arrmul24_and4_9[0], h_u_arrmul24_fa5_8_xor1[0], h_u_arrmul24_fa3_9_or0[0], h_u_arrmul24_fa4_9_xor1, h_u_arrmul24_fa4_9_or0);
  and_gate and_gate_h_u_arrmul24_and5_9(a[5], b[9], h_u_arrmul24_and5_9);
  fa fa_h_u_arrmul24_fa5_9_out(h_u_arrmul24_and5_9[0], h_u_arrmul24_fa6_8_xor1[0], h_u_arrmul24_fa4_9_or0[0], h_u_arrmul24_fa5_9_xor1, h_u_arrmul24_fa5_9_or0);
  and_gate and_gate_h_u_arrmul24_and6_9(a[6], b[9], h_u_arrmul24_and6_9);
  fa fa_h_u_arrmul24_fa6_9_out(h_u_arrmul24_and6_9[0], h_u_arrmul24_fa7_8_xor1[0], h_u_arrmul24_fa5_9_or0[0], h_u_arrmul24_fa6_9_xor1, h_u_arrmul24_fa6_9_or0);
  and_gate and_gate_h_u_arrmul24_and7_9(a[7], b[9], h_u_arrmul24_and7_9);
  fa fa_h_u_arrmul24_fa7_9_out(h_u_arrmul24_and7_9[0], h_u_arrmul24_fa8_8_xor1[0], h_u_arrmul24_fa6_9_or0[0], h_u_arrmul24_fa7_9_xor1, h_u_arrmul24_fa7_9_or0);
  and_gate and_gate_h_u_arrmul24_and8_9(a[8], b[9], h_u_arrmul24_and8_9);
  fa fa_h_u_arrmul24_fa8_9_out(h_u_arrmul24_and8_9[0], h_u_arrmul24_fa9_8_xor1[0], h_u_arrmul24_fa7_9_or0[0], h_u_arrmul24_fa8_9_xor1, h_u_arrmul24_fa8_9_or0);
  and_gate and_gate_h_u_arrmul24_and9_9(a[9], b[9], h_u_arrmul24_and9_9);
  fa fa_h_u_arrmul24_fa9_9_out(h_u_arrmul24_and9_9[0], h_u_arrmul24_fa10_8_xor1[0], h_u_arrmul24_fa8_9_or0[0], h_u_arrmul24_fa9_9_xor1, h_u_arrmul24_fa9_9_or0);
  and_gate and_gate_h_u_arrmul24_and10_9(a[10], b[9], h_u_arrmul24_and10_9);
  fa fa_h_u_arrmul24_fa10_9_out(h_u_arrmul24_and10_9[0], h_u_arrmul24_fa11_8_xor1[0], h_u_arrmul24_fa9_9_or0[0], h_u_arrmul24_fa10_9_xor1, h_u_arrmul24_fa10_9_or0);
  and_gate and_gate_h_u_arrmul24_and11_9(a[11], b[9], h_u_arrmul24_and11_9);
  fa fa_h_u_arrmul24_fa11_9_out(h_u_arrmul24_and11_9[0], h_u_arrmul24_fa12_8_xor1[0], h_u_arrmul24_fa10_9_or0[0], h_u_arrmul24_fa11_9_xor1, h_u_arrmul24_fa11_9_or0);
  and_gate and_gate_h_u_arrmul24_and12_9(a[12], b[9], h_u_arrmul24_and12_9);
  fa fa_h_u_arrmul24_fa12_9_out(h_u_arrmul24_and12_9[0], h_u_arrmul24_fa13_8_xor1[0], h_u_arrmul24_fa11_9_or0[0], h_u_arrmul24_fa12_9_xor1, h_u_arrmul24_fa12_9_or0);
  and_gate and_gate_h_u_arrmul24_and13_9(a[13], b[9], h_u_arrmul24_and13_9);
  fa fa_h_u_arrmul24_fa13_9_out(h_u_arrmul24_and13_9[0], h_u_arrmul24_fa14_8_xor1[0], h_u_arrmul24_fa12_9_or0[0], h_u_arrmul24_fa13_9_xor1, h_u_arrmul24_fa13_9_or0);
  and_gate and_gate_h_u_arrmul24_and14_9(a[14], b[9], h_u_arrmul24_and14_9);
  fa fa_h_u_arrmul24_fa14_9_out(h_u_arrmul24_and14_9[0], h_u_arrmul24_fa15_8_xor1[0], h_u_arrmul24_fa13_9_or0[0], h_u_arrmul24_fa14_9_xor1, h_u_arrmul24_fa14_9_or0);
  and_gate and_gate_h_u_arrmul24_and15_9(a[15], b[9], h_u_arrmul24_and15_9);
  fa fa_h_u_arrmul24_fa15_9_out(h_u_arrmul24_and15_9[0], h_u_arrmul24_fa16_8_xor1[0], h_u_arrmul24_fa14_9_or0[0], h_u_arrmul24_fa15_9_xor1, h_u_arrmul24_fa15_9_or0);
  and_gate and_gate_h_u_arrmul24_and16_9(a[16], b[9], h_u_arrmul24_and16_9);
  fa fa_h_u_arrmul24_fa16_9_out(h_u_arrmul24_and16_9[0], h_u_arrmul24_fa17_8_xor1[0], h_u_arrmul24_fa15_9_or0[0], h_u_arrmul24_fa16_9_xor1, h_u_arrmul24_fa16_9_or0);
  and_gate and_gate_h_u_arrmul24_and17_9(a[17], b[9], h_u_arrmul24_and17_9);
  fa fa_h_u_arrmul24_fa17_9_out(h_u_arrmul24_and17_9[0], h_u_arrmul24_fa18_8_xor1[0], h_u_arrmul24_fa16_9_or0[0], h_u_arrmul24_fa17_9_xor1, h_u_arrmul24_fa17_9_or0);
  and_gate and_gate_h_u_arrmul24_and18_9(a[18], b[9], h_u_arrmul24_and18_9);
  fa fa_h_u_arrmul24_fa18_9_out(h_u_arrmul24_and18_9[0], h_u_arrmul24_fa19_8_xor1[0], h_u_arrmul24_fa17_9_or0[0], h_u_arrmul24_fa18_9_xor1, h_u_arrmul24_fa18_9_or0);
  and_gate and_gate_h_u_arrmul24_and19_9(a[19], b[9], h_u_arrmul24_and19_9);
  fa fa_h_u_arrmul24_fa19_9_out(h_u_arrmul24_and19_9[0], h_u_arrmul24_fa20_8_xor1[0], h_u_arrmul24_fa18_9_or0[0], h_u_arrmul24_fa19_9_xor1, h_u_arrmul24_fa19_9_or0);
  and_gate and_gate_h_u_arrmul24_and20_9(a[20], b[9], h_u_arrmul24_and20_9);
  fa fa_h_u_arrmul24_fa20_9_out(h_u_arrmul24_and20_9[0], h_u_arrmul24_fa21_8_xor1[0], h_u_arrmul24_fa19_9_or0[0], h_u_arrmul24_fa20_9_xor1, h_u_arrmul24_fa20_9_or0);
  and_gate and_gate_h_u_arrmul24_and21_9(a[21], b[9], h_u_arrmul24_and21_9);
  fa fa_h_u_arrmul24_fa21_9_out(h_u_arrmul24_and21_9[0], h_u_arrmul24_fa22_8_xor1[0], h_u_arrmul24_fa20_9_or0[0], h_u_arrmul24_fa21_9_xor1, h_u_arrmul24_fa21_9_or0);
  and_gate and_gate_h_u_arrmul24_and22_9(a[22], b[9], h_u_arrmul24_and22_9);
  fa fa_h_u_arrmul24_fa22_9_out(h_u_arrmul24_and22_9[0], h_u_arrmul24_fa23_8_xor1[0], h_u_arrmul24_fa21_9_or0[0], h_u_arrmul24_fa22_9_xor1, h_u_arrmul24_fa22_9_or0);
  and_gate and_gate_h_u_arrmul24_and23_9(a[23], b[9], h_u_arrmul24_and23_9);
  fa fa_h_u_arrmul24_fa23_9_out(h_u_arrmul24_and23_9[0], h_u_arrmul24_fa23_8_or0[0], h_u_arrmul24_fa22_9_or0[0], h_u_arrmul24_fa23_9_xor1, h_u_arrmul24_fa23_9_or0);
  and_gate and_gate_h_u_arrmul24_and0_10(a[0], b[10], h_u_arrmul24_and0_10);
  ha ha_h_u_arrmul24_ha0_10_out(h_u_arrmul24_and0_10[0], h_u_arrmul24_fa1_9_xor1[0], h_u_arrmul24_ha0_10_xor0, h_u_arrmul24_ha0_10_and0);
  and_gate and_gate_h_u_arrmul24_and1_10(a[1], b[10], h_u_arrmul24_and1_10);
  fa fa_h_u_arrmul24_fa1_10_out(h_u_arrmul24_and1_10[0], h_u_arrmul24_fa2_9_xor1[0], h_u_arrmul24_ha0_10_and0[0], h_u_arrmul24_fa1_10_xor1, h_u_arrmul24_fa1_10_or0);
  and_gate and_gate_h_u_arrmul24_and2_10(a[2], b[10], h_u_arrmul24_and2_10);
  fa fa_h_u_arrmul24_fa2_10_out(h_u_arrmul24_and2_10[0], h_u_arrmul24_fa3_9_xor1[0], h_u_arrmul24_fa1_10_or0[0], h_u_arrmul24_fa2_10_xor1, h_u_arrmul24_fa2_10_or0);
  and_gate and_gate_h_u_arrmul24_and3_10(a[3], b[10], h_u_arrmul24_and3_10);
  fa fa_h_u_arrmul24_fa3_10_out(h_u_arrmul24_and3_10[0], h_u_arrmul24_fa4_9_xor1[0], h_u_arrmul24_fa2_10_or0[0], h_u_arrmul24_fa3_10_xor1, h_u_arrmul24_fa3_10_or0);
  and_gate and_gate_h_u_arrmul24_and4_10(a[4], b[10], h_u_arrmul24_and4_10);
  fa fa_h_u_arrmul24_fa4_10_out(h_u_arrmul24_and4_10[0], h_u_arrmul24_fa5_9_xor1[0], h_u_arrmul24_fa3_10_or0[0], h_u_arrmul24_fa4_10_xor1, h_u_arrmul24_fa4_10_or0);
  and_gate and_gate_h_u_arrmul24_and5_10(a[5], b[10], h_u_arrmul24_and5_10);
  fa fa_h_u_arrmul24_fa5_10_out(h_u_arrmul24_and5_10[0], h_u_arrmul24_fa6_9_xor1[0], h_u_arrmul24_fa4_10_or0[0], h_u_arrmul24_fa5_10_xor1, h_u_arrmul24_fa5_10_or0);
  and_gate and_gate_h_u_arrmul24_and6_10(a[6], b[10], h_u_arrmul24_and6_10);
  fa fa_h_u_arrmul24_fa6_10_out(h_u_arrmul24_and6_10[0], h_u_arrmul24_fa7_9_xor1[0], h_u_arrmul24_fa5_10_or0[0], h_u_arrmul24_fa6_10_xor1, h_u_arrmul24_fa6_10_or0);
  and_gate and_gate_h_u_arrmul24_and7_10(a[7], b[10], h_u_arrmul24_and7_10);
  fa fa_h_u_arrmul24_fa7_10_out(h_u_arrmul24_and7_10[0], h_u_arrmul24_fa8_9_xor1[0], h_u_arrmul24_fa6_10_or0[0], h_u_arrmul24_fa7_10_xor1, h_u_arrmul24_fa7_10_or0);
  and_gate and_gate_h_u_arrmul24_and8_10(a[8], b[10], h_u_arrmul24_and8_10);
  fa fa_h_u_arrmul24_fa8_10_out(h_u_arrmul24_and8_10[0], h_u_arrmul24_fa9_9_xor1[0], h_u_arrmul24_fa7_10_or0[0], h_u_arrmul24_fa8_10_xor1, h_u_arrmul24_fa8_10_or0);
  and_gate and_gate_h_u_arrmul24_and9_10(a[9], b[10], h_u_arrmul24_and9_10);
  fa fa_h_u_arrmul24_fa9_10_out(h_u_arrmul24_and9_10[0], h_u_arrmul24_fa10_9_xor1[0], h_u_arrmul24_fa8_10_or0[0], h_u_arrmul24_fa9_10_xor1, h_u_arrmul24_fa9_10_or0);
  and_gate and_gate_h_u_arrmul24_and10_10(a[10], b[10], h_u_arrmul24_and10_10);
  fa fa_h_u_arrmul24_fa10_10_out(h_u_arrmul24_and10_10[0], h_u_arrmul24_fa11_9_xor1[0], h_u_arrmul24_fa9_10_or0[0], h_u_arrmul24_fa10_10_xor1, h_u_arrmul24_fa10_10_or0);
  and_gate and_gate_h_u_arrmul24_and11_10(a[11], b[10], h_u_arrmul24_and11_10);
  fa fa_h_u_arrmul24_fa11_10_out(h_u_arrmul24_and11_10[0], h_u_arrmul24_fa12_9_xor1[0], h_u_arrmul24_fa10_10_or0[0], h_u_arrmul24_fa11_10_xor1, h_u_arrmul24_fa11_10_or0);
  and_gate and_gate_h_u_arrmul24_and12_10(a[12], b[10], h_u_arrmul24_and12_10);
  fa fa_h_u_arrmul24_fa12_10_out(h_u_arrmul24_and12_10[0], h_u_arrmul24_fa13_9_xor1[0], h_u_arrmul24_fa11_10_or0[0], h_u_arrmul24_fa12_10_xor1, h_u_arrmul24_fa12_10_or0);
  and_gate and_gate_h_u_arrmul24_and13_10(a[13], b[10], h_u_arrmul24_and13_10);
  fa fa_h_u_arrmul24_fa13_10_out(h_u_arrmul24_and13_10[0], h_u_arrmul24_fa14_9_xor1[0], h_u_arrmul24_fa12_10_or0[0], h_u_arrmul24_fa13_10_xor1, h_u_arrmul24_fa13_10_or0);
  and_gate and_gate_h_u_arrmul24_and14_10(a[14], b[10], h_u_arrmul24_and14_10);
  fa fa_h_u_arrmul24_fa14_10_out(h_u_arrmul24_and14_10[0], h_u_arrmul24_fa15_9_xor1[0], h_u_arrmul24_fa13_10_or0[0], h_u_arrmul24_fa14_10_xor1, h_u_arrmul24_fa14_10_or0);
  and_gate and_gate_h_u_arrmul24_and15_10(a[15], b[10], h_u_arrmul24_and15_10);
  fa fa_h_u_arrmul24_fa15_10_out(h_u_arrmul24_and15_10[0], h_u_arrmul24_fa16_9_xor1[0], h_u_arrmul24_fa14_10_or0[0], h_u_arrmul24_fa15_10_xor1, h_u_arrmul24_fa15_10_or0);
  and_gate and_gate_h_u_arrmul24_and16_10(a[16], b[10], h_u_arrmul24_and16_10);
  fa fa_h_u_arrmul24_fa16_10_out(h_u_arrmul24_and16_10[0], h_u_arrmul24_fa17_9_xor1[0], h_u_arrmul24_fa15_10_or0[0], h_u_arrmul24_fa16_10_xor1, h_u_arrmul24_fa16_10_or0);
  and_gate and_gate_h_u_arrmul24_and17_10(a[17], b[10], h_u_arrmul24_and17_10);
  fa fa_h_u_arrmul24_fa17_10_out(h_u_arrmul24_and17_10[0], h_u_arrmul24_fa18_9_xor1[0], h_u_arrmul24_fa16_10_or0[0], h_u_arrmul24_fa17_10_xor1, h_u_arrmul24_fa17_10_or0);
  and_gate and_gate_h_u_arrmul24_and18_10(a[18], b[10], h_u_arrmul24_and18_10);
  fa fa_h_u_arrmul24_fa18_10_out(h_u_arrmul24_and18_10[0], h_u_arrmul24_fa19_9_xor1[0], h_u_arrmul24_fa17_10_or0[0], h_u_arrmul24_fa18_10_xor1, h_u_arrmul24_fa18_10_or0);
  and_gate and_gate_h_u_arrmul24_and19_10(a[19], b[10], h_u_arrmul24_and19_10);
  fa fa_h_u_arrmul24_fa19_10_out(h_u_arrmul24_and19_10[0], h_u_arrmul24_fa20_9_xor1[0], h_u_arrmul24_fa18_10_or0[0], h_u_arrmul24_fa19_10_xor1, h_u_arrmul24_fa19_10_or0);
  and_gate and_gate_h_u_arrmul24_and20_10(a[20], b[10], h_u_arrmul24_and20_10);
  fa fa_h_u_arrmul24_fa20_10_out(h_u_arrmul24_and20_10[0], h_u_arrmul24_fa21_9_xor1[0], h_u_arrmul24_fa19_10_or0[0], h_u_arrmul24_fa20_10_xor1, h_u_arrmul24_fa20_10_or0);
  and_gate and_gate_h_u_arrmul24_and21_10(a[21], b[10], h_u_arrmul24_and21_10);
  fa fa_h_u_arrmul24_fa21_10_out(h_u_arrmul24_and21_10[0], h_u_arrmul24_fa22_9_xor1[0], h_u_arrmul24_fa20_10_or0[0], h_u_arrmul24_fa21_10_xor1, h_u_arrmul24_fa21_10_or0);
  and_gate and_gate_h_u_arrmul24_and22_10(a[22], b[10], h_u_arrmul24_and22_10);
  fa fa_h_u_arrmul24_fa22_10_out(h_u_arrmul24_and22_10[0], h_u_arrmul24_fa23_9_xor1[0], h_u_arrmul24_fa21_10_or0[0], h_u_arrmul24_fa22_10_xor1, h_u_arrmul24_fa22_10_or0);
  and_gate and_gate_h_u_arrmul24_and23_10(a[23], b[10], h_u_arrmul24_and23_10);
  fa fa_h_u_arrmul24_fa23_10_out(h_u_arrmul24_and23_10[0], h_u_arrmul24_fa23_9_or0[0], h_u_arrmul24_fa22_10_or0[0], h_u_arrmul24_fa23_10_xor1, h_u_arrmul24_fa23_10_or0);
  and_gate and_gate_h_u_arrmul24_and0_11(a[0], b[11], h_u_arrmul24_and0_11);
  ha ha_h_u_arrmul24_ha0_11_out(h_u_arrmul24_and0_11[0], h_u_arrmul24_fa1_10_xor1[0], h_u_arrmul24_ha0_11_xor0, h_u_arrmul24_ha0_11_and0);
  and_gate and_gate_h_u_arrmul24_and1_11(a[1], b[11], h_u_arrmul24_and1_11);
  fa fa_h_u_arrmul24_fa1_11_out(h_u_arrmul24_and1_11[0], h_u_arrmul24_fa2_10_xor1[0], h_u_arrmul24_ha0_11_and0[0], h_u_arrmul24_fa1_11_xor1, h_u_arrmul24_fa1_11_or0);
  and_gate and_gate_h_u_arrmul24_and2_11(a[2], b[11], h_u_arrmul24_and2_11);
  fa fa_h_u_arrmul24_fa2_11_out(h_u_arrmul24_and2_11[0], h_u_arrmul24_fa3_10_xor1[0], h_u_arrmul24_fa1_11_or0[0], h_u_arrmul24_fa2_11_xor1, h_u_arrmul24_fa2_11_or0);
  and_gate and_gate_h_u_arrmul24_and3_11(a[3], b[11], h_u_arrmul24_and3_11);
  fa fa_h_u_arrmul24_fa3_11_out(h_u_arrmul24_and3_11[0], h_u_arrmul24_fa4_10_xor1[0], h_u_arrmul24_fa2_11_or0[0], h_u_arrmul24_fa3_11_xor1, h_u_arrmul24_fa3_11_or0);
  and_gate and_gate_h_u_arrmul24_and4_11(a[4], b[11], h_u_arrmul24_and4_11);
  fa fa_h_u_arrmul24_fa4_11_out(h_u_arrmul24_and4_11[0], h_u_arrmul24_fa5_10_xor1[0], h_u_arrmul24_fa3_11_or0[0], h_u_arrmul24_fa4_11_xor1, h_u_arrmul24_fa4_11_or0);
  and_gate and_gate_h_u_arrmul24_and5_11(a[5], b[11], h_u_arrmul24_and5_11);
  fa fa_h_u_arrmul24_fa5_11_out(h_u_arrmul24_and5_11[0], h_u_arrmul24_fa6_10_xor1[0], h_u_arrmul24_fa4_11_or0[0], h_u_arrmul24_fa5_11_xor1, h_u_arrmul24_fa5_11_or0);
  and_gate and_gate_h_u_arrmul24_and6_11(a[6], b[11], h_u_arrmul24_and6_11);
  fa fa_h_u_arrmul24_fa6_11_out(h_u_arrmul24_and6_11[0], h_u_arrmul24_fa7_10_xor1[0], h_u_arrmul24_fa5_11_or0[0], h_u_arrmul24_fa6_11_xor1, h_u_arrmul24_fa6_11_or0);
  and_gate and_gate_h_u_arrmul24_and7_11(a[7], b[11], h_u_arrmul24_and7_11);
  fa fa_h_u_arrmul24_fa7_11_out(h_u_arrmul24_and7_11[0], h_u_arrmul24_fa8_10_xor1[0], h_u_arrmul24_fa6_11_or0[0], h_u_arrmul24_fa7_11_xor1, h_u_arrmul24_fa7_11_or0);
  and_gate and_gate_h_u_arrmul24_and8_11(a[8], b[11], h_u_arrmul24_and8_11);
  fa fa_h_u_arrmul24_fa8_11_out(h_u_arrmul24_and8_11[0], h_u_arrmul24_fa9_10_xor1[0], h_u_arrmul24_fa7_11_or0[0], h_u_arrmul24_fa8_11_xor1, h_u_arrmul24_fa8_11_or0);
  and_gate and_gate_h_u_arrmul24_and9_11(a[9], b[11], h_u_arrmul24_and9_11);
  fa fa_h_u_arrmul24_fa9_11_out(h_u_arrmul24_and9_11[0], h_u_arrmul24_fa10_10_xor1[0], h_u_arrmul24_fa8_11_or0[0], h_u_arrmul24_fa9_11_xor1, h_u_arrmul24_fa9_11_or0);
  and_gate and_gate_h_u_arrmul24_and10_11(a[10], b[11], h_u_arrmul24_and10_11);
  fa fa_h_u_arrmul24_fa10_11_out(h_u_arrmul24_and10_11[0], h_u_arrmul24_fa11_10_xor1[0], h_u_arrmul24_fa9_11_or0[0], h_u_arrmul24_fa10_11_xor1, h_u_arrmul24_fa10_11_or0);
  and_gate and_gate_h_u_arrmul24_and11_11(a[11], b[11], h_u_arrmul24_and11_11);
  fa fa_h_u_arrmul24_fa11_11_out(h_u_arrmul24_and11_11[0], h_u_arrmul24_fa12_10_xor1[0], h_u_arrmul24_fa10_11_or0[0], h_u_arrmul24_fa11_11_xor1, h_u_arrmul24_fa11_11_or0);
  and_gate and_gate_h_u_arrmul24_and12_11(a[12], b[11], h_u_arrmul24_and12_11);
  fa fa_h_u_arrmul24_fa12_11_out(h_u_arrmul24_and12_11[0], h_u_arrmul24_fa13_10_xor1[0], h_u_arrmul24_fa11_11_or0[0], h_u_arrmul24_fa12_11_xor1, h_u_arrmul24_fa12_11_or0);
  and_gate and_gate_h_u_arrmul24_and13_11(a[13], b[11], h_u_arrmul24_and13_11);
  fa fa_h_u_arrmul24_fa13_11_out(h_u_arrmul24_and13_11[0], h_u_arrmul24_fa14_10_xor1[0], h_u_arrmul24_fa12_11_or0[0], h_u_arrmul24_fa13_11_xor1, h_u_arrmul24_fa13_11_or0);
  and_gate and_gate_h_u_arrmul24_and14_11(a[14], b[11], h_u_arrmul24_and14_11);
  fa fa_h_u_arrmul24_fa14_11_out(h_u_arrmul24_and14_11[0], h_u_arrmul24_fa15_10_xor1[0], h_u_arrmul24_fa13_11_or0[0], h_u_arrmul24_fa14_11_xor1, h_u_arrmul24_fa14_11_or0);
  and_gate and_gate_h_u_arrmul24_and15_11(a[15], b[11], h_u_arrmul24_and15_11);
  fa fa_h_u_arrmul24_fa15_11_out(h_u_arrmul24_and15_11[0], h_u_arrmul24_fa16_10_xor1[0], h_u_arrmul24_fa14_11_or0[0], h_u_arrmul24_fa15_11_xor1, h_u_arrmul24_fa15_11_or0);
  and_gate and_gate_h_u_arrmul24_and16_11(a[16], b[11], h_u_arrmul24_and16_11);
  fa fa_h_u_arrmul24_fa16_11_out(h_u_arrmul24_and16_11[0], h_u_arrmul24_fa17_10_xor1[0], h_u_arrmul24_fa15_11_or0[0], h_u_arrmul24_fa16_11_xor1, h_u_arrmul24_fa16_11_or0);
  and_gate and_gate_h_u_arrmul24_and17_11(a[17], b[11], h_u_arrmul24_and17_11);
  fa fa_h_u_arrmul24_fa17_11_out(h_u_arrmul24_and17_11[0], h_u_arrmul24_fa18_10_xor1[0], h_u_arrmul24_fa16_11_or0[0], h_u_arrmul24_fa17_11_xor1, h_u_arrmul24_fa17_11_or0);
  and_gate and_gate_h_u_arrmul24_and18_11(a[18], b[11], h_u_arrmul24_and18_11);
  fa fa_h_u_arrmul24_fa18_11_out(h_u_arrmul24_and18_11[0], h_u_arrmul24_fa19_10_xor1[0], h_u_arrmul24_fa17_11_or0[0], h_u_arrmul24_fa18_11_xor1, h_u_arrmul24_fa18_11_or0);
  and_gate and_gate_h_u_arrmul24_and19_11(a[19], b[11], h_u_arrmul24_and19_11);
  fa fa_h_u_arrmul24_fa19_11_out(h_u_arrmul24_and19_11[0], h_u_arrmul24_fa20_10_xor1[0], h_u_arrmul24_fa18_11_or0[0], h_u_arrmul24_fa19_11_xor1, h_u_arrmul24_fa19_11_or0);
  and_gate and_gate_h_u_arrmul24_and20_11(a[20], b[11], h_u_arrmul24_and20_11);
  fa fa_h_u_arrmul24_fa20_11_out(h_u_arrmul24_and20_11[0], h_u_arrmul24_fa21_10_xor1[0], h_u_arrmul24_fa19_11_or0[0], h_u_arrmul24_fa20_11_xor1, h_u_arrmul24_fa20_11_or0);
  and_gate and_gate_h_u_arrmul24_and21_11(a[21], b[11], h_u_arrmul24_and21_11);
  fa fa_h_u_arrmul24_fa21_11_out(h_u_arrmul24_and21_11[0], h_u_arrmul24_fa22_10_xor1[0], h_u_arrmul24_fa20_11_or0[0], h_u_arrmul24_fa21_11_xor1, h_u_arrmul24_fa21_11_or0);
  and_gate and_gate_h_u_arrmul24_and22_11(a[22], b[11], h_u_arrmul24_and22_11);
  fa fa_h_u_arrmul24_fa22_11_out(h_u_arrmul24_and22_11[0], h_u_arrmul24_fa23_10_xor1[0], h_u_arrmul24_fa21_11_or0[0], h_u_arrmul24_fa22_11_xor1, h_u_arrmul24_fa22_11_or0);
  and_gate and_gate_h_u_arrmul24_and23_11(a[23], b[11], h_u_arrmul24_and23_11);
  fa fa_h_u_arrmul24_fa23_11_out(h_u_arrmul24_and23_11[0], h_u_arrmul24_fa23_10_or0[0], h_u_arrmul24_fa22_11_or0[0], h_u_arrmul24_fa23_11_xor1, h_u_arrmul24_fa23_11_or0);
  and_gate and_gate_h_u_arrmul24_and0_12(a[0], b[12], h_u_arrmul24_and0_12);
  ha ha_h_u_arrmul24_ha0_12_out(h_u_arrmul24_and0_12[0], h_u_arrmul24_fa1_11_xor1[0], h_u_arrmul24_ha0_12_xor0, h_u_arrmul24_ha0_12_and0);
  and_gate and_gate_h_u_arrmul24_and1_12(a[1], b[12], h_u_arrmul24_and1_12);
  fa fa_h_u_arrmul24_fa1_12_out(h_u_arrmul24_and1_12[0], h_u_arrmul24_fa2_11_xor1[0], h_u_arrmul24_ha0_12_and0[0], h_u_arrmul24_fa1_12_xor1, h_u_arrmul24_fa1_12_or0);
  and_gate and_gate_h_u_arrmul24_and2_12(a[2], b[12], h_u_arrmul24_and2_12);
  fa fa_h_u_arrmul24_fa2_12_out(h_u_arrmul24_and2_12[0], h_u_arrmul24_fa3_11_xor1[0], h_u_arrmul24_fa1_12_or0[0], h_u_arrmul24_fa2_12_xor1, h_u_arrmul24_fa2_12_or0);
  and_gate and_gate_h_u_arrmul24_and3_12(a[3], b[12], h_u_arrmul24_and3_12);
  fa fa_h_u_arrmul24_fa3_12_out(h_u_arrmul24_and3_12[0], h_u_arrmul24_fa4_11_xor1[0], h_u_arrmul24_fa2_12_or0[0], h_u_arrmul24_fa3_12_xor1, h_u_arrmul24_fa3_12_or0);
  and_gate and_gate_h_u_arrmul24_and4_12(a[4], b[12], h_u_arrmul24_and4_12);
  fa fa_h_u_arrmul24_fa4_12_out(h_u_arrmul24_and4_12[0], h_u_arrmul24_fa5_11_xor1[0], h_u_arrmul24_fa3_12_or0[0], h_u_arrmul24_fa4_12_xor1, h_u_arrmul24_fa4_12_or0);
  and_gate and_gate_h_u_arrmul24_and5_12(a[5], b[12], h_u_arrmul24_and5_12);
  fa fa_h_u_arrmul24_fa5_12_out(h_u_arrmul24_and5_12[0], h_u_arrmul24_fa6_11_xor1[0], h_u_arrmul24_fa4_12_or0[0], h_u_arrmul24_fa5_12_xor1, h_u_arrmul24_fa5_12_or0);
  and_gate and_gate_h_u_arrmul24_and6_12(a[6], b[12], h_u_arrmul24_and6_12);
  fa fa_h_u_arrmul24_fa6_12_out(h_u_arrmul24_and6_12[0], h_u_arrmul24_fa7_11_xor1[0], h_u_arrmul24_fa5_12_or0[0], h_u_arrmul24_fa6_12_xor1, h_u_arrmul24_fa6_12_or0);
  and_gate and_gate_h_u_arrmul24_and7_12(a[7], b[12], h_u_arrmul24_and7_12);
  fa fa_h_u_arrmul24_fa7_12_out(h_u_arrmul24_and7_12[0], h_u_arrmul24_fa8_11_xor1[0], h_u_arrmul24_fa6_12_or0[0], h_u_arrmul24_fa7_12_xor1, h_u_arrmul24_fa7_12_or0);
  and_gate and_gate_h_u_arrmul24_and8_12(a[8], b[12], h_u_arrmul24_and8_12);
  fa fa_h_u_arrmul24_fa8_12_out(h_u_arrmul24_and8_12[0], h_u_arrmul24_fa9_11_xor1[0], h_u_arrmul24_fa7_12_or0[0], h_u_arrmul24_fa8_12_xor1, h_u_arrmul24_fa8_12_or0);
  and_gate and_gate_h_u_arrmul24_and9_12(a[9], b[12], h_u_arrmul24_and9_12);
  fa fa_h_u_arrmul24_fa9_12_out(h_u_arrmul24_and9_12[0], h_u_arrmul24_fa10_11_xor1[0], h_u_arrmul24_fa8_12_or0[0], h_u_arrmul24_fa9_12_xor1, h_u_arrmul24_fa9_12_or0);
  and_gate and_gate_h_u_arrmul24_and10_12(a[10], b[12], h_u_arrmul24_and10_12);
  fa fa_h_u_arrmul24_fa10_12_out(h_u_arrmul24_and10_12[0], h_u_arrmul24_fa11_11_xor1[0], h_u_arrmul24_fa9_12_or0[0], h_u_arrmul24_fa10_12_xor1, h_u_arrmul24_fa10_12_or0);
  and_gate and_gate_h_u_arrmul24_and11_12(a[11], b[12], h_u_arrmul24_and11_12);
  fa fa_h_u_arrmul24_fa11_12_out(h_u_arrmul24_and11_12[0], h_u_arrmul24_fa12_11_xor1[0], h_u_arrmul24_fa10_12_or0[0], h_u_arrmul24_fa11_12_xor1, h_u_arrmul24_fa11_12_or0);
  and_gate and_gate_h_u_arrmul24_and12_12(a[12], b[12], h_u_arrmul24_and12_12);
  fa fa_h_u_arrmul24_fa12_12_out(h_u_arrmul24_and12_12[0], h_u_arrmul24_fa13_11_xor1[0], h_u_arrmul24_fa11_12_or0[0], h_u_arrmul24_fa12_12_xor1, h_u_arrmul24_fa12_12_or0);
  and_gate and_gate_h_u_arrmul24_and13_12(a[13], b[12], h_u_arrmul24_and13_12);
  fa fa_h_u_arrmul24_fa13_12_out(h_u_arrmul24_and13_12[0], h_u_arrmul24_fa14_11_xor1[0], h_u_arrmul24_fa12_12_or0[0], h_u_arrmul24_fa13_12_xor1, h_u_arrmul24_fa13_12_or0);
  and_gate and_gate_h_u_arrmul24_and14_12(a[14], b[12], h_u_arrmul24_and14_12);
  fa fa_h_u_arrmul24_fa14_12_out(h_u_arrmul24_and14_12[0], h_u_arrmul24_fa15_11_xor1[0], h_u_arrmul24_fa13_12_or0[0], h_u_arrmul24_fa14_12_xor1, h_u_arrmul24_fa14_12_or0);
  and_gate and_gate_h_u_arrmul24_and15_12(a[15], b[12], h_u_arrmul24_and15_12);
  fa fa_h_u_arrmul24_fa15_12_out(h_u_arrmul24_and15_12[0], h_u_arrmul24_fa16_11_xor1[0], h_u_arrmul24_fa14_12_or0[0], h_u_arrmul24_fa15_12_xor1, h_u_arrmul24_fa15_12_or0);
  and_gate and_gate_h_u_arrmul24_and16_12(a[16], b[12], h_u_arrmul24_and16_12);
  fa fa_h_u_arrmul24_fa16_12_out(h_u_arrmul24_and16_12[0], h_u_arrmul24_fa17_11_xor1[0], h_u_arrmul24_fa15_12_or0[0], h_u_arrmul24_fa16_12_xor1, h_u_arrmul24_fa16_12_or0);
  and_gate and_gate_h_u_arrmul24_and17_12(a[17], b[12], h_u_arrmul24_and17_12);
  fa fa_h_u_arrmul24_fa17_12_out(h_u_arrmul24_and17_12[0], h_u_arrmul24_fa18_11_xor1[0], h_u_arrmul24_fa16_12_or0[0], h_u_arrmul24_fa17_12_xor1, h_u_arrmul24_fa17_12_or0);
  and_gate and_gate_h_u_arrmul24_and18_12(a[18], b[12], h_u_arrmul24_and18_12);
  fa fa_h_u_arrmul24_fa18_12_out(h_u_arrmul24_and18_12[0], h_u_arrmul24_fa19_11_xor1[0], h_u_arrmul24_fa17_12_or0[0], h_u_arrmul24_fa18_12_xor1, h_u_arrmul24_fa18_12_or0);
  and_gate and_gate_h_u_arrmul24_and19_12(a[19], b[12], h_u_arrmul24_and19_12);
  fa fa_h_u_arrmul24_fa19_12_out(h_u_arrmul24_and19_12[0], h_u_arrmul24_fa20_11_xor1[0], h_u_arrmul24_fa18_12_or0[0], h_u_arrmul24_fa19_12_xor1, h_u_arrmul24_fa19_12_or0);
  and_gate and_gate_h_u_arrmul24_and20_12(a[20], b[12], h_u_arrmul24_and20_12);
  fa fa_h_u_arrmul24_fa20_12_out(h_u_arrmul24_and20_12[0], h_u_arrmul24_fa21_11_xor1[0], h_u_arrmul24_fa19_12_or0[0], h_u_arrmul24_fa20_12_xor1, h_u_arrmul24_fa20_12_or0);
  and_gate and_gate_h_u_arrmul24_and21_12(a[21], b[12], h_u_arrmul24_and21_12);
  fa fa_h_u_arrmul24_fa21_12_out(h_u_arrmul24_and21_12[0], h_u_arrmul24_fa22_11_xor1[0], h_u_arrmul24_fa20_12_or0[0], h_u_arrmul24_fa21_12_xor1, h_u_arrmul24_fa21_12_or0);
  and_gate and_gate_h_u_arrmul24_and22_12(a[22], b[12], h_u_arrmul24_and22_12);
  fa fa_h_u_arrmul24_fa22_12_out(h_u_arrmul24_and22_12[0], h_u_arrmul24_fa23_11_xor1[0], h_u_arrmul24_fa21_12_or0[0], h_u_arrmul24_fa22_12_xor1, h_u_arrmul24_fa22_12_or0);
  and_gate and_gate_h_u_arrmul24_and23_12(a[23], b[12], h_u_arrmul24_and23_12);
  fa fa_h_u_arrmul24_fa23_12_out(h_u_arrmul24_and23_12[0], h_u_arrmul24_fa23_11_or0[0], h_u_arrmul24_fa22_12_or0[0], h_u_arrmul24_fa23_12_xor1, h_u_arrmul24_fa23_12_or0);
  and_gate and_gate_h_u_arrmul24_and0_13(a[0], b[13], h_u_arrmul24_and0_13);
  ha ha_h_u_arrmul24_ha0_13_out(h_u_arrmul24_and0_13[0], h_u_arrmul24_fa1_12_xor1[0], h_u_arrmul24_ha0_13_xor0, h_u_arrmul24_ha0_13_and0);
  and_gate and_gate_h_u_arrmul24_and1_13(a[1], b[13], h_u_arrmul24_and1_13);
  fa fa_h_u_arrmul24_fa1_13_out(h_u_arrmul24_and1_13[0], h_u_arrmul24_fa2_12_xor1[0], h_u_arrmul24_ha0_13_and0[0], h_u_arrmul24_fa1_13_xor1, h_u_arrmul24_fa1_13_or0);
  and_gate and_gate_h_u_arrmul24_and2_13(a[2], b[13], h_u_arrmul24_and2_13);
  fa fa_h_u_arrmul24_fa2_13_out(h_u_arrmul24_and2_13[0], h_u_arrmul24_fa3_12_xor1[0], h_u_arrmul24_fa1_13_or0[0], h_u_arrmul24_fa2_13_xor1, h_u_arrmul24_fa2_13_or0);
  and_gate and_gate_h_u_arrmul24_and3_13(a[3], b[13], h_u_arrmul24_and3_13);
  fa fa_h_u_arrmul24_fa3_13_out(h_u_arrmul24_and3_13[0], h_u_arrmul24_fa4_12_xor1[0], h_u_arrmul24_fa2_13_or0[0], h_u_arrmul24_fa3_13_xor1, h_u_arrmul24_fa3_13_or0);
  and_gate and_gate_h_u_arrmul24_and4_13(a[4], b[13], h_u_arrmul24_and4_13);
  fa fa_h_u_arrmul24_fa4_13_out(h_u_arrmul24_and4_13[0], h_u_arrmul24_fa5_12_xor1[0], h_u_arrmul24_fa3_13_or0[0], h_u_arrmul24_fa4_13_xor1, h_u_arrmul24_fa4_13_or0);
  and_gate and_gate_h_u_arrmul24_and5_13(a[5], b[13], h_u_arrmul24_and5_13);
  fa fa_h_u_arrmul24_fa5_13_out(h_u_arrmul24_and5_13[0], h_u_arrmul24_fa6_12_xor1[0], h_u_arrmul24_fa4_13_or0[0], h_u_arrmul24_fa5_13_xor1, h_u_arrmul24_fa5_13_or0);
  and_gate and_gate_h_u_arrmul24_and6_13(a[6], b[13], h_u_arrmul24_and6_13);
  fa fa_h_u_arrmul24_fa6_13_out(h_u_arrmul24_and6_13[0], h_u_arrmul24_fa7_12_xor1[0], h_u_arrmul24_fa5_13_or0[0], h_u_arrmul24_fa6_13_xor1, h_u_arrmul24_fa6_13_or0);
  and_gate and_gate_h_u_arrmul24_and7_13(a[7], b[13], h_u_arrmul24_and7_13);
  fa fa_h_u_arrmul24_fa7_13_out(h_u_arrmul24_and7_13[0], h_u_arrmul24_fa8_12_xor1[0], h_u_arrmul24_fa6_13_or0[0], h_u_arrmul24_fa7_13_xor1, h_u_arrmul24_fa7_13_or0);
  and_gate and_gate_h_u_arrmul24_and8_13(a[8], b[13], h_u_arrmul24_and8_13);
  fa fa_h_u_arrmul24_fa8_13_out(h_u_arrmul24_and8_13[0], h_u_arrmul24_fa9_12_xor1[0], h_u_arrmul24_fa7_13_or0[0], h_u_arrmul24_fa8_13_xor1, h_u_arrmul24_fa8_13_or0);
  and_gate and_gate_h_u_arrmul24_and9_13(a[9], b[13], h_u_arrmul24_and9_13);
  fa fa_h_u_arrmul24_fa9_13_out(h_u_arrmul24_and9_13[0], h_u_arrmul24_fa10_12_xor1[0], h_u_arrmul24_fa8_13_or0[0], h_u_arrmul24_fa9_13_xor1, h_u_arrmul24_fa9_13_or0);
  and_gate and_gate_h_u_arrmul24_and10_13(a[10], b[13], h_u_arrmul24_and10_13);
  fa fa_h_u_arrmul24_fa10_13_out(h_u_arrmul24_and10_13[0], h_u_arrmul24_fa11_12_xor1[0], h_u_arrmul24_fa9_13_or0[0], h_u_arrmul24_fa10_13_xor1, h_u_arrmul24_fa10_13_or0);
  and_gate and_gate_h_u_arrmul24_and11_13(a[11], b[13], h_u_arrmul24_and11_13);
  fa fa_h_u_arrmul24_fa11_13_out(h_u_arrmul24_and11_13[0], h_u_arrmul24_fa12_12_xor1[0], h_u_arrmul24_fa10_13_or0[0], h_u_arrmul24_fa11_13_xor1, h_u_arrmul24_fa11_13_or0);
  and_gate and_gate_h_u_arrmul24_and12_13(a[12], b[13], h_u_arrmul24_and12_13);
  fa fa_h_u_arrmul24_fa12_13_out(h_u_arrmul24_and12_13[0], h_u_arrmul24_fa13_12_xor1[0], h_u_arrmul24_fa11_13_or0[0], h_u_arrmul24_fa12_13_xor1, h_u_arrmul24_fa12_13_or0);
  and_gate and_gate_h_u_arrmul24_and13_13(a[13], b[13], h_u_arrmul24_and13_13);
  fa fa_h_u_arrmul24_fa13_13_out(h_u_arrmul24_and13_13[0], h_u_arrmul24_fa14_12_xor1[0], h_u_arrmul24_fa12_13_or0[0], h_u_arrmul24_fa13_13_xor1, h_u_arrmul24_fa13_13_or0);
  and_gate and_gate_h_u_arrmul24_and14_13(a[14], b[13], h_u_arrmul24_and14_13);
  fa fa_h_u_arrmul24_fa14_13_out(h_u_arrmul24_and14_13[0], h_u_arrmul24_fa15_12_xor1[0], h_u_arrmul24_fa13_13_or0[0], h_u_arrmul24_fa14_13_xor1, h_u_arrmul24_fa14_13_or0);
  and_gate and_gate_h_u_arrmul24_and15_13(a[15], b[13], h_u_arrmul24_and15_13);
  fa fa_h_u_arrmul24_fa15_13_out(h_u_arrmul24_and15_13[0], h_u_arrmul24_fa16_12_xor1[0], h_u_arrmul24_fa14_13_or0[0], h_u_arrmul24_fa15_13_xor1, h_u_arrmul24_fa15_13_or0);
  and_gate and_gate_h_u_arrmul24_and16_13(a[16], b[13], h_u_arrmul24_and16_13);
  fa fa_h_u_arrmul24_fa16_13_out(h_u_arrmul24_and16_13[0], h_u_arrmul24_fa17_12_xor1[0], h_u_arrmul24_fa15_13_or0[0], h_u_arrmul24_fa16_13_xor1, h_u_arrmul24_fa16_13_or0);
  and_gate and_gate_h_u_arrmul24_and17_13(a[17], b[13], h_u_arrmul24_and17_13);
  fa fa_h_u_arrmul24_fa17_13_out(h_u_arrmul24_and17_13[0], h_u_arrmul24_fa18_12_xor1[0], h_u_arrmul24_fa16_13_or0[0], h_u_arrmul24_fa17_13_xor1, h_u_arrmul24_fa17_13_or0);
  and_gate and_gate_h_u_arrmul24_and18_13(a[18], b[13], h_u_arrmul24_and18_13);
  fa fa_h_u_arrmul24_fa18_13_out(h_u_arrmul24_and18_13[0], h_u_arrmul24_fa19_12_xor1[0], h_u_arrmul24_fa17_13_or0[0], h_u_arrmul24_fa18_13_xor1, h_u_arrmul24_fa18_13_or0);
  and_gate and_gate_h_u_arrmul24_and19_13(a[19], b[13], h_u_arrmul24_and19_13);
  fa fa_h_u_arrmul24_fa19_13_out(h_u_arrmul24_and19_13[0], h_u_arrmul24_fa20_12_xor1[0], h_u_arrmul24_fa18_13_or0[0], h_u_arrmul24_fa19_13_xor1, h_u_arrmul24_fa19_13_or0);
  and_gate and_gate_h_u_arrmul24_and20_13(a[20], b[13], h_u_arrmul24_and20_13);
  fa fa_h_u_arrmul24_fa20_13_out(h_u_arrmul24_and20_13[0], h_u_arrmul24_fa21_12_xor1[0], h_u_arrmul24_fa19_13_or0[0], h_u_arrmul24_fa20_13_xor1, h_u_arrmul24_fa20_13_or0);
  and_gate and_gate_h_u_arrmul24_and21_13(a[21], b[13], h_u_arrmul24_and21_13);
  fa fa_h_u_arrmul24_fa21_13_out(h_u_arrmul24_and21_13[0], h_u_arrmul24_fa22_12_xor1[0], h_u_arrmul24_fa20_13_or0[0], h_u_arrmul24_fa21_13_xor1, h_u_arrmul24_fa21_13_or0);
  and_gate and_gate_h_u_arrmul24_and22_13(a[22], b[13], h_u_arrmul24_and22_13);
  fa fa_h_u_arrmul24_fa22_13_out(h_u_arrmul24_and22_13[0], h_u_arrmul24_fa23_12_xor1[0], h_u_arrmul24_fa21_13_or0[0], h_u_arrmul24_fa22_13_xor1, h_u_arrmul24_fa22_13_or0);
  and_gate and_gate_h_u_arrmul24_and23_13(a[23], b[13], h_u_arrmul24_and23_13);
  fa fa_h_u_arrmul24_fa23_13_out(h_u_arrmul24_and23_13[0], h_u_arrmul24_fa23_12_or0[0], h_u_arrmul24_fa22_13_or0[0], h_u_arrmul24_fa23_13_xor1, h_u_arrmul24_fa23_13_or0);
  and_gate and_gate_h_u_arrmul24_and0_14(a[0], b[14], h_u_arrmul24_and0_14);
  ha ha_h_u_arrmul24_ha0_14_out(h_u_arrmul24_and0_14[0], h_u_arrmul24_fa1_13_xor1[0], h_u_arrmul24_ha0_14_xor0, h_u_arrmul24_ha0_14_and0);
  and_gate and_gate_h_u_arrmul24_and1_14(a[1], b[14], h_u_arrmul24_and1_14);
  fa fa_h_u_arrmul24_fa1_14_out(h_u_arrmul24_and1_14[0], h_u_arrmul24_fa2_13_xor1[0], h_u_arrmul24_ha0_14_and0[0], h_u_arrmul24_fa1_14_xor1, h_u_arrmul24_fa1_14_or0);
  and_gate and_gate_h_u_arrmul24_and2_14(a[2], b[14], h_u_arrmul24_and2_14);
  fa fa_h_u_arrmul24_fa2_14_out(h_u_arrmul24_and2_14[0], h_u_arrmul24_fa3_13_xor1[0], h_u_arrmul24_fa1_14_or0[0], h_u_arrmul24_fa2_14_xor1, h_u_arrmul24_fa2_14_or0);
  and_gate and_gate_h_u_arrmul24_and3_14(a[3], b[14], h_u_arrmul24_and3_14);
  fa fa_h_u_arrmul24_fa3_14_out(h_u_arrmul24_and3_14[0], h_u_arrmul24_fa4_13_xor1[0], h_u_arrmul24_fa2_14_or0[0], h_u_arrmul24_fa3_14_xor1, h_u_arrmul24_fa3_14_or0);
  and_gate and_gate_h_u_arrmul24_and4_14(a[4], b[14], h_u_arrmul24_and4_14);
  fa fa_h_u_arrmul24_fa4_14_out(h_u_arrmul24_and4_14[0], h_u_arrmul24_fa5_13_xor1[0], h_u_arrmul24_fa3_14_or0[0], h_u_arrmul24_fa4_14_xor1, h_u_arrmul24_fa4_14_or0);
  and_gate and_gate_h_u_arrmul24_and5_14(a[5], b[14], h_u_arrmul24_and5_14);
  fa fa_h_u_arrmul24_fa5_14_out(h_u_arrmul24_and5_14[0], h_u_arrmul24_fa6_13_xor1[0], h_u_arrmul24_fa4_14_or0[0], h_u_arrmul24_fa5_14_xor1, h_u_arrmul24_fa5_14_or0);
  and_gate and_gate_h_u_arrmul24_and6_14(a[6], b[14], h_u_arrmul24_and6_14);
  fa fa_h_u_arrmul24_fa6_14_out(h_u_arrmul24_and6_14[0], h_u_arrmul24_fa7_13_xor1[0], h_u_arrmul24_fa5_14_or0[0], h_u_arrmul24_fa6_14_xor1, h_u_arrmul24_fa6_14_or0);
  and_gate and_gate_h_u_arrmul24_and7_14(a[7], b[14], h_u_arrmul24_and7_14);
  fa fa_h_u_arrmul24_fa7_14_out(h_u_arrmul24_and7_14[0], h_u_arrmul24_fa8_13_xor1[0], h_u_arrmul24_fa6_14_or0[0], h_u_arrmul24_fa7_14_xor1, h_u_arrmul24_fa7_14_or0);
  and_gate and_gate_h_u_arrmul24_and8_14(a[8], b[14], h_u_arrmul24_and8_14);
  fa fa_h_u_arrmul24_fa8_14_out(h_u_arrmul24_and8_14[0], h_u_arrmul24_fa9_13_xor1[0], h_u_arrmul24_fa7_14_or0[0], h_u_arrmul24_fa8_14_xor1, h_u_arrmul24_fa8_14_or0);
  and_gate and_gate_h_u_arrmul24_and9_14(a[9], b[14], h_u_arrmul24_and9_14);
  fa fa_h_u_arrmul24_fa9_14_out(h_u_arrmul24_and9_14[0], h_u_arrmul24_fa10_13_xor1[0], h_u_arrmul24_fa8_14_or0[0], h_u_arrmul24_fa9_14_xor1, h_u_arrmul24_fa9_14_or0);
  and_gate and_gate_h_u_arrmul24_and10_14(a[10], b[14], h_u_arrmul24_and10_14);
  fa fa_h_u_arrmul24_fa10_14_out(h_u_arrmul24_and10_14[0], h_u_arrmul24_fa11_13_xor1[0], h_u_arrmul24_fa9_14_or0[0], h_u_arrmul24_fa10_14_xor1, h_u_arrmul24_fa10_14_or0);
  and_gate and_gate_h_u_arrmul24_and11_14(a[11], b[14], h_u_arrmul24_and11_14);
  fa fa_h_u_arrmul24_fa11_14_out(h_u_arrmul24_and11_14[0], h_u_arrmul24_fa12_13_xor1[0], h_u_arrmul24_fa10_14_or0[0], h_u_arrmul24_fa11_14_xor1, h_u_arrmul24_fa11_14_or0);
  and_gate and_gate_h_u_arrmul24_and12_14(a[12], b[14], h_u_arrmul24_and12_14);
  fa fa_h_u_arrmul24_fa12_14_out(h_u_arrmul24_and12_14[0], h_u_arrmul24_fa13_13_xor1[0], h_u_arrmul24_fa11_14_or0[0], h_u_arrmul24_fa12_14_xor1, h_u_arrmul24_fa12_14_or0);
  and_gate and_gate_h_u_arrmul24_and13_14(a[13], b[14], h_u_arrmul24_and13_14);
  fa fa_h_u_arrmul24_fa13_14_out(h_u_arrmul24_and13_14[0], h_u_arrmul24_fa14_13_xor1[0], h_u_arrmul24_fa12_14_or0[0], h_u_arrmul24_fa13_14_xor1, h_u_arrmul24_fa13_14_or0);
  and_gate and_gate_h_u_arrmul24_and14_14(a[14], b[14], h_u_arrmul24_and14_14);
  fa fa_h_u_arrmul24_fa14_14_out(h_u_arrmul24_and14_14[0], h_u_arrmul24_fa15_13_xor1[0], h_u_arrmul24_fa13_14_or0[0], h_u_arrmul24_fa14_14_xor1, h_u_arrmul24_fa14_14_or0);
  and_gate and_gate_h_u_arrmul24_and15_14(a[15], b[14], h_u_arrmul24_and15_14);
  fa fa_h_u_arrmul24_fa15_14_out(h_u_arrmul24_and15_14[0], h_u_arrmul24_fa16_13_xor1[0], h_u_arrmul24_fa14_14_or0[0], h_u_arrmul24_fa15_14_xor1, h_u_arrmul24_fa15_14_or0);
  and_gate and_gate_h_u_arrmul24_and16_14(a[16], b[14], h_u_arrmul24_and16_14);
  fa fa_h_u_arrmul24_fa16_14_out(h_u_arrmul24_and16_14[0], h_u_arrmul24_fa17_13_xor1[0], h_u_arrmul24_fa15_14_or0[0], h_u_arrmul24_fa16_14_xor1, h_u_arrmul24_fa16_14_or0);
  and_gate and_gate_h_u_arrmul24_and17_14(a[17], b[14], h_u_arrmul24_and17_14);
  fa fa_h_u_arrmul24_fa17_14_out(h_u_arrmul24_and17_14[0], h_u_arrmul24_fa18_13_xor1[0], h_u_arrmul24_fa16_14_or0[0], h_u_arrmul24_fa17_14_xor1, h_u_arrmul24_fa17_14_or0);
  and_gate and_gate_h_u_arrmul24_and18_14(a[18], b[14], h_u_arrmul24_and18_14);
  fa fa_h_u_arrmul24_fa18_14_out(h_u_arrmul24_and18_14[0], h_u_arrmul24_fa19_13_xor1[0], h_u_arrmul24_fa17_14_or0[0], h_u_arrmul24_fa18_14_xor1, h_u_arrmul24_fa18_14_or0);
  and_gate and_gate_h_u_arrmul24_and19_14(a[19], b[14], h_u_arrmul24_and19_14);
  fa fa_h_u_arrmul24_fa19_14_out(h_u_arrmul24_and19_14[0], h_u_arrmul24_fa20_13_xor1[0], h_u_arrmul24_fa18_14_or0[0], h_u_arrmul24_fa19_14_xor1, h_u_arrmul24_fa19_14_or0);
  and_gate and_gate_h_u_arrmul24_and20_14(a[20], b[14], h_u_arrmul24_and20_14);
  fa fa_h_u_arrmul24_fa20_14_out(h_u_arrmul24_and20_14[0], h_u_arrmul24_fa21_13_xor1[0], h_u_arrmul24_fa19_14_or0[0], h_u_arrmul24_fa20_14_xor1, h_u_arrmul24_fa20_14_or0);
  and_gate and_gate_h_u_arrmul24_and21_14(a[21], b[14], h_u_arrmul24_and21_14);
  fa fa_h_u_arrmul24_fa21_14_out(h_u_arrmul24_and21_14[0], h_u_arrmul24_fa22_13_xor1[0], h_u_arrmul24_fa20_14_or0[0], h_u_arrmul24_fa21_14_xor1, h_u_arrmul24_fa21_14_or0);
  and_gate and_gate_h_u_arrmul24_and22_14(a[22], b[14], h_u_arrmul24_and22_14);
  fa fa_h_u_arrmul24_fa22_14_out(h_u_arrmul24_and22_14[0], h_u_arrmul24_fa23_13_xor1[0], h_u_arrmul24_fa21_14_or0[0], h_u_arrmul24_fa22_14_xor1, h_u_arrmul24_fa22_14_or0);
  and_gate and_gate_h_u_arrmul24_and23_14(a[23], b[14], h_u_arrmul24_and23_14);
  fa fa_h_u_arrmul24_fa23_14_out(h_u_arrmul24_and23_14[0], h_u_arrmul24_fa23_13_or0[0], h_u_arrmul24_fa22_14_or0[0], h_u_arrmul24_fa23_14_xor1, h_u_arrmul24_fa23_14_or0);
  and_gate and_gate_h_u_arrmul24_and0_15(a[0], b[15], h_u_arrmul24_and0_15);
  ha ha_h_u_arrmul24_ha0_15_out(h_u_arrmul24_and0_15[0], h_u_arrmul24_fa1_14_xor1[0], h_u_arrmul24_ha0_15_xor0, h_u_arrmul24_ha0_15_and0);
  and_gate and_gate_h_u_arrmul24_and1_15(a[1], b[15], h_u_arrmul24_and1_15);
  fa fa_h_u_arrmul24_fa1_15_out(h_u_arrmul24_and1_15[0], h_u_arrmul24_fa2_14_xor1[0], h_u_arrmul24_ha0_15_and0[0], h_u_arrmul24_fa1_15_xor1, h_u_arrmul24_fa1_15_or0);
  and_gate and_gate_h_u_arrmul24_and2_15(a[2], b[15], h_u_arrmul24_and2_15);
  fa fa_h_u_arrmul24_fa2_15_out(h_u_arrmul24_and2_15[0], h_u_arrmul24_fa3_14_xor1[0], h_u_arrmul24_fa1_15_or0[0], h_u_arrmul24_fa2_15_xor1, h_u_arrmul24_fa2_15_or0);
  and_gate and_gate_h_u_arrmul24_and3_15(a[3], b[15], h_u_arrmul24_and3_15);
  fa fa_h_u_arrmul24_fa3_15_out(h_u_arrmul24_and3_15[0], h_u_arrmul24_fa4_14_xor1[0], h_u_arrmul24_fa2_15_or0[0], h_u_arrmul24_fa3_15_xor1, h_u_arrmul24_fa3_15_or0);
  and_gate and_gate_h_u_arrmul24_and4_15(a[4], b[15], h_u_arrmul24_and4_15);
  fa fa_h_u_arrmul24_fa4_15_out(h_u_arrmul24_and4_15[0], h_u_arrmul24_fa5_14_xor1[0], h_u_arrmul24_fa3_15_or0[0], h_u_arrmul24_fa4_15_xor1, h_u_arrmul24_fa4_15_or0);
  and_gate and_gate_h_u_arrmul24_and5_15(a[5], b[15], h_u_arrmul24_and5_15);
  fa fa_h_u_arrmul24_fa5_15_out(h_u_arrmul24_and5_15[0], h_u_arrmul24_fa6_14_xor1[0], h_u_arrmul24_fa4_15_or0[0], h_u_arrmul24_fa5_15_xor1, h_u_arrmul24_fa5_15_or0);
  and_gate and_gate_h_u_arrmul24_and6_15(a[6], b[15], h_u_arrmul24_and6_15);
  fa fa_h_u_arrmul24_fa6_15_out(h_u_arrmul24_and6_15[0], h_u_arrmul24_fa7_14_xor1[0], h_u_arrmul24_fa5_15_or0[0], h_u_arrmul24_fa6_15_xor1, h_u_arrmul24_fa6_15_or0);
  and_gate and_gate_h_u_arrmul24_and7_15(a[7], b[15], h_u_arrmul24_and7_15);
  fa fa_h_u_arrmul24_fa7_15_out(h_u_arrmul24_and7_15[0], h_u_arrmul24_fa8_14_xor1[0], h_u_arrmul24_fa6_15_or0[0], h_u_arrmul24_fa7_15_xor1, h_u_arrmul24_fa7_15_or0);
  and_gate and_gate_h_u_arrmul24_and8_15(a[8], b[15], h_u_arrmul24_and8_15);
  fa fa_h_u_arrmul24_fa8_15_out(h_u_arrmul24_and8_15[0], h_u_arrmul24_fa9_14_xor1[0], h_u_arrmul24_fa7_15_or0[0], h_u_arrmul24_fa8_15_xor1, h_u_arrmul24_fa8_15_or0);
  and_gate and_gate_h_u_arrmul24_and9_15(a[9], b[15], h_u_arrmul24_and9_15);
  fa fa_h_u_arrmul24_fa9_15_out(h_u_arrmul24_and9_15[0], h_u_arrmul24_fa10_14_xor1[0], h_u_arrmul24_fa8_15_or0[0], h_u_arrmul24_fa9_15_xor1, h_u_arrmul24_fa9_15_or0);
  and_gate and_gate_h_u_arrmul24_and10_15(a[10], b[15], h_u_arrmul24_and10_15);
  fa fa_h_u_arrmul24_fa10_15_out(h_u_arrmul24_and10_15[0], h_u_arrmul24_fa11_14_xor1[0], h_u_arrmul24_fa9_15_or0[0], h_u_arrmul24_fa10_15_xor1, h_u_arrmul24_fa10_15_or0);
  and_gate and_gate_h_u_arrmul24_and11_15(a[11], b[15], h_u_arrmul24_and11_15);
  fa fa_h_u_arrmul24_fa11_15_out(h_u_arrmul24_and11_15[0], h_u_arrmul24_fa12_14_xor1[0], h_u_arrmul24_fa10_15_or0[0], h_u_arrmul24_fa11_15_xor1, h_u_arrmul24_fa11_15_or0);
  and_gate and_gate_h_u_arrmul24_and12_15(a[12], b[15], h_u_arrmul24_and12_15);
  fa fa_h_u_arrmul24_fa12_15_out(h_u_arrmul24_and12_15[0], h_u_arrmul24_fa13_14_xor1[0], h_u_arrmul24_fa11_15_or0[0], h_u_arrmul24_fa12_15_xor1, h_u_arrmul24_fa12_15_or0);
  and_gate and_gate_h_u_arrmul24_and13_15(a[13], b[15], h_u_arrmul24_and13_15);
  fa fa_h_u_arrmul24_fa13_15_out(h_u_arrmul24_and13_15[0], h_u_arrmul24_fa14_14_xor1[0], h_u_arrmul24_fa12_15_or0[0], h_u_arrmul24_fa13_15_xor1, h_u_arrmul24_fa13_15_or0);
  and_gate and_gate_h_u_arrmul24_and14_15(a[14], b[15], h_u_arrmul24_and14_15);
  fa fa_h_u_arrmul24_fa14_15_out(h_u_arrmul24_and14_15[0], h_u_arrmul24_fa15_14_xor1[0], h_u_arrmul24_fa13_15_or0[0], h_u_arrmul24_fa14_15_xor1, h_u_arrmul24_fa14_15_or0);
  and_gate and_gate_h_u_arrmul24_and15_15(a[15], b[15], h_u_arrmul24_and15_15);
  fa fa_h_u_arrmul24_fa15_15_out(h_u_arrmul24_and15_15[0], h_u_arrmul24_fa16_14_xor1[0], h_u_arrmul24_fa14_15_or0[0], h_u_arrmul24_fa15_15_xor1, h_u_arrmul24_fa15_15_or0);
  and_gate and_gate_h_u_arrmul24_and16_15(a[16], b[15], h_u_arrmul24_and16_15);
  fa fa_h_u_arrmul24_fa16_15_out(h_u_arrmul24_and16_15[0], h_u_arrmul24_fa17_14_xor1[0], h_u_arrmul24_fa15_15_or0[0], h_u_arrmul24_fa16_15_xor1, h_u_arrmul24_fa16_15_or0);
  and_gate and_gate_h_u_arrmul24_and17_15(a[17], b[15], h_u_arrmul24_and17_15);
  fa fa_h_u_arrmul24_fa17_15_out(h_u_arrmul24_and17_15[0], h_u_arrmul24_fa18_14_xor1[0], h_u_arrmul24_fa16_15_or0[0], h_u_arrmul24_fa17_15_xor1, h_u_arrmul24_fa17_15_or0);
  and_gate and_gate_h_u_arrmul24_and18_15(a[18], b[15], h_u_arrmul24_and18_15);
  fa fa_h_u_arrmul24_fa18_15_out(h_u_arrmul24_and18_15[0], h_u_arrmul24_fa19_14_xor1[0], h_u_arrmul24_fa17_15_or0[0], h_u_arrmul24_fa18_15_xor1, h_u_arrmul24_fa18_15_or0);
  and_gate and_gate_h_u_arrmul24_and19_15(a[19], b[15], h_u_arrmul24_and19_15);
  fa fa_h_u_arrmul24_fa19_15_out(h_u_arrmul24_and19_15[0], h_u_arrmul24_fa20_14_xor1[0], h_u_arrmul24_fa18_15_or0[0], h_u_arrmul24_fa19_15_xor1, h_u_arrmul24_fa19_15_or0);
  and_gate and_gate_h_u_arrmul24_and20_15(a[20], b[15], h_u_arrmul24_and20_15);
  fa fa_h_u_arrmul24_fa20_15_out(h_u_arrmul24_and20_15[0], h_u_arrmul24_fa21_14_xor1[0], h_u_arrmul24_fa19_15_or0[0], h_u_arrmul24_fa20_15_xor1, h_u_arrmul24_fa20_15_or0);
  and_gate and_gate_h_u_arrmul24_and21_15(a[21], b[15], h_u_arrmul24_and21_15);
  fa fa_h_u_arrmul24_fa21_15_out(h_u_arrmul24_and21_15[0], h_u_arrmul24_fa22_14_xor1[0], h_u_arrmul24_fa20_15_or0[0], h_u_arrmul24_fa21_15_xor1, h_u_arrmul24_fa21_15_or0);
  and_gate and_gate_h_u_arrmul24_and22_15(a[22], b[15], h_u_arrmul24_and22_15);
  fa fa_h_u_arrmul24_fa22_15_out(h_u_arrmul24_and22_15[0], h_u_arrmul24_fa23_14_xor1[0], h_u_arrmul24_fa21_15_or0[0], h_u_arrmul24_fa22_15_xor1, h_u_arrmul24_fa22_15_or0);
  and_gate and_gate_h_u_arrmul24_and23_15(a[23], b[15], h_u_arrmul24_and23_15);
  fa fa_h_u_arrmul24_fa23_15_out(h_u_arrmul24_and23_15[0], h_u_arrmul24_fa23_14_or0[0], h_u_arrmul24_fa22_15_or0[0], h_u_arrmul24_fa23_15_xor1, h_u_arrmul24_fa23_15_or0);
  and_gate and_gate_h_u_arrmul24_and0_16(a[0], b[16], h_u_arrmul24_and0_16);
  ha ha_h_u_arrmul24_ha0_16_out(h_u_arrmul24_and0_16[0], h_u_arrmul24_fa1_15_xor1[0], h_u_arrmul24_ha0_16_xor0, h_u_arrmul24_ha0_16_and0);
  and_gate and_gate_h_u_arrmul24_and1_16(a[1], b[16], h_u_arrmul24_and1_16);
  fa fa_h_u_arrmul24_fa1_16_out(h_u_arrmul24_and1_16[0], h_u_arrmul24_fa2_15_xor1[0], h_u_arrmul24_ha0_16_and0[0], h_u_arrmul24_fa1_16_xor1, h_u_arrmul24_fa1_16_or0);
  and_gate and_gate_h_u_arrmul24_and2_16(a[2], b[16], h_u_arrmul24_and2_16);
  fa fa_h_u_arrmul24_fa2_16_out(h_u_arrmul24_and2_16[0], h_u_arrmul24_fa3_15_xor1[0], h_u_arrmul24_fa1_16_or0[0], h_u_arrmul24_fa2_16_xor1, h_u_arrmul24_fa2_16_or0);
  and_gate and_gate_h_u_arrmul24_and3_16(a[3], b[16], h_u_arrmul24_and3_16);
  fa fa_h_u_arrmul24_fa3_16_out(h_u_arrmul24_and3_16[0], h_u_arrmul24_fa4_15_xor1[0], h_u_arrmul24_fa2_16_or0[0], h_u_arrmul24_fa3_16_xor1, h_u_arrmul24_fa3_16_or0);
  and_gate and_gate_h_u_arrmul24_and4_16(a[4], b[16], h_u_arrmul24_and4_16);
  fa fa_h_u_arrmul24_fa4_16_out(h_u_arrmul24_and4_16[0], h_u_arrmul24_fa5_15_xor1[0], h_u_arrmul24_fa3_16_or0[0], h_u_arrmul24_fa4_16_xor1, h_u_arrmul24_fa4_16_or0);
  and_gate and_gate_h_u_arrmul24_and5_16(a[5], b[16], h_u_arrmul24_and5_16);
  fa fa_h_u_arrmul24_fa5_16_out(h_u_arrmul24_and5_16[0], h_u_arrmul24_fa6_15_xor1[0], h_u_arrmul24_fa4_16_or0[0], h_u_arrmul24_fa5_16_xor1, h_u_arrmul24_fa5_16_or0);
  and_gate and_gate_h_u_arrmul24_and6_16(a[6], b[16], h_u_arrmul24_and6_16);
  fa fa_h_u_arrmul24_fa6_16_out(h_u_arrmul24_and6_16[0], h_u_arrmul24_fa7_15_xor1[0], h_u_arrmul24_fa5_16_or0[0], h_u_arrmul24_fa6_16_xor1, h_u_arrmul24_fa6_16_or0);
  and_gate and_gate_h_u_arrmul24_and7_16(a[7], b[16], h_u_arrmul24_and7_16);
  fa fa_h_u_arrmul24_fa7_16_out(h_u_arrmul24_and7_16[0], h_u_arrmul24_fa8_15_xor1[0], h_u_arrmul24_fa6_16_or0[0], h_u_arrmul24_fa7_16_xor1, h_u_arrmul24_fa7_16_or0);
  and_gate and_gate_h_u_arrmul24_and8_16(a[8], b[16], h_u_arrmul24_and8_16);
  fa fa_h_u_arrmul24_fa8_16_out(h_u_arrmul24_and8_16[0], h_u_arrmul24_fa9_15_xor1[0], h_u_arrmul24_fa7_16_or0[0], h_u_arrmul24_fa8_16_xor1, h_u_arrmul24_fa8_16_or0);
  and_gate and_gate_h_u_arrmul24_and9_16(a[9], b[16], h_u_arrmul24_and9_16);
  fa fa_h_u_arrmul24_fa9_16_out(h_u_arrmul24_and9_16[0], h_u_arrmul24_fa10_15_xor1[0], h_u_arrmul24_fa8_16_or0[0], h_u_arrmul24_fa9_16_xor1, h_u_arrmul24_fa9_16_or0);
  and_gate and_gate_h_u_arrmul24_and10_16(a[10], b[16], h_u_arrmul24_and10_16);
  fa fa_h_u_arrmul24_fa10_16_out(h_u_arrmul24_and10_16[0], h_u_arrmul24_fa11_15_xor1[0], h_u_arrmul24_fa9_16_or0[0], h_u_arrmul24_fa10_16_xor1, h_u_arrmul24_fa10_16_or0);
  and_gate and_gate_h_u_arrmul24_and11_16(a[11], b[16], h_u_arrmul24_and11_16);
  fa fa_h_u_arrmul24_fa11_16_out(h_u_arrmul24_and11_16[0], h_u_arrmul24_fa12_15_xor1[0], h_u_arrmul24_fa10_16_or0[0], h_u_arrmul24_fa11_16_xor1, h_u_arrmul24_fa11_16_or0);
  and_gate and_gate_h_u_arrmul24_and12_16(a[12], b[16], h_u_arrmul24_and12_16);
  fa fa_h_u_arrmul24_fa12_16_out(h_u_arrmul24_and12_16[0], h_u_arrmul24_fa13_15_xor1[0], h_u_arrmul24_fa11_16_or0[0], h_u_arrmul24_fa12_16_xor1, h_u_arrmul24_fa12_16_or0);
  and_gate and_gate_h_u_arrmul24_and13_16(a[13], b[16], h_u_arrmul24_and13_16);
  fa fa_h_u_arrmul24_fa13_16_out(h_u_arrmul24_and13_16[0], h_u_arrmul24_fa14_15_xor1[0], h_u_arrmul24_fa12_16_or0[0], h_u_arrmul24_fa13_16_xor1, h_u_arrmul24_fa13_16_or0);
  and_gate and_gate_h_u_arrmul24_and14_16(a[14], b[16], h_u_arrmul24_and14_16);
  fa fa_h_u_arrmul24_fa14_16_out(h_u_arrmul24_and14_16[0], h_u_arrmul24_fa15_15_xor1[0], h_u_arrmul24_fa13_16_or0[0], h_u_arrmul24_fa14_16_xor1, h_u_arrmul24_fa14_16_or0);
  and_gate and_gate_h_u_arrmul24_and15_16(a[15], b[16], h_u_arrmul24_and15_16);
  fa fa_h_u_arrmul24_fa15_16_out(h_u_arrmul24_and15_16[0], h_u_arrmul24_fa16_15_xor1[0], h_u_arrmul24_fa14_16_or0[0], h_u_arrmul24_fa15_16_xor1, h_u_arrmul24_fa15_16_or0);
  and_gate and_gate_h_u_arrmul24_and16_16(a[16], b[16], h_u_arrmul24_and16_16);
  fa fa_h_u_arrmul24_fa16_16_out(h_u_arrmul24_and16_16[0], h_u_arrmul24_fa17_15_xor1[0], h_u_arrmul24_fa15_16_or0[0], h_u_arrmul24_fa16_16_xor1, h_u_arrmul24_fa16_16_or0);
  and_gate and_gate_h_u_arrmul24_and17_16(a[17], b[16], h_u_arrmul24_and17_16);
  fa fa_h_u_arrmul24_fa17_16_out(h_u_arrmul24_and17_16[0], h_u_arrmul24_fa18_15_xor1[0], h_u_arrmul24_fa16_16_or0[0], h_u_arrmul24_fa17_16_xor1, h_u_arrmul24_fa17_16_or0);
  and_gate and_gate_h_u_arrmul24_and18_16(a[18], b[16], h_u_arrmul24_and18_16);
  fa fa_h_u_arrmul24_fa18_16_out(h_u_arrmul24_and18_16[0], h_u_arrmul24_fa19_15_xor1[0], h_u_arrmul24_fa17_16_or0[0], h_u_arrmul24_fa18_16_xor1, h_u_arrmul24_fa18_16_or0);
  and_gate and_gate_h_u_arrmul24_and19_16(a[19], b[16], h_u_arrmul24_and19_16);
  fa fa_h_u_arrmul24_fa19_16_out(h_u_arrmul24_and19_16[0], h_u_arrmul24_fa20_15_xor1[0], h_u_arrmul24_fa18_16_or0[0], h_u_arrmul24_fa19_16_xor1, h_u_arrmul24_fa19_16_or0);
  and_gate and_gate_h_u_arrmul24_and20_16(a[20], b[16], h_u_arrmul24_and20_16);
  fa fa_h_u_arrmul24_fa20_16_out(h_u_arrmul24_and20_16[0], h_u_arrmul24_fa21_15_xor1[0], h_u_arrmul24_fa19_16_or0[0], h_u_arrmul24_fa20_16_xor1, h_u_arrmul24_fa20_16_or0);
  and_gate and_gate_h_u_arrmul24_and21_16(a[21], b[16], h_u_arrmul24_and21_16);
  fa fa_h_u_arrmul24_fa21_16_out(h_u_arrmul24_and21_16[0], h_u_arrmul24_fa22_15_xor1[0], h_u_arrmul24_fa20_16_or0[0], h_u_arrmul24_fa21_16_xor1, h_u_arrmul24_fa21_16_or0);
  and_gate and_gate_h_u_arrmul24_and22_16(a[22], b[16], h_u_arrmul24_and22_16);
  fa fa_h_u_arrmul24_fa22_16_out(h_u_arrmul24_and22_16[0], h_u_arrmul24_fa23_15_xor1[0], h_u_arrmul24_fa21_16_or0[0], h_u_arrmul24_fa22_16_xor1, h_u_arrmul24_fa22_16_or0);
  and_gate and_gate_h_u_arrmul24_and23_16(a[23], b[16], h_u_arrmul24_and23_16);
  fa fa_h_u_arrmul24_fa23_16_out(h_u_arrmul24_and23_16[0], h_u_arrmul24_fa23_15_or0[0], h_u_arrmul24_fa22_16_or0[0], h_u_arrmul24_fa23_16_xor1, h_u_arrmul24_fa23_16_or0);
  and_gate and_gate_h_u_arrmul24_and0_17(a[0], b[17], h_u_arrmul24_and0_17);
  ha ha_h_u_arrmul24_ha0_17_out(h_u_arrmul24_and0_17[0], h_u_arrmul24_fa1_16_xor1[0], h_u_arrmul24_ha0_17_xor0, h_u_arrmul24_ha0_17_and0);
  and_gate and_gate_h_u_arrmul24_and1_17(a[1], b[17], h_u_arrmul24_and1_17);
  fa fa_h_u_arrmul24_fa1_17_out(h_u_arrmul24_and1_17[0], h_u_arrmul24_fa2_16_xor1[0], h_u_arrmul24_ha0_17_and0[0], h_u_arrmul24_fa1_17_xor1, h_u_arrmul24_fa1_17_or0);
  and_gate and_gate_h_u_arrmul24_and2_17(a[2], b[17], h_u_arrmul24_and2_17);
  fa fa_h_u_arrmul24_fa2_17_out(h_u_arrmul24_and2_17[0], h_u_arrmul24_fa3_16_xor1[0], h_u_arrmul24_fa1_17_or0[0], h_u_arrmul24_fa2_17_xor1, h_u_arrmul24_fa2_17_or0);
  and_gate and_gate_h_u_arrmul24_and3_17(a[3], b[17], h_u_arrmul24_and3_17);
  fa fa_h_u_arrmul24_fa3_17_out(h_u_arrmul24_and3_17[0], h_u_arrmul24_fa4_16_xor1[0], h_u_arrmul24_fa2_17_or0[0], h_u_arrmul24_fa3_17_xor1, h_u_arrmul24_fa3_17_or0);
  and_gate and_gate_h_u_arrmul24_and4_17(a[4], b[17], h_u_arrmul24_and4_17);
  fa fa_h_u_arrmul24_fa4_17_out(h_u_arrmul24_and4_17[0], h_u_arrmul24_fa5_16_xor1[0], h_u_arrmul24_fa3_17_or0[0], h_u_arrmul24_fa4_17_xor1, h_u_arrmul24_fa4_17_or0);
  and_gate and_gate_h_u_arrmul24_and5_17(a[5], b[17], h_u_arrmul24_and5_17);
  fa fa_h_u_arrmul24_fa5_17_out(h_u_arrmul24_and5_17[0], h_u_arrmul24_fa6_16_xor1[0], h_u_arrmul24_fa4_17_or0[0], h_u_arrmul24_fa5_17_xor1, h_u_arrmul24_fa5_17_or0);
  and_gate and_gate_h_u_arrmul24_and6_17(a[6], b[17], h_u_arrmul24_and6_17);
  fa fa_h_u_arrmul24_fa6_17_out(h_u_arrmul24_and6_17[0], h_u_arrmul24_fa7_16_xor1[0], h_u_arrmul24_fa5_17_or0[0], h_u_arrmul24_fa6_17_xor1, h_u_arrmul24_fa6_17_or0);
  and_gate and_gate_h_u_arrmul24_and7_17(a[7], b[17], h_u_arrmul24_and7_17);
  fa fa_h_u_arrmul24_fa7_17_out(h_u_arrmul24_and7_17[0], h_u_arrmul24_fa8_16_xor1[0], h_u_arrmul24_fa6_17_or0[0], h_u_arrmul24_fa7_17_xor1, h_u_arrmul24_fa7_17_or0);
  and_gate and_gate_h_u_arrmul24_and8_17(a[8], b[17], h_u_arrmul24_and8_17);
  fa fa_h_u_arrmul24_fa8_17_out(h_u_arrmul24_and8_17[0], h_u_arrmul24_fa9_16_xor1[0], h_u_arrmul24_fa7_17_or0[0], h_u_arrmul24_fa8_17_xor1, h_u_arrmul24_fa8_17_or0);
  and_gate and_gate_h_u_arrmul24_and9_17(a[9], b[17], h_u_arrmul24_and9_17);
  fa fa_h_u_arrmul24_fa9_17_out(h_u_arrmul24_and9_17[0], h_u_arrmul24_fa10_16_xor1[0], h_u_arrmul24_fa8_17_or0[0], h_u_arrmul24_fa9_17_xor1, h_u_arrmul24_fa9_17_or0);
  and_gate and_gate_h_u_arrmul24_and10_17(a[10], b[17], h_u_arrmul24_and10_17);
  fa fa_h_u_arrmul24_fa10_17_out(h_u_arrmul24_and10_17[0], h_u_arrmul24_fa11_16_xor1[0], h_u_arrmul24_fa9_17_or0[0], h_u_arrmul24_fa10_17_xor1, h_u_arrmul24_fa10_17_or0);
  and_gate and_gate_h_u_arrmul24_and11_17(a[11], b[17], h_u_arrmul24_and11_17);
  fa fa_h_u_arrmul24_fa11_17_out(h_u_arrmul24_and11_17[0], h_u_arrmul24_fa12_16_xor1[0], h_u_arrmul24_fa10_17_or0[0], h_u_arrmul24_fa11_17_xor1, h_u_arrmul24_fa11_17_or0);
  and_gate and_gate_h_u_arrmul24_and12_17(a[12], b[17], h_u_arrmul24_and12_17);
  fa fa_h_u_arrmul24_fa12_17_out(h_u_arrmul24_and12_17[0], h_u_arrmul24_fa13_16_xor1[0], h_u_arrmul24_fa11_17_or0[0], h_u_arrmul24_fa12_17_xor1, h_u_arrmul24_fa12_17_or0);
  and_gate and_gate_h_u_arrmul24_and13_17(a[13], b[17], h_u_arrmul24_and13_17);
  fa fa_h_u_arrmul24_fa13_17_out(h_u_arrmul24_and13_17[0], h_u_arrmul24_fa14_16_xor1[0], h_u_arrmul24_fa12_17_or0[0], h_u_arrmul24_fa13_17_xor1, h_u_arrmul24_fa13_17_or0);
  and_gate and_gate_h_u_arrmul24_and14_17(a[14], b[17], h_u_arrmul24_and14_17);
  fa fa_h_u_arrmul24_fa14_17_out(h_u_arrmul24_and14_17[0], h_u_arrmul24_fa15_16_xor1[0], h_u_arrmul24_fa13_17_or0[0], h_u_arrmul24_fa14_17_xor1, h_u_arrmul24_fa14_17_or0);
  and_gate and_gate_h_u_arrmul24_and15_17(a[15], b[17], h_u_arrmul24_and15_17);
  fa fa_h_u_arrmul24_fa15_17_out(h_u_arrmul24_and15_17[0], h_u_arrmul24_fa16_16_xor1[0], h_u_arrmul24_fa14_17_or0[0], h_u_arrmul24_fa15_17_xor1, h_u_arrmul24_fa15_17_or0);
  and_gate and_gate_h_u_arrmul24_and16_17(a[16], b[17], h_u_arrmul24_and16_17);
  fa fa_h_u_arrmul24_fa16_17_out(h_u_arrmul24_and16_17[0], h_u_arrmul24_fa17_16_xor1[0], h_u_arrmul24_fa15_17_or0[0], h_u_arrmul24_fa16_17_xor1, h_u_arrmul24_fa16_17_or0);
  and_gate and_gate_h_u_arrmul24_and17_17(a[17], b[17], h_u_arrmul24_and17_17);
  fa fa_h_u_arrmul24_fa17_17_out(h_u_arrmul24_and17_17[0], h_u_arrmul24_fa18_16_xor1[0], h_u_arrmul24_fa16_17_or0[0], h_u_arrmul24_fa17_17_xor1, h_u_arrmul24_fa17_17_or0);
  and_gate and_gate_h_u_arrmul24_and18_17(a[18], b[17], h_u_arrmul24_and18_17);
  fa fa_h_u_arrmul24_fa18_17_out(h_u_arrmul24_and18_17[0], h_u_arrmul24_fa19_16_xor1[0], h_u_arrmul24_fa17_17_or0[0], h_u_arrmul24_fa18_17_xor1, h_u_arrmul24_fa18_17_or0);
  and_gate and_gate_h_u_arrmul24_and19_17(a[19], b[17], h_u_arrmul24_and19_17);
  fa fa_h_u_arrmul24_fa19_17_out(h_u_arrmul24_and19_17[0], h_u_arrmul24_fa20_16_xor1[0], h_u_arrmul24_fa18_17_or0[0], h_u_arrmul24_fa19_17_xor1, h_u_arrmul24_fa19_17_or0);
  and_gate and_gate_h_u_arrmul24_and20_17(a[20], b[17], h_u_arrmul24_and20_17);
  fa fa_h_u_arrmul24_fa20_17_out(h_u_arrmul24_and20_17[0], h_u_arrmul24_fa21_16_xor1[0], h_u_arrmul24_fa19_17_or0[0], h_u_arrmul24_fa20_17_xor1, h_u_arrmul24_fa20_17_or0);
  and_gate and_gate_h_u_arrmul24_and21_17(a[21], b[17], h_u_arrmul24_and21_17);
  fa fa_h_u_arrmul24_fa21_17_out(h_u_arrmul24_and21_17[0], h_u_arrmul24_fa22_16_xor1[0], h_u_arrmul24_fa20_17_or0[0], h_u_arrmul24_fa21_17_xor1, h_u_arrmul24_fa21_17_or0);
  and_gate and_gate_h_u_arrmul24_and22_17(a[22], b[17], h_u_arrmul24_and22_17);
  fa fa_h_u_arrmul24_fa22_17_out(h_u_arrmul24_and22_17[0], h_u_arrmul24_fa23_16_xor1[0], h_u_arrmul24_fa21_17_or0[0], h_u_arrmul24_fa22_17_xor1, h_u_arrmul24_fa22_17_or0);
  and_gate and_gate_h_u_arrmul24_and23_17(a[23], b[17], h_u_arrmul24_and23_17);
  fa fa_h_u_arrmul24_fa23_17_out(h_u_arrmul24_and23_17[0], h_u_arrmul24_fa23_16_or0[0], h_u_arrmul24_fa22_17_or0[0], h_u_arrmul24_fa23_17_xor1, h_u_arrmul24_fa23_17_or0);
  and_gate and_gate_h_u_arrmul24_and0_18(a[0], b[18], h_u_arrmul24_and0_18);
  ha ha_h_u_arrmul24_ha0_18_out(h_u_arrmul24_and0_18[0], h_u_arrmul24_fa1_17_xor1[0], h_u_arrmul24_ha0_18_xor0, h_u_arrmul24_ha0_18_and0);
  and_gate and_gate_h_u_arrmul24_and1_18(a[1], b[18], h_u_arrmul24_and1_18);
  fa fa_h_u_arrmul24_fa1_18_out(h_u_arrmul24_and1_18[0], h_u_arrmul24_fa2_17_xor1[0], h_u_arrmul24_ha0_18_and0[0], h_u_arrmul24_fa1_18_xor1, h_u_arrmul24_fa1_18_or0);
  and_gate and_gate_h_u_arrmul24_and2_18(a[2], b[18], h_u_arrmul24_and2_18);
  fa fa_h_u_arrmul24_fa2_18_out(h_u_arrmul24_and2_18[0], h_u_arrmul24_fa3_17_xor1[0], h_u_arrmul24_fa1_18_or0[0], h_u_arrmul24_fa2_18_xor1, h_u_arrmul24_fa2_18_or0);
  and_gate and_gate_h_u_arrmul24_and3_18(a[3], b[18], h_u_arrmul24_and3_18);
  fa fa_h_u_arrmul24_fa3_18_out(h_u_arrmul24_and3_18[0], h_u_arrmul24_fa4_17_xor1[0], h_u_arrmul24_fa2_18_or0[0], h_u_arrmul24_fa3_18_xor1, h_u_arrmul24_fa3_18_or0);
  and_gate and_gate_h_u_arrmul24_and4_18(a[4], b[18], h_u_arrmul24_and4_18);
  fa fa_h_u_arrmul24_fa4_18_out(h_u_arrmul24_and4_18[0], h_u_arrmul24_fa5_17_xor1[0], h_u_arrmul24_fa3_18_or0[0], h_u_arrmul24_fa4_18_xor1, h_u_arrmul24_fa4_18_or0);
  and_gate and_gate_h_u_arrmul24_and5_18(a[5], b[18], h_u_arrmul24_and5_18);
  fa fa_h_u_arrmul24_fa5_18_out(h_u_arrmul24_and5_18[0], h_u_arrmul24_fa6_17_xor1[0], h_u_arrmul24_fa4_18_or0[0], h_u_arrmul24_fa5_18_xor1, h_u_arrmul24_fa5_18_or0);
  and_gate and_gate_h_u_arrmul24_and6_18(a[6], b[18], h_u_arrmul24_and6_18);
  fa fa_h_u_arrmul24_fa6_18_out(h_u_arrmul24_and6_18[0], h_u_arrmul24_fa7_17_xor1[0], h_u_arrmul24_fa5_18_or0[0], h_u_arrmul24_fa6_18_xor1, h_u_arrmul24_fa6_18_or0);
  and_gate and_gate_h_u_arrmul24_and7_18(a[7], b[18], h_u_arrmul24_and7_18);
  fa fa_h_u_arrmul24_fa7_18_out(h_u_arrmul24_and7_18[0], h_u_arrmul24_fa8_17_xor1[0], h_u_arrmul24_fa6_18_or0[0], h_u_arrmul24_fa7_18_xor1, h_u_arrmul24_fa7_18_or0);
  and_gate and_gate_h_u_arrmul24_and8_18(a[8], b[18], h_u_arrmul24_and8_18);
  fa fa_h_u_arrmul24_fa8_18_out(h_u_arrmul24_and8_18[0], h_u_arrmul24_fa9_17_xor1[0], h_u_arrmul24_fa7_18_or0[0], h_u_arrmul24_fa8_18_xor1, h_u_arrmul24_fa8_18_or0);
  and_gate and_gate_h_u_arrmul24_and9_18(a[9], b[18], h_u_arrmul24_and9_18);
  fa fa_h_u_arrmul24_fa9_18_out(h_u_arrmul24_and9_18[0], h_u_arrmul24_fa10_17_xor1[0], h_u_arrmul24_fa8_18_or0[0], h_u_arrmul24_fa9_18_xor1, h_u_arrmul24_fa9_18_or0);
  and_gate and_gate_h_u_arrmul24_and10_18(a[10], b[18], h_u_arrmul24_and10_18);
  fa fa_h_u_arrmul24_fa10_18_out(h_u_arrmul24_and10_18[0], h_u_arrmul24_fa11_17_xor1[0], h_u_arrmul24_fa9_18_or0[0], h_u_arrmul24_fa10_18_xor1, h_u_arrmul24_fa10_18_or0);
  and_gate and_gate_h_u_arrmul24_and11_18(a[11], b[18], h_u_arrmul24_and11_18);
  fa fa_h_u_arrmul24_fa11_18_out(h_u_arrmul24_and11_18[0], h_u_arrmul24_fa12_17_xor1[0], h_u_arrmul24_fa10_18_or0[0], h_u_arrmul24_fa11_18_xor1, h_u_arrmul24_fa11_18_or0);
  and_gate and_gate_h_u_arrmul24_and12_18(a[12], b[18], h_u_arrmul24_and12_18);
  fa fa_h_u_arrmul24_fa12_18_out(h_u_arrmul24_and12_18[0], h_u_arrmul24_fa13_17_xor1[0], h_u_arrmul24_fa11_18_or0[0], h_u_arrmul24_fa12_18_xor1, h_u_arrmul24_fa12_18_or0);
  and_gate and_gate_h_u_arrmul24_and13_18(a[13], b[18], h_u_arrmul24_and13_18);
  fa fa_h_u_arrmul24_fa13_18_out(h_u_arrmul24_and13_18[0], h_u_arrmul24_fa14_17_xor1[0], h_u_arrmul24_fa12_18_or0[0], h_u_arrmul24_fa13_18_xor1, h_u_arrmul24_fa13_18_or0);
  and_gate and_gate_h_u_arrmul24_and14_18(a[14], b[18], h_u_arrmul24_and14_18);
  fa fa_h_u_arrmul24_fa14_18_out(h_u_arrmul24_and14_18[0], h_u_arrmul24_fa15_17_xor1[0], h_u_arrmul24_fa13_18_or0[0], h_u_arrmul24_fa14_18_xor1, h_u_arrmul24_fa14_18_or0);
  and_gate and_gate_h_u_arrmul24_and15_18(a[15], b[18], h_u_arrmul24_and15_18);
  fa fa_h_u_arrmul24_fa15_18_out(h_u_arrmul24_and15_18[0], h_u_arrmul24_fa16_17_xor1[0], h_u_arrmul24_fa14_18_or0[0], h_u_arrmul24_fa15_18_xor1, h_u_arrmul24_fa15_18_or0);
  and_gate and_gate_h_u_arrmul24_and16_18(a[16], b[18], h_u_arrmul24_and16_18);
  fa fa_h_u_arrmul24_fa16_18_out(h_u_arrmul24_and16_18[0], h_u_arrmul24_fa17_17_xor1[0], h_u_arrmul24_fa15_18_or0[0], h_u_arrmul24_fa16_18_xor1, h_u_arrmul24_fa16_18_or0);
  and_gate and_gate_h_u_arrmul24_and17_18(a[17], b[18], h_u_arrmul24_and17_18);
  fa fa_h_u_arrmul24_fa17_18_out(h_u_arrmul24_and17_18[0], h_u_arrmul24_fa18_17_xor1[0], h_u_arrmul24_fa16_18_or0[0], h_u_arrmul24_fa17_18_xor1, h_u_arrmul24_fa17_18_or0);
  and_gate and_gate_h_u_arrmul24_and18_18(a[18], b[18], h_u_arrmul24_and18_18);
  fa fa_h_u_arrmul24_fa18_18_out(h_u_arrmul24_and18_18[0], h_u_arrmul24_fa19_17_xor1[0], h_u_arrmul24_fa17_18_or0[0], h_u_arrmul24_fa18_18_xor1, h_u_arrmul24_fa18_18_or0);
  and_gate and_gate_h_u_arrmul24_and19_18(a[19], b[18], h_u_arrmul24_and19_18);
  fa fa_h_u_arrmul24_fa19_18_out(h_u_arrmul24_and19_18[0], h_u_arrmul24_fa20_17_xor1[0], h_u_arrmul24_fa18_18_or0[0], h_u_arrmul24_fa19_18_xor1, h_u_arrmul24_fa19_18_or0);
  and_gate and_gate_h_u_arrmul24_and20_18(a[20], b[18], h_u_arrmul24_and20_18);
  fa fa_h_u_arrmul24_fa20_18_out(h_u_arrmul24_and20_18[0], h_u_arrmul24_fa21_17_xor1[0], h_u_arrmul24_fa19_18_or0[0], h_u_arrmul24_fa20_18_xor1, h_u_arrmul24_fa20_18_or0);
  and_gate and_gate_h_u_arrmul24_and21_18(a[21], b[18], h_u_arrmul24_and21_18);
  fa fa_h_u_arrmul24_fa21_18_out(h_u_arrmul24_and21_18[0], h_u_arrmul24_fa22_17_xor1[0], h_u_arrmul24_fa20_18_or0[0], h_u_arrmul24_fa21_18_xor1, h_u_arrmul24_fa21_18_or0);
  and_gate and_gate_h_u_arrmul24_and22_18(a[22], b[18], h_u_arrmul24_and22_18);
  fa fa_h_u_arrmul24_fa22_18_out(h_u_arrmul24_and22_18[0], h_u_arrmul24_fa23_17_xor1[0], h_u_arrmul24_fa21_18_or0[0], h_u_arrmul24_fa22_18_xor1, h_u_arrmul24_fa22_18_or0);
  and_gate and_gate_h_u_arrmul24_and23_18(a[23], b[18], h_u_arrmul24_and23_18);
  fa fa_h_u_arrmul24_fa23_18_out(h_u_arrmul24_and23_18[0], h_u_arrmul24_fa23_17_or0[0], h_u_arrmul24_fa22_18_or0[0], h_u_arrmul24_fa23_18_xor1, h_u_arrmul24_fa23_18_or0);
  and_gate and_gate_h_u_arrmul24_and0_19(a[0], b[19], h_u_arrmul24_and0_19);
  ha ha_h_u_arrmul24_ha0_19_out(h_u_arrmul24_and0_19[0], h_u_arrmul24_fa1_18_xor1[0], h_u_arrmul24_ha0_19_xor0, h_u_arrmul24_ha0_19_and0);
  and_gate and_gate_h_u_arrmul24_and1_19(a[1], b[19], h_u_arrmul24_and1_19);
  fa fa_h_u_arrmul24_fa1_19_out(h_u_arrmul24_and1_19[0], h_u_arrmul24_fa2_18_xor1[0], h_u_arrmul24_ha0_19_and0[0], h_u_arrmul24_fa1_19_xor1, h_u_arrmul24_fa1_19_or0);
  and_gate and_gate_h_u_arrmul24_and2_19(a[2], b[19], h_u_arrmul24_and2_19);
  fa fa_h_u_arrmul24_fa2_19_out(h_u_arrmul24_and2_19[0], h_u_arrmul24_fa3_18_xor1[0], h_u_arrmul24_fa1_19_or0[0], h_u_arrmul24_fa2_19_xor1, h_u_arrmul24_fa2_19_or0);
  and_gate and_gate_h_u_arrmul24_and3_19(a[3], b[19], h_u_arrmul24_and3_19);
  fa fa_h_u_arrmul24_fa3_19_out(h_u_arrmul24_and3_19[0], h_u_arrmul24_fa4_18_xor1[0], h_u_arrmul24_fa2_19_or0[0], h_u_arrmul24_fa3_19_xor1, h_u_arrmul24_fa3_19_or0);
  and_gate and_gate_h_u_arrmul24_and4_19(a[4], b[19], h_u_arrmul24_and4_19);
  fa fa_h_u_arrmul24_fa4_19_out(h_u_arrmul24_and4_19[0], h_u_arrmul24_fa5_18_xor1[0], h_u_arrmul24_fa3_19_or0[0], h_u_arrmul24_fa4_19_xor1, h_u_arrmul24_fa4_19_or0);
  and_gate and_gate_h_u_arrmul24_and5_19(a[5], b[19], h_u_arrmul24_and5_19);
  fa fa_h_u_arrmul24_fa5_19_out(h_u_arrmul24_and5_19[0], h_u_arrmul24_fa6_18_xor1[0], h_u_arrmul24_fa4_19_or0[0], h_u_arrmul24_fa5_19_xor1, h_u_arrmul24_fa5_19_or0);
  and_gate and_gate_h_u_arrmul24_and6_19(a[6], b[19], h_u_arrmul24_and6_19);
  fa fa_h_u_arrmul24_fa6_19_out(h_u_arrmul24_and6_19[0], h_u_arrmul24_fa7_18_xor1[0], h_u_arrmul24_fa5_19_or0[0], h_u_arrmul24_fa6_19_xor1, h_u_arrmul24_fa6_19_or0);
  and_gate and_gate_h_u_arrmul24_and7_19(a[7], b[19], h_u_arrmul24_and7_19);
  fa fa_h_u_arrmul24_fa7_19_out(h_u_arrmul24_and7_19[0], h_u_arrmul24_fa8_18_xor1[0], h_u_arrmul24_fa6_19_or0[0], h_u_arrmul24_fa7_19_xor1, h_u_arrmul24_fa7_19_or0);
  and_gate and_gate_h_u_arrmul24_and8_19(a[8], b[19], h_u_arrmul24_and8_19);
  fa fa_h_u_arrmul24_fa8_19_out(h_u_arrmul24_and8_19[0], h_u_arrmul24_fa9_18_xor1[0], h_u_arrmul24_fa7_19_or0[0], h_u_arrmul24_fa8_19_xor1, h_u_arrmul24_fa8_19_or0);
  and_gate and_gate_h_u_arrmul24_and9_19(a[9], b[19], h_u_arrmul24_and9_19);
  fa fa_h_u_arrmul24_fa9_19_out(h_u_arrmul24_and9_19[0], h_u_arrmul24_fa10_18_xor1[0], h_u_arrmul24_fa8_19_or0[0], h_u_arrmul24_fa9_19_xor1, h_u_arrmul24_fa9_19_or0);
  and_gate and_gate_h_u_arrmul24_and10_19(a[10], b[19], h_u_arrmul24_and10_19);
  fa fa_h_u_arrmul24_fa10_19_out(h_u_arrmul24_and10_19[0], h_u_arrmul24_fa11_18_xor1[0], h_u_arrmul24_fa9_19_or0[0], h_u_arrmul24_fa10_19_xor1, h_u_arrmul24_fa10_19_or0);
  and_gate and_gate_h_u_arrmul24_and11_19(a[11], b[19], h_u_arrmul24_and11_19);
  fa fa_h_u_arrmul24_fa11_19_out(h_u_arrmul24_and11_19[0], h_u_arrmul24_fa12_18_xor1[0], h_u_arrmul24_fa10_19_or0[0], h_u_arrmul24_fa11_19_xor1, h_u_arrmul24_fa11_19_or0);
  and_gate and_gate_h_u_arrmul24_and12_19(a[12], b[19], h_u_arrmul24_and12_19);
  fa fa_h_u_arrmul24_fa12_19_out(h_u_arrmul24_and12_19[0], h_u_arrmul24_fa13_18_xor1[0], h_u_arrmul24_fa11_19_or0[0], h_u_arrmul24_fa12_19_xor1, h_u_arrmul24_fa12_19_or0);
  and_gate and_gate_h_u_arrmul24_and13_19(a[13], b[19], h_u_arrmul24_and13_19);
  fa fa_h_u_arrmul24_fa13_19_out(h_u_arrmul24_and13_19[0], h_u_arrmul24_fa14_18_xor1[0], h_u_arrmul24_fa12_19_or0[0], h_u_arrmul24_fa13_19_xor1, h_u_arrmul24_fa13_19_or0);
  and_gate and_gate_h_u_arrmul24_and14_19(a[14], b[19], h_u_arrmul24_and14_19);
  fa fa_h_u_arrmul24_fa14_19_out(h_u_arrmul24_and14_19[0], h_u_arrmul24_fa15_18_xor1[0], h_u_arrmul24_fa13_19_or0[0], h_u_arrmul24_fa14_19_xor1, h_u_arrmul24_fa14_19_or0);
  and_gate and_gate_h_u_arrmul24_and15_19(a[15], b[19], h_u_arrmul24_and15_19);
  fa fa_h_u_arrmul24_fa15_19_out(h_u_arrmul24_and15_19[0], h_u_arrmul24_fa16_18_xor1[0], h_u_arrmul24_fa14_19_or0[0], h_u_arrmul24_fa15_19_xor1, h_u_arrmul24_fa15_19_or0);
  and_gate and_gate_h_u_arrmul24_and16_19(a[16], b[19], h_u_arrmul24_and16_19);
  fa fa_h_u_arrmul24_fa16_19_out(h_u_arrmul24_and16_19[0], h_u_arrmul24_fa17_18_xor1[0], h_u_arrmul24_fa15_19_or0[0], h_u_arrmul24_fa16_19_xor1, h_u_arrmul24_fa16_19_or0);
  and_gate and_gate_h_u_arrmul24_and17_19(a[17], b[19], h_u_arrmul24_and17_19);
  fa fa_h_u_arrmul24_fa17_19_out(h_u_arrmul24_and17_19[0], h_u_arrmul24_fa18_18_xor1[0], h_u_arrmul24_fa16_19_or0[0], h_u_arrmul24_fa17_19_xor1, h_u_arrmul24_fa17_19_or0);
  and_gate and_gate_h_u_arrmul24_and18_19(a[18], b[19], h_u_arrmul24_and18_19);
  fa fa_h_u_arrmul24_fa18_19_out(h_u_arrmul24_and18_19[0], h_u_arrmul24_fa19_18_xor1[0], h_u_arrmul24_fa17_19_or0[0], h_u_arrmul24_fa18_19_xor1, h_u_arrmul24_fa18_19_or0);
  and_gate and_gate_h_u_arrmul24_and19_19(a[19], b[19], h_u_arrmul24_and19_19);
  fa fa_h_u_arrmul24_fa19_19_out(h_u_arrmul24_and19_19[0], h_u_arrmul24_fa20_18_xor1[0], h_u_arrmul24_fa18_19_or0[0], h_u_arrmul24_fa19_19_xor1, h_u_arrmul24_fa19_19_or0);
  and_gate and_gate_h_u_arrmul24_and20_19(a[20], b[19], h_u_arrmul24_and20_19);
  fa fa_h_u_arrmul24_fa20_19_out(h_u_arrmul24_and20_19[0], h_u_arrmul24_fa21_18_xor1[0], h_u_arrmul24_fa19_19_or0[0], h_u_arrmul24_fa20_19_xor1, h_u_arrmul24_fa20_19_or0);
  and_gate and_gate_h_u_arrmul24_and21_19(a[21], b[19], h_u_arrmul24_and21_19);
  fa fa_h_u_arrmul24_fa21_19_out(h_u_arrmul24_and21_19[0], h_u_arrmul24_fa22_18_xor1[0], h_u_arrmul24_fa20_19_or0[0], h_u_arrmul24_fa21_19_xor1, h_u_arrmul24_fa21_19_or0);
  and_gate and_gate_h_u_arrmul24_and22_19(a[22], b[19], h_u_arrmul24_and22_19);
  fa fa_h_u_arrmul24_fa22_19_out(h_u_arrmul24_and22_19[0], h_u_arrmul24_fa23_18_xor1[0], h_u_arrmul24_fa21_19_or0[0], h_u_arrmul24_fa22_19_xor1, h_u_arrmul24_fa22_19_or0);
  and_gate and_gate_h_u_arrmul24_and23_19(a[23], b[19], h_u_arrmul24_and23_19);
  fa fa_h_u_arrmul24_fa23_19_out(h_u_arrmul24_and23_19[0], h_u_arrmul24_fa23_18_or0[0], h_u_arrmul24_fa22_19_or0[0], h_u_arrmul24_fa23_19_xor1, h_u_arrmul24_fa23_19_or0);
  and_gate and_gate_h_u_arrmul24_and0_20(a[0], b[20], h_u_arrmul24_and0_20);
  ha ha_h_u_arrmul24_ha0_20_out(h_u_arrmul24_and0_20[0], h_u_arrmul24_fa1_19_xor1[0], h_u_arrmul24_ha0_20_xor0, h_u_arrmul24_ha0_20_and0);
  and_gate and_gate_h_u_arrmul24_and1_20(a[1], b[20], h_u_arrmul24_and1_20);
  fa fa_h_u_arrmul24_fa1_20_out(h_u_arrmul24_and1_20[0], h_u_arrmul24_fa2_19_xor1[0], h_u_arrmul24_ha0_20_and0[0], h_u_arrmul24_fa1_20_xor1, h_u_arrmul24_fa1_20_or0);
  and_gate and_gate_h_u_arrmul24_and2_20(a[2], b[20], h_u_arrmul24_and2_20);
  fa fa_h_u_arrmul24_fa2_20_out(h_u_arrmul24_and2_20[0], h_u_arrmul24_fa3_19_xor1[0], h_u_arrmul24_fa1_20_or0[0], h_u_arrmul24_fa2_20_xor1, h_u_arrmul24_fa2_20_or0);
  and_gate and_gate_h_u_arrmul24_and3_20(a[3], b[20], h_u_arrmul24_and3_20);
  fa fa_h_u_arrmul24_fa3_20_out(h_u_arrmul24_and3_20[0], h_u_arrmul24_fa4_19_xor1[0], h_u_arrmul24_fa2_20_or0[0], h_u_arrmul24_fa3_20_xor1, h_u_arrmul24_fa3_20_or0);
  and_gate and_gate_h_u_arrmul24_and4_20(a[4], b[20], h_u_arrmul24_and4_20);
  fa fa_h_u_arrmul24_fa4_20_out(h_u_arrmul24_and4_20[0], h_u_arrmul24_fa5_19_xor1[0], h_u_arrmul24_fa3_20_or0[0], h_u_arrmul24_fa4_20_xor1, h_u_arrmul24_fa4_20_or0);
  and_gate and_gate_h_u_arrmul24_and5_20(a[5], b[20], h_u_arrmul24_and5_20);
  fa fa_h_u_arrmul24_fa5_20_out(h_u_arrmul24_and5_20[0], h_u_arrmul24_fa6_19_xor1[0], h_u_arrmul24_fa4_20_or0[0], h_u_arrmul24_fa5_20_xor1, h_u_arrmul24_fa5_20_or0);
  and_gate and_gate_h_u_arrmul24_and6_20(a[6], b[20], h_u_arrmul24_and6_20);
  fa fa_h_u_arrmul24_fa6_20_out(h_u_arrmul24_and6_20[0], h_u_arrmul24_fa7_19_xor1[0], h_u_arrmul24_fa5_20_or0[0], h_u_arrmul24_fa6_20_xor1, h_u_arrmul24_fa6_20_or0);
  and_gate and_gate_h_u_arrmul24_and7_20(a[7], b[20], h_u_arrmul24_and7_20);
  fa fa_h_u_arrmul24_fa7_20_out(h_u_arrmul24_and7_20[0], h_u_arrmul24_fa8_19_xor1[0], h_u_arrmul24_fa6_20_or0[0], h_u_arrmul24_fa7_20_xor1, h_u_arrmul24_fa7_20_or0);
  and_gate and_gate_h_u_arrmul24_and8_20(a[8], b[20], h_u_arrmul24_and8_20);
  fa fa_h_u_arrmul24_fa8_20_out(h_u_arrmul24_and8_20[0], h_u_arrmul24_fa9_19_xor1[0], h_u_arrmul24_fa7_20_or0[0], h_u_arrmul24_fa8_20_xor1, h_u_arrmul24_fa8_20_or0);
  and_gate and_gate_h_u_arrmul24_and9_20(a[9], b[20], h_u_arrmul24_and9_20);
  fa fa_h_u_arrmul24_fa9_20_out(h_u_arrmul24_and9_20[0], h_u_arrmul24_fa10_19_xor1[0], h_u_arrmul24_fa8_20_or0[0], h_u_arrmul24_fa9_20_xor1, h_u_arrmul24_fa9_20_or0);
  and_gate and_gate_h_u_arrmul24_and10_20(a[10], b[20], h_u_arrmul24_and10_20);
  fa fa_h_u_arrmul24_fa10_20_out(h_u_arrmul24_and10_20[0], h_u_arrmul24_fa11_19_xor1[0], h_u_arrmul24_fa9_20_or0[0], h_u_arrmul24_fa10_20_xor1, h_u_arrmul24_fa10_20_or0);
  and_gate and_gate_h_u_arrmul24_and11_20(a[11], b[20], h_u_arrmul24_and11_20);
  fa fa_h_u_arrmul24_fa11_20_out(h_u_arrmul24_and11_20[0], h_u_arrmul24_fa12_19_xor1[0], h_u_arrmul24_fa10_20_or0[0], h_u_arrmul24_fa11_20_xor1, h_u_arrmul24_fa11_20_or0);
  and_gate and_gate_h_u_arrmul24_and12_20(a[12], b[20], h_u_arrmul24_and12_20);
  fa fa_h_u_arrmul24_fa12_20_out(h_u_arrmul24_and12_20[0], h_u_arrmul24_fa13_19_xor1[0], h_u_arrmul24_fa11_20_or0[0], h_u_arrmul24_fa12_20_xor1, h_u_arrmul24_fa12_20_or0);
  and_gate and_gate_h_u_arrmul24_and13_20(a[13], b[20], h_u_arrmul24_and13_20);
  fa fa_h_u_arrmul24_fa13_20_out(h_u_arrmul24_and13_20[0], h_u_arrmul24_fa14_19_xor1[0], h_u_arrmul24_fa12_20_or0[0], h_u_arrmul24_fa13_20_xor1, h_u_arrmul24_fa13_20_or0);
  and_gate and_gate_h_u_arrmul24_and14_20(a[14], b[20], h_u_arrmul24_and14_20);
  fa fa_h_u_arrmul24_fa14_20_out(h_u_arrmul24_and14_20[0], h_u_arrmul24_fa15_19_xor1[0], h_u_arrmul24_fa13_20_or0[0], h_u_arrmul24_fa14_20_xor1, h_u_arrmul24_fa14_20_or0);
  and_gate and_gate_h_u_arrmul24_and15_20(a[15], b[20], h_u_arrmul24_and15_20);
  fa fa_h_u_arrmul24_fa15_20_out(h_u_arrmul24_and15_20[0], h_u_arrmul24_fa16_19_xor1[0], h_u_arrmul24_fa14_20_or0[0], h_u_arrmul24_fa15_20_xor1, h_u_arrmul24_fa15_20_or0);
  and_gate and_gate_h_u_arrmul24_and16_20(a[16], b[20], h_u_arrmul24_and16_20);
  fa fa_h_u_arrmul24_fa16_20_out(h_u_arrmul24_and16_20[0], h_u_arrmul24_fa17_19_xor1[0], h_u_arrmul24_fa15_20_or0[0], h_u_arrmul24_fa16_20_xor1, h_u_arrmul24_fa16_20_or0);
  and_gate and_gate_h_u_arrmul24_and17_20(a[17], b[20], h_u_arrmul24_and17_20);
  fa fa_h_u_arrmul24_fa17_20_out(h_u_arrmul24_and17_20[0], h_u_arrmul24_fa18_19_xor1[0], h_u_arrmul24_fa16_20_or0[0], h_u_arrmul24_fa17_20_xor1, h_u_arrmul24_fa17_20_or0);
  and_gate and_gate_h_u_arrmul24_and18_20(a[18], b[20], h_u_arrmul24_and18_20);
  fa fa_h_u_arrmul24_fa18_20_out(h_u_arrmul24_and18_20[0], h_u_arrmul24_fa19_19_xor1[0], h_u_arrmul24_fa17_20_or0[0], h_u_arrmul24_fa18_20_xor1, h_u_arrmul24_fa18_20_or0);
  and_gate and_gate_h_u_arrmul24_and19_20(a[19], b[20], h_u_arrmul24_and19_20);
  fa fa_h_u_arrmul24_fa19_20_out(h_u_arrmul24_and19_20[0], h_u_arrmul24_fa20_19_xor1[0], h_u_arrmul24_fa18_20_or0[0], h_u_arrmul24_fa19_20_xor1, h_u_arrmul24_fa19_20_or0);
  and_gate and_gate_h_u_arrmul24_and20_20(a[20], b[20], h_u_arrmul24_and20_20);
  fa fa_h_u_arrmul24_fa20_20_out(h_u_arrmul24_and20_20[0], h_u_arrmul24_fa21_19_xor1[0], h_u_arrmul24_fa19_20_or0[0], h_u_arrmul24_fa20_20_xor1, h_u_arrmul24_fa20_20_or0);
  and_gate and_gate_h_u_arrmul24_and21_20(a[21], b[20], h_u_arrmul24_and21_20);
  fa fa_h_u_arrmul24_fa21_20_out(h_u_arrmul24_and21_20[0], h_u_arrmul24_fa22_19_xor1[0], h_u_arrmul24_fa20_20_or0[0], h_u_arrmul24_fa21_20_xor1, h_u_arrmul24_fa21_20_or0);
  and_gate and_gate_h_u_arrmul24_and22_20(a[22], b[20], h_u_arrmul24_and22_20);
  fa fa_h_u_arrmul24_fa22_20_out(h_u_arrmul24_and22_20[0], h_u_arrmul24_fa23_19_xor1[0], h_u_arrmul24_fa21_20_or0[0], h_u_arrmul24_fa22_20_xor1, h_u_arrmul24_fa22_20_or0);
  and_gate and_gate_h_u_arrmul24_and23_20(a[23], b[20], h_u_arrmul24_and23_20);
  fa fa_h_u_arrmul24_fa23_20_out(h_u_arrmul24_and23_20[0], h_u_arrmul24_fa23_19_or0[0], h_u_arrmul24_fa22_20_or0[0], h_u_arrmul24_fa23_20_xor1, h_u_arrmul24_fa23_20_or0);
  and_gate and_gate_h_u_arrmul24_and0_21(a[0], b[21], h_u_arrmul24_and0_21);
  ha ha_h_u_arrmul24_ha0_21_out(h_u_arrmul24_and0_21[0], h_u_arrmul24_fa1_20_xor1[0], h_u_arrmul24_ha0_21_xor0, h_u_arrmul24_ha0_21_and0);
  and_gate and_gate_h_u_arrmul24_and1_21(a[1], b[21], h_u_arrmul24_and1_21);
  fa fa_h_u_arrmul24_fa1_21_out(h_u_arrmul24_and1_21[0], h_u_arrmul24_fa2_20_xor1[0], h_u_arrmul24_ha0_21_and0[0], h_u_arrmul24_fa1_21_xor1, h_u_arrmul24_fa1_21_or0);
  and_gate and_gate_h_u_arrmul24_and2_21(a[2], b[21], h_u_arrmul24_and2_21);
  fa fa_h_u_arrmul24_fa2_21_out(h_u_arrmul24_and2_21[0], h_u_arrmul24_fa3_20_xor1[0], h_u_arrmul24_fa1_21_or0[0], h_u_arrmul24_fa2_21_xor1, h_u_arrmul24_fa2_21_or0);
  and_gate and_gate_h_u_arrmul24_and3_21(a[3], b[21], h_u_arrmul24_and3_21);
  fa fa_h_u_arrmul24_fa3_21_out(h_u_arrmul24_and3_21[0], h_u_arrmul24_fa4_20_xor1[0], h_u_arrmul24_fa2_21_or0[0], h_u_arrmul24_fa3_21_xor1, h_u_arrmul24_fa3_21_or0);
  and_gate and_gate_h_u_arrmul24_and4_21(a[4], b[21], h_u_arrmul24_and4_21);
  fa fa_h_u_arrmul24_fa4_21_out(h_u_arrmul24_and4_21[0], h_u_arrmul24_fa5_20_xor1[0], h_u_arrmul24_fa3_21_or0[0], h_u_arrmul24_fa4_21_xor1, h_u_arrmul24_fa4_21_or0);
  and_gate and_gate_h_u_arrmul24_and5_21(a[5], b[21], h_u_arrmul24_and5_21);
  fa fa_h_u_arrmul24_fa5_21_out(h_u_arrmul24_and5_21[0], h_u_arrmul24_fa6_20_xor1[0], h_u_arrmul24_fa4_21_or0[0], h_u_arrmul24_fa5_21_xor1, h_u_arrmul24_fa5_21_or0);
  and_gate and_gate_h_u_arrmul24_and6_21(a[6], b[21], h_u_arrmul24_and6_21);
  fa fa_h_u_arrmul24_fa6_21_out(h_u_arrmul24_and6_21[0], h_u_arrmul24_fa7_20_xor1[0], h_u_arrmul24_fa5_21_or0[0], h_u_arrmul24_fa6_21_xor1, h_u_arrmul24_fa6_21_or0);
  and_gate and_gate_h_u_arrmul24_and7_21(a[7], b[21], h_u_arrmul24_and7_21);
  fa fa_h_u_arrmul24_fa7_21_out(h_u_arrmul24_and7_21[0], h_u_arrmul24_fa8_20_xor1[0], h_u_arrmul24_fa6_21_or0[0], h_u_arrmul24_fa7_21_xor1, h_u_arrmul24_fa7_21_or0);
  and_gate and_gate_h_u_arrmul24_and8_21(a[8], b[21], h_u_arrmul24_and8_21);
  fa fa_h_u_arrmul24_fa8_21_out(h_u_arrmul24_and8_21[0], h_u_arrmul24_fa9_20_xor1[0], h_u_arrmul24_fa7_21_or0[0], h_u_arrmul24_fa8_21_xor1, h_u_arrmul24_fa8_21_or0);
  and_gate and_gate_h_u_arrmul24_and9_21(a[9], b[21], h_u_arrmul24_and9_21);
  fa fa_h_u_arrmul24_fa9_21_out(h_u_arrmul24_and9_21[0], h_u_arrmul24_fa10_20_xor1[0], h_u_arrmul24_fa8_21_or0[0], h_u_arrmul24_fa9_21_xor1, h_u_arrmul24_fa9_21_or0);
  and_gate and_gate_h_u_arrmul24_and10_21(a[10], b[21], h_u_arrmul24_and10_21);
  fa fa_h_u_arrmul24_fa10_21_out(h_u_arrmul24_and10_21[0], h_u_arrmul24_fa11_20_xor1[0], h_u_arrmul24_fa9_21_or0[0], h_u_arrmul24_fa10_21_xor1, h_u_arrmul24_fa10_21_or0);
  and_gate and_gate_h_u_arrmul24_and11_21(a[11], b[21], h_u_arrmul24_and11_21);
  fa fa_h_u_arrmul24_fa11_21_out(h_u_arrmul24_and11_21[0], h_u_arrmul24_fa12_20_xor1[0], h_u_arrmul24_fa10_21_or0[0], h_u_arrmul24_fa11_21_xor1, h_u_arrmul24_fa11_21_or0);
  and_gate and_gate_h_u_arrmul24_and12_21(a[12], b[21], h_u_arrmul24_and12_21);
  fa fa_h_u_arrmul24_fa12_21_out(h_u_arrmul24_and12_21[0], h_u_arrmul24_fa13_20_xor1[0], h_u_arrmul24_fa11_21_or0[0], h_u_arrmul24_fa12_21_xor1, h_u_arrmul24_fa12_21_or0);
  and_gate and_gate_h_u_arrmul24_and13_21(a[13], b[21], h_u_arrmul24_and13_21);
  fa fa_h_u_arrmul24_fa13_21_out(h_u_arrmul24_and13_21[0], h_u_arrmul24_fa14_20_xor1[0], h_u_arrmul24_fa12_21_or0[0], h_u_arrmul24_fa13_21_xor1, h_u_arrmul24_fa13_21_or0);
  and_gate and_gate_h_u_arrmul24_and14_21(a[14], b[21], h_u_arrmul24_and14_21);
  fa fa_h_u_arrmul24_fa14_21_out(h_u_arrmul24_and14_21[0], h_u_arrmul24_fa15_20_xor1[0], h_u_arrmul24_fa13_21_or0[0], h_u_arrmul24_fa14_21_xor1, h_u_arrmul24_fa14_21_or0);
  and_gate and_gate_h_u_arrmul24_and15_21(a[15], b[21], h_u_arrmul24_and15_21);
  fa fa_h_u_arrmul24_fa15_21_out(h_u_arrmul24_and15_21[0], h_u_arrmul24_fa16_20_xor1[0], h_u_arrmul24_fa14_21_or0[0], h_u_arrmul24_fa15_21_xor1, h_u_arrmul24_fa15_21_or0);
  and_gate and_gate_h_u_arrmul24_and16_21(a[16], b[21], h_u_arrmul24_and16_21);
  fa fa_h_u_arrmul24_fa16_21_out(h_u_arrmul24_and16_21[0], h_u_arrmul24_fa17_20_xor1[0], h_u_arrmul24_fa15_21_or0[0], h_u_arrmul24_fa16_21_xor1, h_u_arrmul24_fa16_21_or0);
  and_gate and_gate_h_u_arrmul24_and17_21(a[17], b[21], h_u_arrmul24_and17_21);
  fa fa_h_u_arrmul24_fa17_21_out(h_u_arrmul24_and17_21[0], h_u_arrmul24_fa18_20_xor1[0], h_u_arrmul24_fa16_21_or0[0], h_u_arrmul24_fa17_21_xor1, h_u_arrmul24_fa17_21_or0);
  and_gate and_gate_h_u_arrmul24_and18_21(a[18], b[21], h_u_arrmul24_and18_21);
  fa fa_h_u_arrmul24_fa18_21_out(h_u_arrmul24_and18_21[0], h_u_arrmul24_fa19_20_xor1[0], h_u_arrmul24_fa17_21_or0[0], h_u_arrmul24_fa18_21_xor1, h_u_arrmul24_fa18_21_or0);
  and_gate and_gate_h_u_arrmul24_and19_21(a[19], b[21], h_u_arrmul24_and19_21);
  fa fa_h_u_arrmul24_fa19_21_out(h_u_arrmul24_and19_21[0], h_u_arrmul24_fa20_20_xor1[0], h_u_arrmul24_fa18_21_or0[0], h_u_arrmul24_fa19_21_xor1, h_u_arrmul24_fa19_21_or0);
  and_gate and_gate_h_u_arrmul24_and20_21(a[20], b[21], h_u_arrmul24_and20_21);
  fa fa_h_u_arrmul24_fa20_21_out(h_u_arrmul24_and20_21[0], h_u_arrmul24_fa21_20_xor1[0], h_u_arrmul24_fa19_21_or0[0], h_u_arrmul24_fa20_21_xor1, h_u_arrmul24_fa20_21_or0);
  and_gate and_gate_h_u_arrmul24_and21_21(a[21], b[21], h_u_arrmul24_and21_21);
  fa fa_h_u_arrmul24_fa21_21_out(h_u_arrmul24_and21_21[0], h_u_arrmul24_fa22_20_xor1[0], h_u_arrmul24_fa20_21_or0[0], h_u_arrmul24_fa21_21_xor1, h_u_arrmul24_fa21_21_or0);
  and_gate and_gate_h_u_arrmul24_and22_21(a[22], b[21], h_u_arrmul24_and22_21);
  fa fa_h_u_arrmul24_fa22_21_out(h_u_arrmul24_and22_21[0], h_u_arrmul24_fa23_20_xor1[0], h_u_arrmul24_fa21_21_or0[0], h_u_arrmul24_fa22_21_xor1, h_u_arrmul24_fa22_21_or0);
  and_gate and_gate_h_u_arrmul24_and23_21(a[23], b[21], h_u_arrmul24_and23_21);
  fa fa_h_u_arrmul24_fa23_21_out(h_u_arrmul24_and23_21[0], h_u_arrmul24_fa23_20_or0[0], h_u_arrmul24_fa22_21_or0[0], h_u_arrmul24_fa23_21_xor1, h_u_arrmul24_fa23_21_or0);
  and_gate and_gate_h_u_arrmul24_and0_22(a[0], b[22], h_u_arrmul24_and0_22);
  ha ha_h_u_arrmul24_ha0_22_out(h_u_arrmul24_and0_22[0], h_u_arrmul24_fa1_21_xor1[0], h_u_arrmul24_ha0_22_xor0, h_u_arrmul24_ha0_22_and0);
  and_gate and_gate_h_u_arrmul24_and1_22(a[1], b[22], h_u_arrmul24_and1_22);
  fa fa_h_u_arrmul24_fa1_22_out(h_u_arrmul24_and1_22[0], h_u_arrmul24_fa2_21_xor1[0], h_u_arrmul24_ha0_22_and0[0], h_u_arrmul24_fa1_22_xor1, h_u_arrmul24_fa1_22_or0);
  and_gate and_gate_h_u_arrmul24_and2_22(a[2], b[22], h_u_arrmul24_and2_22);
  fa fa_h_u_arrmul24_fa2_22_out(h_u_arrmul24_and2_22[0], h_u_arrmul24_fa3_21_xor1[0], h_u_arrmul24_fa1_22_or0[0], h_u_arrmul24_fa2_22_xor1, h_u_arrmul24_fa2_22_or0);
  and_gate and_gate_h_u_arrmul24_and3_22(a[3], b[22], h_u_arrmul24_and3_22);
  fa fa_h_u_arrmul24_fa3_22_out(h_u_arrmul24_and3_22[0], h_u_arrmul24_fa4_21_xor1[0], h_u_arrmul24_fa2_22_or0[0], h_u_arrmul24_fa3_22_xor1, h_u_arrmul24_fa3_22_or0);
  and_gate and_gate_h_u_arrmul24_and4_22(a[4], b[22], h_u_arrmul24_and4_22);
  fa fa_h_u_arrmul24_fa4_22_out(h_u_arrmul24_and4_22[0], h_u_arrmul24_fa5_21_xor1[0], h_u_arrmul24_fa3_22_or0[0], h_u_arrmul24_fa4_22_xor1, h_u_arrmul24_fa4_22_or0);
  and_gate and_gate_h_u_arrmul24_and5_22(a[5], b[22], h_u_arrmul24_and5_22);
  fa fa_h_u_arrmul24_fa5_22_out(h_u_arrmul24_and5_22[0], h_u_arrmul24_fa6_21_xor1[0], h_u_arrmul24_fa4_22_or0[0], h_u_arrmul24_fa5_22_xor1, h_u_arrmul24_fa5_22_or0);
  and_gate and_gate_h_u_arrmul24_and6_22(a[6], b[22], h_u_arrmul24_and6_22);
  fa fa_h_u_arrmul24_fa6_22_out(h_u_arrmul24_and6_22[0], h_u_arrmul24_fa7_21_xor1[0], h_u_arrmul24_fa5_22_or0[0], h_u_arrmul24_fa6_22_xor1, h_u_arrmul24_fa6_22_or0);
  and_gate and_gate_h_u_arrmul24_and7_22(a[7], b[22], h_u_arrmul24_and7_22);
  fa fa_h_u_arrmul24_fa7_22_out(h_u_arrmul24_and7_22[0], h_u_arrmul24_fa8_21_xor1[0], h_u_arrmul24_fa6_22_or0[0], h_u_arrmul24_fa7_22_xor1, h_u_arrmul24_fa7_22_or0);
  and_gate and_gate_h_u_arrmul24_and8_22(a[8], b[22], h_u_arrmul24_and8_22);
  fa fa_h_u_arrmul24_fa8_22_out(h_u_arrmul24_and8_22[0], h_u_arrmul24_fa9_21_xor1[0], h_u_arrmul24_fa7_22_or0[0], h_u_arrmul24_fa8_22_xor1, h_u_arrmul24_fa8_22_or0);
  and_gate and_gate_h_u_arrmul24_and9_22(a[9], b[22], h_u_arrmul24_and9_22);
  fa fa_h_u_arrmul24_fa9_22_out(h_u_arrmul24_and9_22[0], h_u_arrmul24_fa10_21_xor1[0], h_u_arrmul24_fa8_22_or0[0], h_u_arrmul24_fa9_22_xor1, h_u_arrmul24_fa9_22_or0);
  and_gate and_gate_h_u_arrmul24_and10_22(a[10], b[22], h_u_arrmul24_and10_22);
  fa fa_h_u_arrmul24_fa10_22_out(h_u_arrmul24_and10_22[0], h_u_arrmul24_fa11_21_xor1[0], h_u_arrmul24_fa9_22_or0[0], h_u_arrmul24_fa10_22_xor1, h_u_arrmul24_fa10_22_or0);
  and_gate and_gate_h_u_arrmul24_and11_22(a[11], b[22], h_u_arrmul24_and11_22);
  fa fa_h_u_arrmul24_fa11_22_out(h_u_arrmul24_and11_22[0], h_u_arrmul24_fa12_21_xor1[0], h_u_arrmul24_fa10_22_or0[0], h_u_arrmul24_fa11_22_xor1, h_u_arrmul24_fa11_22_or0);
  and_gate and_gate_h_u_arrmul24_and12_22(a[12], b[22], h_u_arrmul24_and12_22);
  fa fa_h_u_arrmul24_fa12_22_out(h_u_arrmul24_and12_22[0], h_u_arrmul24_fa13_21_xor1[0], h_u_arrmul24_fa11_22_or0[0], h_u_arrmul24_fa12_22_xor1, h_u_arrmul24_fa12_22_or0);
  and_gate and_gate_h_u_arrmul24_and13_22(a[13], b[22], h_u_arrmul24_and13_22);
  fa fa_h_u_arrmul24_fa13_22_out(h_u_arrmul24_and13_22[0], h_u_arrmul24_fa14_21_xor1[0], h_u_arrmul24_fa12_22_or0[0], h_u_arrmul24_fa13_22_xor1, h_u_arrmul24_fa13_22_or0);
  and_gate and_gate_h_u_arrmul24_and14_22(a[14], b[22], h_u_arrmul24_and14_22);
  fa fa_h_u_arrmul24_fa14_22_out(h_u_arrmul24_and14_22[0], h_u_arrmul24_fa15_21_xor1[0], h_u_arrmul24_fa13_22_or0[0], h_u_arrmul24_fa14_22_xor1, h_u_arrmul24_fa14_22_or0);
  and_gate and_gate_h_u_arrmul24_and15_22(a[15], b[22], h_u_arrmul24_and15_22);
  fa fa_h_u_arrmul24_fa15_22_out(h_u_arrmul24_and15_22[0], h_u_arrmul24_fa16_21_xor1[0], h_u_arrmul24_fa14_22_or0[0], h_u_arrmul24_fa15_22_xor1, h_u_arrmul24_fa15_22_or0);
  and_gate and_gate_h_u_arrmul24_and16_22(a[16], b[22], h_u_arrmul24_and16_22);
  fa fa_h_u_arrmul24_fa16_22_out(h_u_arrmul24_and16_22[0], h_u_arrmul24_fa17_21_xor1[0], h_u_arrmul24_fa15_22_or0[0], h_u_arrmul24_fa16_22_xor1, h_u_arrmul24_fa16_22_or0);
  and_gate and_gate_h_u_arrmul24_and17_22(a[17], b[22], h_u_arrmul24_and17_22);
  fa fa_h_u_arrmul24_fa17_22_out(h_u_arrmul24_and17_22[0], h_u_arrmul24_fa18_21_xor1[0], h_u_arrmul24_fa16_22_or0[0], h_u_arrmul24_fa17_22_xor1, h_u_arrmul24_fa17_22_or0);
  and_gate and_gate_h_u_arrmul24_and18_22(a[18], b[22], h_u_arrmul24_and18_22);
  fa fa_h_u_arrmul24_fa18_22_out(h_u_arrmul24_and18_22[0], h_u_arrmul24_fa19_21_xor1[0], h_u_arrmul24_fa17_22_or0[0], h_u_arrmul24_fa18_22_xor1, h_u_arrmul24_fa18_22_or0);
  and_gate and_gate_h_u_arrmul24_and19_22(a[19], b[22], h_u_arrmul24_and19_22);
  fa fa_h_u_arrmul24_fa19_22_out(h_u_arrmul24_and19_22[0], h_u_arrmul24_fa20_21_xor1[0], h_u_arrmul24_fa18_22_or0[0], h_u_arrmul24_fa19_22_xor1, h_u_arrmul24_fa19_22_or0);
  and_gate and_gate_h_u_arrmul24_and20_22(a[20], b[22], h_u_arrmul24_and20_22);
  fa fa_h_u_arrmul24_fa20_22_out(h_u_arrmul24_and20_22[0], h_u_arrmul24_fa21_21_xor1[0], h_u_arrmul24_fa19_22_or0[0], h_u_arrmul24_fa20_22_xor1, h_u_arrmul24_fa20_22_or0);
  and_gate and_gate_h_u_arrmul24_and21_22(a[21], b[22], h_u_arrmul24_and21_22);
  fa fa_h_u_arrmul24_fa21_22_out(h_u_arrmul24_and21_22[0], h_u_arrmul24_fa22_21_xor1[0], h_u_arrmul24_fa20_22_or0[0], h_u_arrmul24_fa21_22_xor1, h_u_arrmul24_fa21_22_or0);
  and_gate and_gate_h_u_arrmul24_and22_22(a[22], b[22], h_u_arrmul24_and22_22);
  fa fa_h_u_arrmul24_fa22_22_out(h_u_arrmul24_and22_22[0], h_u_arrmul24_fa23_21_xor1[0], h_u_arrmul24_fa21_22_or0[0], h_u_arrmul24_fa22_22_xor1, h_u_arrmul24_fa22_22_or0);
  and_gate and_gate_h_u_arrmul24_and23_22(a[23], b[22], h_u_arrmul24_and23_22);
  fa fa_h_u_arrmul24_fa23_22_out(h_u_arrmul24_and23_22[0], h_u_arrmul24_fa23_21_or0[0], h_u_arrmul24_fa22_22_or0[0], h_u_arrmul24_fa23_22_xor1, h_u_arrmul24_fa23_22_or0);
  and_gate and_gate_h_u_arrmul24_and0_23(a[0], b[23], h_u_arrmul24_and0_23);
  ha ha_h_u_arrmul24_ha0_23_out(h_u_arrmul24_and0_23[0], h_u_arrmul24_fa1_22_xor1[0], h_u_arrmul24_ha0_23_xor0, h_u_arrmul24_ha0_23_and0);
  and_gate and_gate_h_u_arrmul24_and1_23(a[1], b[23], h_u_arrmul24_and1_23);
  fa fa_h_u_arrmul24_fa1_23_out(h_u_arrmul24_and1_23[0], h_u_arrmul24_fa2_22_xor1[0], h_u_arrmul24_ha0_23_and0[0], h_u_arrmul24_fa1_23_xor1, h_u_arrmul24_fa1_23_or0);
  and_gate and_gate_h_u_arrmul24_and2_23(a[2], b[23], h_u_arrmul24_and2_23);
  fa fa_h_u_arrmul24_fa2_23_out(h_u_arrmul24_and2_23[0], h_u_arrmul24_fa3_22_xor1[0], h_u_arrmul24_fa1_23_or0[0], h_u_arrmul24_fa2_23_xor1, h_u_arrmul24_fa2_23_or0);
  and_gate and_gate_h_u_arrmul24_and3_23(a[3], b[23], h_u_arrmul24_and3_23);
  fa fa_h_u_arrmul24_fa3_23_out(h_u_arrmul24_and3_23[0], h_u_arrmul24_fa4_22_xor1[0], h_u_arrmul24_fa2_23_or0[0], h_u_arrmul24_fa3_23_xor1, h_u_arrmul24_fa3_23_or0);
  and_gate and_gate_h_u_arrmul24_and4_23(a[4], b[23], h_u_arrmul24_and4_23);
  fa fa_h_u_arrmul24_fa4_23_out(h_u_arrmul24_and4_23[0], h_u_arrmul24_fa5_22_xor1[0], h_u_arrmul24_fa3_23_or0[0], h_u_arrmul24_fa4_23_xor1, h_u_arrmul24_fa4_23_or0);
  and_gate and_gate_h_u_arrmul24_and5_23(a[5], b[23], h_u_arrmul24_and5_23);
  fa fa_h_u_arrmul24_fa5_23_out(h_u_arrmul24_and5_23[0], h_u_arrmul24_fa6_22_xor1[0], h_u_arrmul24_fa4_23_or0[0], h_u_arrmul24_fa5_23_xor1, h_u_arrmul24_fa5_23_or0);
  and_gate and_gate_h_u_arrmul24_and6_23(a[6], b[23], h_u_arrmul24_and6_23);
  fa fa_h_u_arrmul24_fa6_23_out(h_u_arrmul24_and6_23[0], h_u_arrmul24_fa7_22_xor1[0], h_u_arrmul24_fa5_23_or0[0], h_u_arrmul24_fa6_23_xor1, h_u_arrmul24_fa6_23_or0);
  and_gate and_gate_h_u_arrmul24_and7_23(a[7], b[23], h_u_arrmul24_and7_23);
  fa fa_h_u_arrmul24_fa7_23_out(h_u_arrmul24_and7_23[0], h_u_arrmul24_fa8_22_xor1[0], h_u_arrmul24_fa6_23_or0[0], h_u_arrmul24_fa7_23_xor1, h_u_arrmul24_fa7_23_or0);
  and_gate and_gate_h_u_arrmul24_and8_23(a[8], b[23], h_u_arrmul24_and8_23);
  fa fa_h_u_arrmul24_fa8_23_out(h_u_arrmul24_and8_23[0], h_u_arrmul24_fa9_22_xor1[0], h_u_arrmul24_fa7_23_or0[0], h_u_arrmul24_fa8_23_xor1, h_u_arrmul24_fa8_23_or0);
  and_gate and_gate_h_u_arrmul24_and9_23(a[9], b[23], h_u_arrmul24_and9_23);
  fa fa_h_u_arrmul24_fa9_23_out(h_u_arrmul24_and9_23[0], h_u_arrmul24_fa10_22_xor1[0], h_u_arrmul24_fa8_23_or0[0], h_u_arrmul24_fa9_23_xor1, h_u_arrmul24_fa9_23_or0);
  and_gate and_gate_h_u_arrmul24_and10_23(a[10], b[23], h_u_arrmul24_and10_23);
  fa fa_h_u_arrmul24_fa10_23_out(h_u_arrmul24_and10_23[0], h_u_arrmul24_fa11_22_xor1[0], h_u_arrmul24_fa9_23_or0[0], h_u_arrmul24_fa10_23_xor1, h_u_arrmul24_fa10_23_or0);
  and_gate and_gate_h_u_arrmul24_and11_23(a[11], b[23], h_u_arrmul24_and11_23);
  fa fa_h_u_arrmul24_fa11_23_out(h_u_arrmul24_and11_23[0], h_u_arrmul24_fa12_22_xor1[0], h_u_arrmul24_fa10_23_or0[0], h_u_arrmul24_fa11_23_xor1, h_u_arrmul24_fa11_23_or0);
  and_gate and_gate_h_u_arrmul24_and12_23(a[12], b[23], h_u_arrmul24_and12_23);
  fa fa_h_u_arrmul24_fa12_23_out(h_u_arrmul24_and12_23[0], h_u_arrmul24_fa13_22_xor1[0], h_u_arrmul24_fa11_23_or0[0], h_u_arrmul24_fa12_23_xor1, h_u_arrmul24_fa12_23_or0);
  and_gate and_gate_h_u_arrmul24_and13_23(a[13], b[23], h_u_arrmul24_and13_23);
  fa fa_h_u_arrmul24_fa13_23_out(h_u_arrmul24_and13_23[0], h_u_arrmul24_fa14_22_xor1[0], h_u_arrmul24_fa12_23_or0[0], h_u_arrmul24_fa13_23_xor1, h_u_arrmul24_fa13_23_or0);
  and_gate and_gate_h_u_arrmul24_and14_23(a[14], b[23], h_u_arrmul24_and14_23);
  fa fa_h_u_arrmul24_fa14_23_out(h_u_arrmul24_and14_23[0], h_u_arrmul24_fa15_22_xor1[0], h_u_arrmul24_fa13_23_or0[0], h_u_arrmul24_fa14_23_xor1, h_u_arrmul24_fa14_23_or0);
  and_gate and_gate_h_u_arrmul24_and15_23(a[15], b[23], h_u_arrmul24_and15_23);
  fa fa_h_u_arrmul24_fa15_23_out(h_u_arrmul24_and15_23[0], h_u_arrmul24_fa16_22_xor1[0], h_u_arrmul24_fa14_23_or0[0], h_u_arrmul24_fa15_23_xor1, h_u_arrmul24_fa15_23_or0);
  and_gate and_gate_h_u_arrmul24_and16_23(a[16], b[23], h_u_arrmul24_and16_23);
  fa fa_h_u_arrmul24_fa16_23_out(h_u_arrmul24_and16_23[0], h_u_arrmul24_fa17_22_xor1[0], h_u_arrmul24_fa15_23_or0[0], h_u_arrmul24_fa16_23_xor1, h_u_arrmul24_fa16_23_or0);
  and_gate and_gate_h_u_arrmul24_and17_23(a[17], b[23], h_u_arrmul24_and17_23);
  fa fa_h_u_arrmul24_fa17_23_out(h_u_arrmul24_and17_23[0], h_u_arrmul24_fa18_22_xor1[0], h_u_arrmul24_fa16_23_or0[0], h_u_arrmul24_fa17_23_xor1, h_u_arrmul24_fa17_23_or0);
  and_gate and_gate_h_u_arrmul24_and18_23(a[18], b[23], h_u_arrmul24_and18_23);
  fa fa_h_u_arrmul24_fa18_23_out(h_u_arrmul24_and18_23[0], h_u_arrmul24_fa19_22_xor1[0], h_u_arrmul24_fa17_23_or0[0], h_u_arrmul24_fa18_23_xor1, h_u_arrmul24_fa18_23_or0);
  and_gate and_gate_h_u_arrmul24_and19_23(a[19], b[23], h_u_arrmul24_and19_23);
  fa fa_h_u_arrmul24_fa19_23_out(h_u_arrmul24_and19_23[0], h_u_arrmul24_fa20_22_xor1[0], h_u_arrmul24_fa18_23_or0[0], h_u_arrmul24_fa19_23_xor1, h_u_arrmul24_fa19_23_or0);
  and_gate and_gate_h_u_arrmul24_and20_23(a[20], b[23], h_u_arrmul24_and20_23);
  fa fa_h_u_arrmul24_fa20_23_out(h_u_arrmul24_and20_23[0], h_u_arrmul24_fa21_22_xor1[0], h_u_arrmul24_fa19_23_or0[0], h_u_arrmul24_fa20_23_xor1, h_u_arrmul24_fa20_23_or0);
  and_gate and_gate_h_u_arrmul24_and21_23(a[21], b[23], h_u_arrmul24_and21_23);
  fa fa_h_u_arrmul24_fa21_23_out(h_u_arrmul24_and21_23[0], h_u_arrmul24_fa22_22_xor1[0], h_u_arrmul24_fa20_23_or0[0], h_u_arrmul24_fa21_23_xor1, h_u_arrmul24_fa21_23_or0);
  and_gate and_gate_h_u_arrmul24_and22_23(a[22], b[23], h_u_arrmul24_and22_23);
  fa fa_h_u_arrmul24_fa22_23_out(h_u_arrmul24_and22_23[0], h_u_arrmul24_fa23_22_xor1[0], h_u_arrmul24_fa21_23_or0[0], h_u_arrmul24_fa22_23_xor1, h_u_arrmul24_fa22_23_or0);
  and_gate and_gate_h_u_arrmul24_and23_23(a[23], b[23], h_u_arrmul24_and23_23);
  fa fa_h_u_arrmul24_fa23_23_out(h_u_arrmul24_and23_23[0], h_u_arrmul24_fa23_22_or0[0], h_u_arrmul24_fa22_23_or0[0], h_u_arrmul24_fa23_23_xor1, h_u_arrmul24_fa23_23_or0);

  assign h_u_arrmul24_out[0] = h_u_arrmul24_and0_0[0];
  assign h_u_arrmul24_out[1] = h_u_arrmul24_ha0_1_xor0[0];
  assign h_u_arrmul24_out[2] = h_u_arrmul24_ha0_2_xor0[0];
  assign h_u_arrmul24_out[3] = h_u_arrmul24_ha0_3_xor0[0];
  assign h_u_arrmul24_out[4] = h_u_arrmul24_ha0_4_xor0[0];
  assign h_u_arrmul24_out[5] = h_u_arrmul24_ha0_5_xor0[0];
  assign h_u_arrmul24_out[6] = h_u_arrmul24_ha0_6_xor0[0];
  assign h_u_arrmul24_out[7] = h_u_arrmul24_ha0_7_xor0[0];
  assign h_u_arrmul24_out[8] = h_u_arrmul24_ha0_8_xor0[0];
  assign h_u_arrmul24_out[9] = h_u_arrmul24_ha0_9_xor0[0];
  assign h_u_arrmul24_out[10] = h_u_arrmul24_ha0_10_xor0[0];
  assign h_u_arrmul24_out[11] = h_u_arrmul24_ha0_11_xor0[0];
  assign h_u_arrmul24_out[12] = h_u_arrmul24_ha0_12_xor0[0];
  assign h_u_arrmul24_out[13] = h_u_arrmul24_ha0_13_xor0[0];
  assign h_u_arrmul24_out[14] = h_u_arrmul24_ha0_14_xor0[0];
  assign h_u_arrmul24_out[15] = h_u_arrmul24_ha0_15_xor0[0];
  assign h_u_arrmul24_out[16] = h_u_arrmul24_ha0_16_xor0[0];
  assign h_u_arrmul24_out[17] = h_u_arrmul24_ha0_17_xor0[0];
  assign h_u_arrmul24_out[18] = h_u_arrmul24_ha0_18_xor0[0];
  assign h_u_arrmul24_out[19] = h_u_arrmul24_ha0_19_xor0[0];
  assign h_u_arrmul24_out[20] = h_u_arrmul24_ha0_20_xor0[0];
  assign h_u_arrmul24_out[21] = h_u_arrmul24_ha0_21_xor0[0];
  assign h_u_arrmul24_out[22] = h_u_arrmul24_ha0_22_xor0[0];
  assign h_u_arrmul24_out[23] = h_u_arrmul24_ha0_23_xor0[0];
  assign h_u_arrmul24_out[24] = h_u_arrmul24_fa1_23_xor1[0];
  assign h_u_arrmul24_out[25] = h_u_arrmul24_fa2_23_xor1[0];
  assign h_u_arrmul24_out[26] = h_u_arrmul24_fa3_23_xor1[0];
  assign h_u_arrmul24_out[27] = h_u_arrmul24_fa4_23_xor1[0];
  assign h_u_arrmul24_out[28] = h_u_arrmul24_fa5_23_xor1[0];
  assign h_u_arrmul24_out[29] = h_u_arrmul24_fa6_23_xor1[0];
  assign h_u_arrmul24_out[30] = h_u_arrmul24_fa7_23_xor1[0];
  assign h_u_arrmul24_out[31] = h_u_arrmul24_fa8_23_xor1[0];
  assign h_u_arrmul24_out[32] = h_u_arrmul24_fa9_23_xor1[0];
  assign h_u_arrmul24_out[33] = h_u_arrmul24_fa10_23_xor1[0];
  assign h_u_arrmul24_out[34] = h_u_arrmul24_fa11_23_xor1[0];
  assign h_u_arrmul24_out[35] = h_u_arrmul24_fa12_23_xor1[0];
  assign h_u_arrmul24_out[36] = h_u_arrmul24_fa13_23_xor1[0];
  assign h_u_arrmul24_out[37] = h_u_arrmul24_fa14_23_xor1[0];
  assign h_u_arrmul24_out[38] = h_u_arrmul24_fa15_23_xor1[0];
  assign h_u_arrmul24_out[39] = h_u_arrmul24_fa16_23_xor1[0];
  assign h_u_arrmul24_out[40] = h_u_arrmul24_fa17_23_xor1[0];
  assign h_u_arrmul24_out[41] = h_u_arrmul24_fa18_23_xor1[0];
  assign h_u_arrmul24_out[42] = h_u_arrmul24_fa19_23_xor1[0];
  assign h_u_arrmul24_out[43] = h_u_arrmul24_fa20_23_xor1[0];
  assign h_u_arrmul24_out[44] = h_u_arrmul24_fa21_23_xor1[0];
  assign h_u_arrmul24_out[45] = h_u_arrmul24_fa22_23_xor1[0];
  assign h_u_arrmul24_out[46] = h_u_arrmul24_fa23_23_xor1[0];
  assign h_u_arrmul24_out[47] = h_u_arrmul24_fa23_23_or0[0];
endmodule