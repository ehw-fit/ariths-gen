module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(.a(a[0]), .b(b[0]), .out(pg_logic_or0));
  and_gate and_gate_pg_logic_and0(.a(a[0]), .b(b[0]), .out(pg_logic_and0));
  xor_gate xor_gate_pg_logic_xor0(.a(a[0]), .b(b[0]), .out(pg_logic_xor0));
endmodule

module u_cla12(input [11:0] a, input [11:0] b, output [12:0] u_cla12_out);
  wire [0:0] u_cla12_pg_logic0_or0;
  wire [0:0] u_cla12_pg_logic0_and0;
  wire [0:0] u_cla12_pg_logic0_xor0;
  wire [0:0] u_cla12_pg_logic1_or0;
  wire [0:0] u_cla12_pg_logic1_and0;
  wire [0:0] u_cla12_pg_logic1_xor0;
  wire [0:0] u_cla12_xor1;
  wire [0:0] u_cla12_and0;
  wire [0:0] u_cla12_or0;
  wire [0:0] u_cla12_pg_logic2_or0;
  wire [0:0] u_cla12_pg_logic2_and0;
  wire [0:0] u_cla12_pg_logic2_xor0;
  wire [0:0] u_cla12_xor2;
  wire [0:0] u_cla12_and1;
  wire [0:0] u_cla12_and2;
  wire [0:0] u_cla12_and3;
  wire [0:0] u_cla12_and4;
  wire [0:0] u_cla12_or1;
  wire [0:0] u_cla12_or2;
  wire [0:0] u_cla12_pg_logic3_or0;
  wire [0:0] u_cla12_pg_logic3_and0;
  wire [0:0] u_cla12_pg_logic3_xor0;
  wire [0:0] u_cla12_xor3;
  wire [0:0] u_cla12_and5;
  wire [0:0] u_cla12_and6;
  wire [0:0] u_cla12_and7;
  wire [0:0] u_cla12_and8;
  wire [0:0] u_cla12_and9;
  wire [0:0] u_cla12_and10;
  wire [0:0] u_cla12_and11;
  wire [0:0] u_cla12_or3;
  wire [0:0] u_cla12_or4;
  wire [0:0] u_cla12_or5;
  wire [0:0] u_cla12_pg_logic4_or0;
  wire [0:0] u_cla12_pg_logic4_and0;
  wire [0:0] u_cla12_pg_logic4_xor0;
  wire [0:0] u_cla12_xor4;
  wire [0:0] u_cla12_and12;
  wire [0:0] u_cla12_or6;
  wire [0:0] u_cla12_pg_logic5_or0;
  wire [0:0] u_cla12_pg_logic5_and0;
  wire [0:0] u_cla12_pg_logic5_xor0;
  wire [0:0] u_cla12_xor5;
  wire [0:0] u_cla12_and13;
  wire [0:0] u_cla12_and14;
  wire [0:0] u_cla12_and15;
  wire [0:0] u_cla12_or7;
  wire [0:0] u_cla12_or8;
  wire [0:0] u_cla12_pg_logic6_or0;
  wire [0:0] u_cla12_pg_logic6_and0;
  wire [0:0] u_cla12_pg_logic6_xor0;
  wire [0:0] u_cla12_xor6;
  wire [0:0] u_cla12_and16;
  wire [0:0] u_cla12_and17;
  wire [0:0] u_cla12_and18;
  wire [0:0] u_cla12_and19;
  wire [0:0] u_cla12_and20;
  wire [0:0] u_cla12_and21;
  wire [0:0] u_cla12_or9;
  wire [0:0] u_cla12_or10;
  wire [0:0] u_cla12_or11;
  wire [0:0] u_cla12_pg_logic7_or0;
  wire [0:0] u_cla12_pg_logic7_and0;
  wire [0:0] u_cla12_pg_logic7_xor0;
  wire [0:0] u_cla12_xor7;
  wire [0:0] u_cla12_and22;
  wire [0:0] u_cla12_and23;
  wire [0:0] u_cla12_and24;
  wire [0:0] u_cla12_and25;
  wire [0:0] u_cla12_and26;
  wire [0:0] u_cla12_and27;
  wire [0:0] u_cla12_and28;
  wire [0:0] u_cla12_and29;
  wire [0:0] u_cla12_and30;
  wire [0:0] u_cla12_and31;
  wire [0:0] u_cla12_or12;
  wire [0:0] u_cla12_or13;
  wire [0:0] u_cla12_or14;
  wire [0:0] u_cla12_or15;
  wire [0:0] u_cla12_pg_logic8_or0;
  wire [0:0] u_cla12_pg_logic8_and0;
  wire [0:0] u_cla12_pg_logic8_xor0;
  wire [0:0] u_cla12_xor8;
  wire [0:0] u_cla12_and32;
  wire [0:0] u_cla12_or16;
  wire [0:0] u_cla12_pg_logic9_or0;
  wire [0:0] u_cla12_pg_logic9_and0;
  wire [0:0] u_cla12_pg_logic9_xor0;
  wire [0:0] u_cla12_xor9;
  wire [0:0] u_cla12_and33;
  wire [0:0] u_cla12_and34;
  wire [0:0] u_cla12_and35;
  wire [0:0] u_cla12_or17;
  wire [0:0] u_cla12_or18;
  wire [0:0] u_cla12_pg_logic10_or0;
  wire [0:0] u_cla12_pg_logic10_and0;
  wire [0:0] u_cla12_pg_logic10_xor0;
  wire [0:0] u_cla12_xor10;
  wire [0:0] u_cla12_and36;
  wire [0:0] u_cla12_and37;
  wire [0:0] u_cla12_and38;
  wire [0:0] u_cla12_and39;
  wire [0:0] u_cla12_and40;
  wire [0:0] u_cla12_and41;
  wire [0:0] u_cla12_or19;
  wire [0:0] u_cla12_or20;
  wire [0:0] u_cla12_or21;
  wire [0:0] u_cla12_pg_logic11_or0;
  wire [0:0] u_cla12_pg_logic11_and0;
  wire [0:0] u_cla12_pg_logic11_xor0;
  wire [0:0] u_cla12_xor11;
  wire [0:0] u_cla12_and42;
  wire [0:0] u_cla12_and43;
  wire [0:0] u_cla12_and44;
  wire [0:0] u_cla12_and45;
  wire [0:0] u_cla12_and46;
  wire [0:0] u_cla12_and47;
  wire [0:0] u_cla12_and48;
  wire [0:0] u_cla12_and49;
  wire [0:0] u_cla12_and50;
  wire [0:0] u_cla12_and51;
  wire [0:0] u_cla12_or22;
  wire [0:0] u_cla12_or23;
  wire [0:0] u_cla12_or24;
  wire [0:0] u_cla12_or25;

  pg_logic pg_logic_u_cla12_pg_logic0_out(.a(a[0]), .b(b[0]), .pg_logic_or0(u_cla12_pg_logic0_or0), .pg_logic_and0(u_cla12_pg_logic0_and0), .pg_logic_xor0(u_cla12_pg_logic0_xor0));
  pg_logic pg_logic_u_cla12_pg_logic1_out(.a(a[1]), .b(b[1]), .pg_logic_or0(u_cla12_pg_logic1_or0), .pg_logic_and0(u_cla12_pg_logic1_and0), .pg_logic_xor0(u_cla12_pg_logic1_xor0));
  xor_gate xor_gate_u_cla12_xor1(.a(u_cla12_pg_logic1_xor0[0]), .b(u_cla12_pg_logic0_and0[0]), .out(u_cla12_xor1));
  and_gate and_gate_u_cla12_and0(.a(u_cla12_pg_logic0_and0[0]), .b(u_cla12_pg_logic1_or0[0]), .out(u_cla12_and0));
  or_gate or_gate_u_cla12_or0(.a(u_cla12_pg_logic1_and0[0]), .b(u_cla12_and0[0]), .out(u_cla12_or0));
  pg_logic pg_logic_u_cla12_pg_logic2_out(.a(a[2]), .b(b[2]), .pg_logic_or0(u_cla12_pg_logic2_or0), .pg_logic_and0(u_cla12_pg_logic2_and0), .pg_logic_xor0(u_cla12_pg_logic2_xor0));
  xor_gate xor_gate_u_cla12_xor2(.a(u_cla12_pg_logic2_xor0[0]), .b(u_cla12_or0[0]), .out(u_cla12_xor2));
  and_gate and_gate_u_cla12_and1(.a(u_cla12_pg_logic2_or0[0]), .b(u_cla12_pg_logic0_or0[0]), .out(u_cla12_and1));
  and_gate and_gate_u_cla12_and2(.a(u_cla12_pg_logic0_and0[0]), .b(u_cla12_pg_logic2_or0[0]), .out(u_cla12_and2));
  and_gate and_gate_u_cla12_and3(.a(u_cla12_and2[0]), .b(u_cla12_pg_logic1_or0[0]), .out(u_cla12_and3));
  and_gate and_gate_u_cla12_and4(.a(u_cla12_pg_logic1_and0[0]), .b(u_cla12_pg_logic2_or0[0]), .out(u_cla12_and4));
  or_gate or_gate_u_cla12_or1(.a(u_cla12_and3[0]), .b(u_cla12_and4[0]), .out(u_cla12_or1));
  or_gate or_gate_u_cla12_or2(.a(u_cla12_pg_logic2_and0[0]), .b(u_cla12_or1[0]), .out(u_cla12_or2));
  pg_logic pg_logic_u_cla12_pg_logic3_out(.a(a[3]), .b(b[3]), .pg_logic_or0(u_cla12_pg_logic3_or0), .pg_logic_and0(u_cla12_pg_logic3_and0), .pg_logic_xor0(u_cla12_pg_logic3_xor0));
  xor_gate xor_gate_u_cla12_xor3(.a(u_cla12_pg_logic3_xor0[0]), .b(u_cla12_or2[0]), .out(u_cla12_xor3));
  and_gate and_gate_u_cla12_and5(.a(u_cla12_pg_logic3_or0[0]), .b(u_cla12_pg_logic1_or0[0]), .out(u_cla12_and5));
  and_gate and_gate_u_cla12_and6(.a(u_cla12_pg_logic0_and0[0]), .b(u_cla12_pg_logic2_or0[0]), .out(u_cla12_and6));
  and_gate and_gate_u_cla12_and7(.a(u_cla12_pg_logic3_or0[0]), .b(u_cla12_pg_logic1_or0[0]), .out(u_cla12_and7));
  and_gate and_gate_u_cla12_and8(.a(u_cla12_and6[0]), .b(u_cla12_and7[0]), .out(u_cla12_and8));
  and_gate and_gate_u_cla12_and9(.a(u_cla12_pg_logic1_and0[0]), .b(u_cla12_pg_logic3_or0[0]), .out(u_cla12_and9));
  and_gate and_gate_u_cla12_and10(.a(u_cla12_and9[0]), .b(u_cla12_pg_logic2_or0[0]), .out(u_cla12_and10));
  and_gate and_gate_u_cla12_and11(.a(u_cla12_pg_logic2_and0[0]), .b(u_cla12_pg_logic3_or0[0]), .out(u_cla12_and11));
  or_gate or_gate_u_cla12_or3(.a(u_cla12_and8[0]), .b(u_cla12_and11[0]), .out(u_cla12_or3));
  or_gate or_gate_u_cla12_or4(.a(u_cla12_and10[0]), .b(u_cla12_or3[0]), .out(u_cla12_or4));
  or_gate or_gate_u_cla12_or5(.a(u_cla12_pg_logic3_and0[0]), .b(u_cla12_or4[0]), .out(u_cla12_or5));
  pg_logic pg_logic_u_cla12_pg_logic4_out(.a(a[4]), .b(b[4]), .pg_logic_or0(u_cla12_pg_logic4_or0), .pg_logic_and0(u_cla12_pg_logic4_and0), .pg_logic_xor0(u_cla12_pg_logic4_xor0));
  xor_gate xor_gate_u_cla12_xor4(.a(u_cla12_pg_logic4_xor0[0]), .b(u_cla12_or5[0]), .out(u_cla12_xor4));
  and_gate and_gate_u_cla12_and12(.a(u_cla12_or5[0]), .b(u_cla12_pg_logic4_or0[0]), .out(u_cla12_and12));
  or_gate or_gate_u_cla12_or6(.a(u_cla12_pg_logic4_and0[0]), .b(u_cla12_and12[0]), .out(u_cla12_or6));
  pg_logic pg_logic_u_cla12_pg_logic5_out(.a(a[5]), .b(b[5]), .pg_logic_or0(u_cla12_pg_logic5_or0), .pg_logic_and0(u_cla12_pg_logic5_and0), .pg_logic_xor0(u_cla12_pg_logic5_xor0));
  xor_gate xor_gate_u_cla12_xor5(.a(u_cla12_pg_logic5_xor0[0]), .b(u_cla12_or6[0]), .out(u_cla12_xor5));
  and_gate and_gate_u_cla12_and13(.a(u_cla12_or5[0]), .b(u_cla12_pg_logic5_or0[0]), .out(u_cla12_and13));
  and_gate and_gate_u_cla12_and14(.a(u_cla12_and13[0]), .b(u_cla12_pg_logic4_or0[0]), .out(u_cla12_and14));
  and_gate and_gate_u_cla12_and15(.a(u_cla12_pg_logic4_and0[0]), .b(u_cla12_pg_logic5_or0[0]), .out(u_cla12_and15));
  or_gate or_gate_u_cla12_or7(.a(u_cla12_and14[0]), .b(u_cla12_and15[0]), .out(u_cla12_or7));
  or_gate or_gate_u_cla12_or8(.a(u_cla12_pg_logic5_and0[0]), .b(u_cla12_or7[0]), .out(u_cla12_or8));
  pg_logic pg_logic_u_cla12_pg_logic6_out(.a(a[6]), .b(b[6]), .pg_logic_or0(u_cla12_pg_logic6_or0), .pg_logic_and0(u_cla12_pg_logic6_and0), .pg_logic_xor0(u_cla12_pg_logic6_xor0));
  xor_gate xor_gate_u_cla12_xor6(.a(u_cla12_pg_logic6_xor0[0]), .b(u_cla12_or8[0]), .out(u_cla12_xor6));
  and_gate and_gate_u_cla12_and16(.a(u_cla12_or5[0]), .b(u_cla12_pg_logic5_or0[0]), .out(u_cla12_and16));
  and_gate and_gate_u_cla12_and17(.a(u_cla12_pg_logic6_or0[0]), .b(u_cla12_pg_logic4_or0[0]), .out(u_cla12_and17));
  and_gate and_gate_u_cla12_and18(.a(u_cla12_and16[0]), .b(u_cla12_and17[0]), .out(u_cla12_and18));
  and_gate and_gate_u_cla12_and19(.a(u_cla12_pg_logic4_and0[0]), .b(u_cla12_pg_logic6_or0[0]), .out(u_cla12_and19));
  and_gate and_gate_u_cla12_and20(.a(u_cla12_and19[0]), .b(u_cla12_pg_logic5_or0[0]), .out(u_cla12_and20));
  and_gate and_gate_u_cla12_and21(.a(u_cla12_pg_logic5_and0[0]), .b(u_cla12_pg_logic6_or0[0]), .out(u_cla12_and21));
  or_gate or_gate_u_cla12_or9(.a(u_cla12_and18[0]), .b(u_cla12_and20[0]), .out(u_cla12_or9));
  or_gate or_gate_u_cla12_or10(.a(u_cla12_or9[0]), .b(u_cla12_and21[0]), .out(u_cla12_or10));
  or_gate or_gate_u_cla12_or11(.a(u_cla12_pg_logic6_and0[0]), .b(u_cla12_or10[0]), .out(u_cla12_or11));
  pg_logic pg_logic_u_cla12_pg_logic7_out(.a(a[7]), .b(b[7]), .pg_logic_or0(u_cla12_pg_logic7_or0), .pg_logic_and0(u_cla12_pg_logic7_and0), .pg_logic_xor0(u_cla12_pg_logic7_xor0));
  xor_gate xor_gate_u_cla12_xor7(.a(u_cla12_pg_logic7_xor0[0]), .b(u_cla12_or11[0]), .out(u_cla12_xor7));
  and_gate and_gate_u_cla12_and22(.a(u_cla12_or5[0]), .b(u_cla12_pg_logic6_or0[0]), .out(u_cla12_and22));
  and_gate and_gate_u_cla12_and23(.a(u_cla12_pg_logic7_or0[0]), .b(u_cla12_pg_logic5_or0[0]), .out(u_cla12_and23));
  and_gate and_gate_u_cla12_and24(.a(u_cla12_and22[0]), .b(u_cla12_and23[0]), .out(u_cla12_and24));
  and_gate and_gate_u_cla12_and25(.a(u_cla12_and24[0]), .b(u_cla12_pg_logic4_or0[0]), .out(u_cla12_and25));
  and_gate and_gate_u_cla12_and26(.a(u_cla12_pg_logic4_and0[0]), .b(u_cla12_pg_logic6_or0[0]), .out(u_cla12_and26));
  and_gate and_gate_u_cla12_and27(.a(u_cla12_pg_logic7_or0[0]), .b(u_cla12_pg_logic5_or0[0]), .out(u_cla12_and27));
  and_gate and_gate_u_cla12_and28(.a(u_cla12_and26[0]), .b(u_cla12_and27[0]), .out(u_cla12_and28));
  and_gate and_gate_u_cla12_and29(.a(u_cla12_pg_logic5_and0[0]), .b(u_cla12_pg_logic7_or0[0]), .out(u_cla12_and29));
  and_gate and_gate_u_cla12_and30(.a(u_cla12_and29[0]), .b(u_cla12_pg_logic6_or0[0]), .out(u_cla12_and30));
  and_gate and_gate_u_cla12_and31(.a(u_cla12_pg_logic6_and0[0]), .b(u_cla12_pg_logic7_or0[0]), .out(u_cla12_and31));
  or_gate or_gate_u_cla12_or12(.a(u_cla12_and25[0]), .b(u_cla12_and30[0]), .out(u_cla12_or12));
  or_gate or_gate_u_cla12_or13(.a(u_cla12_and28[0]), .b(u_cla12_and31[0]), .out(u_cla12_or13));
  or_gate or_gate_u_cla12_or14(.a(u_cla12_or12[0]), .b(u_cla12_or13[0]), .out(u_cla12_or14));
  or_gate or_gate_u_cla12_or15(.a(u_cla12_pg_logic7_and0[0]), .b(u_cla12_or14[0]), .out(u_cla12_or15));
  pg_logic pg_logic_u_cla12_pg_logic8_out(.a(a[8]), .b(b[8]), .pg_logic_or0(u_cla12_pg_logic8_or0), .pg_logic_and0(u_cla12_pg_logic8_and0), .pg_logic_xor0(u_cla12_pg_logic8_xor0));
  xor_gate xor_gate_u_cla12_xor8(.a(u_cla12_pg_logic8_xor0[0]), .b(u_cla12_or15[0]), .out(u_cla12_xor8));
  and_gate and_gate_u_cla12_and32(.a(u_cla12_or15[0]), .b(u_cla12_pg_logic8_or0[0]), .out(u_cla12_and32));
  or_gate or_gate_u_cla12_or16(.a(u_cla12_pg_logic8_and0[0]), .b(u_cla12_and32[0]), .out(u_cla12_or16));
  pg_logic pg_logic_u_cla12_pg_logic9_out(.a(a[9]), .b(b[9]), .pg_logic_or0(u_cla12_pg_logic9_or0), .pg_logic_and0(u_cla12_pg_logic9_and0), .pg_logic_xor0(u_cla12_pg_logic9_xor0));
  xor_gate xor_gate_u_cla12_xor9(.a(u_cla12_pg_logic9_xor0[0]), .b(u_cla12_or16[0]), .out(u_cla12_xor9));
  and_gate and_gate_u_cla12_and33(.a(u_cla12_or15[0]), .b(u_cla12_pg_logic9_or0[0]), .out(u_cla12_and33));
  and_gate and_gate_u_cla12_and34(.a(u_cla12_and33[0]), .b(u_cla12_pg_logic8_or0[0]), .out(u_cla12_and34));
  and_gate and_gate_u_cla12_and35(.a(u_cla12_pg_logic8_and0[0]), .b(u_cla12_pg_logic9_or0[0]), .out(u_cla12_and35));
  or_gate or_gate_u_cla12_or17(.a(u_cla12_and34[0]), .b(u_cla12_and35[0]), .out(u_cla12_or17));
  or_gate or_gate_u_cla12_or18(.a(u_cla12_pg_logic9_and0[0]), .b(u_cla12_or17[0]), .out(u_cla12_or18));
  pg_logic pg_logic_u_cla12_pg_logic10_out(.a(a[10]), .b(b[10]), .pg_logic_or0(u_cla12_pg_logic10_or0), .pg_logic_and0(u_cla12_pg_logic10_and0), .pg_logic_xor0(u_cla12_pg_logic10_xor0));
  xor_gate xor_gate_u_cla12_xor10(.a(u_cla12_pg_logic10_xor0[0]), .b(u_cla12_or18[0]), .out(u_cla12_xor10));
  and_gate and_gate_u_cla12_and36(.a(u_cla12_or15[0]), .b(u_cla12_pg_logic9_or0[0]), .out(u_cla12_and36));
  and_gate and_gate_u_cla12_and37(.a(u_cla12_pg_logic10_or0[0]), .b(u_cla12_pg_logic8_or0[0]), .out(u_cla12_and37));
  and_gate and_gate_u_cla12_and38(.a(u_cla12_and36[0]), .b(u_cla12_and37[0]), .out(u_cla12_and38));
  and_gate and_gate_u_cla12_and39(.a(u_cla12_pg_logic8_and0[0]), .b(u_cla12_pg_logic10_or0[0]), .out(u_cla12_and39));
  and_gate and_gate_u_cla12_and40(.a(u_cla12_and39[0]), .b(u_cla12_pg_logic9_or0[0]), .out(u_cla12_and40));
  and_gate and_gate_u_cla12_and41(.a(u_cla12_pg_logic9_and0[0]), .b(u_cla12_pg_logic10_or0[0]), .out(u_cla12_and41));
  or_gate or_gate_u_cla12_or19(.a(u_cla12_and38[0]), .b(u_cla12_and40[0]), .out(u_cla12_or19));
  or_gate or_gate_u_cla12_or20(.a(u_cla12_or19[0]), .b(u_cla12_and41[0]), .out(u_cla12_or20));
  or_gate or_gate_u_cla12_or21(.a(u_cla12_pg_logic10_and0[0]), .b(u_cla12_or20[0]), .out(u_cla12_or21));
  pg_logic pg_logic_u_cla12_pg_logic11_out(.a(a[11]), .b(b[11]), .pg_logic_or0(u_cla12_pg_logic11_or0), .pg_logic_and0(u_cla12_pg_logic11_and0), .pg_logic_xor0(u_cla12_pg_logic11_xor0));
  xor_gate xor_gate_u_cla12_xor11(.a(u_cla12_pg_logic11_xor0[0]), .b(u_cla12_or21[0]), .out(u_cla12_xor11));
  and_gate and_gate_u_cla12_and42(.a(u_cla12_or15[0]), .b(u_cla12_pg_logic10_or0[0]), .out(u_cla12_and42));
  and_gate and_gate_u_cla12_and43(.a(u_cla12_pg_logic11_or0[0]), .b(u_cla12_pg_logic9_or0[0]), .out(u_cla12_and43));
  and_gate and_gate_u_cla12_and44(.a(u_cla12_and42[0]), .b(u_cla12_and43[0]), .out(u_cla12_and44));
  and_gate and_gate_u_cla12_and45(.a(u_cla12_and44[0]), .b(u_cla12_pg_logic8_or0[0]), .out(u_cla12_and45));
  and_gate and_gate_u_cla12_and46(.a(u_cla12_pg_logic8_and0[0]), .b(u_cla12_pg_logic10_or0[0]), .out(u_cla12_and46));
  and_gate and_gate_u_cla12_and47(.a(u_cla12_pg_logic11_or0[0]), .b(u_cla12_pg_logic9_or0[0]), .out(u_cla12_and47));
  and_gate and_gate_u_cla12_and48(.a(u_cla12_and46[0]), .b(u_cla12_and47[0]), .out(u_cla12_and48));
  and_gate and_gate_u_cla12_and49(.a(u_cla12_pg_logic9_and0[0]), .b(u_cla12_pg_logic11_or0[0]), .out(u_cla12_and49));
  and_gate and_gate_u_cla12_and50(.a(u_cla12_and49[0]), .b(u_cla12_pg_logic10_or0[0]), .out(u_cla12_and50));
  and_gate and_gate_u_cla12_and51(.a(u_cla12_pg_logic10_and0[0]), .b(u_cla12_pg_logic11_or0[0]), .out(u_cla12_and51));
  or_gate or_gate_u_cla12_or22(.a(u_cla12_and45[0]), .b(u_cla12_and50[0]), .out(u_cla12_or22));
  or_gate or_gate_u_cla12_or23(.a(u_cla12_and48[0]), .b(u_cla12_and51[0]), .out(u_cla12_or23));
  or_gate or_gate_u_cla12_or24(.a(u_cla12_or22[0]), .b(u_cla12_or23[0]), .out(u_cla12_or24));
  or_gate or_gate_u_cla12_or25(.a(u_cla12_pg_logic11_and0[0]), .b(u_cla12_or24[0]), .out(u_cla12_or25));

  assign u_cla12_out[0] = u_cla12_pg_logic0_xor0[0];
  assign u_cla12_out[1] = u_cla12_xor1[0];
  assign u_cla12_out[2] = u_cla12_xor2[0];
  assign u_cla12_out[3] = u_cla12_xor3[0];
  assign u_cla12_out[4] = u_cla12_xor4[0];
  assign u_cla12_out[5] = u_cla12_xor5[0];
  assign u_cla12_out[6] = u_cla12_xor6[0];
  assign u_cla12_out[7] = u_cla12_xor7[0];
  assign u_cla12_out[8] = u_cla12_xor8[0];
  assign u_cla12_out[9] = u_cla12_xor9[0];
  assign u_cla12_out[10] = u_cla12_xor10[0];
  assign u_cla12_out[11] = u_cla12_xor11[0];
  assign u_cla12_out[12] = u_cla12_or25[0];
endmodule

module s_csamul_cla12(input [11:0] a, input [11:0] b, output [23:0] s_csamul_cla12_out);
  wire [0:0] s_csamul_cla12_and0_0;
  wire [0:0] s_csamul_cla12_and1_0;
  wire [0:0] s_csamul_cla12_and2_0;
  wire [0:0] s_csamul_cla12_and3_0;
  wire [0:0] s_csamul_cla12_and4_0;
  wire [0:0] s_csamul_cla12_and5_0;
  wire [0:0] s_csamul_cla12_and6_0;
  wire [0:0] s_csamul_cla12_and7_0;
  wire [0:0] s_csamul_cla12_and8_0;
  wire [0:0] s_csamul_cla12_and9_0;
  wire [0:0] s_csamul_cla12_and10_0;
  wire [0:0] s_csamul_cla12_nand11_0;
  wire [0:0] s_csamul_cla12_and0_1;
  wire [0:0] s_csamul_cla12_ha0_1_xor0;
  wire [0:0] s_csamul_cla12_ha0_1_and0;
  wire [0:0] s_csamul_cla12_and1_1;
  wire [0:0] s_csamul_cla12_ha1_1_xor0;
  wire [0:0] s_csamul_cla12_ha1_1_and0;
  wire [0:0] s_csamul_cla12_and2_1;
  wire [0:0] s_csamul_cla12_ha2_1_xor0;
  wire [0:0] s_csamul_cla12_ha2_1_and0;
  wire [0:0] s_csamul_cla12_and3_1;
  wire [0:0] s_csamul_cla12_ha3_1_xor0;
  wire [0:0] s_csamul_cla12_ha3_1_and0;
  wire [0:0] s_csamul_cla12_and4_1;
  wire [0:0] s_csamul_cla12_ha4_1_xor0;
  wire [0:0] s_csamul_cla12_ha4_1_and0;
  wire [0:0] s_csamul_cla12_and5_1;
  wire [0:0] s_csamul_cla12_ha5_1_xor0;
  wire [0:0] s_csamul_cla12_ha5_1_and0;
  wire [0:0] s_csamul_cla12_and6_1;
  wire [0:0] s_csamul_cla12_ha6_1_xor0;
  wire [0:0] s_csamul_cla12_ha6_1_and0;
  wire [0:0] s_csamul_cla12_and7_1;
  wire [0:0] s_csamul_cla12_ha7_1_xor0;
  wire [0:0] s_csamul_cla12_ha7_1_and0;
  wire [0:0] s_csamul_cla12_and8_1;
  wire [0:0] s_csamul_cla12_ha8_1_xor0;
  wire [0:0] s_csamul_cla12_ha8_1_and0;
  wire [0:0] s_csamul_cla12_and9_1;
  wire [0:0] s_csamul_cla12_ha9_1_xor0;
  wire [0:0] s_csamul_cla12_ha9_1_and0;
  wire [0:0] s_csamul_cla12_and10_1;
  wire [0:0] s_csamul_cla12_ha10_1_xor0;
  wire [0:0] s_csamul_cla12_ha10_1_and0;
  wire [0:0] s_csamul_cla12_nand11_1;
  wire [0:0] s_csamul_cla12_ha11_1_xor0;
  wire [0:0] s_csamul_cla12_and0_2;
  wire [0:0] s_csamul_cla12_fa0_2_xor1;
  wire [0:0] s_csamul_cla12_fa0_2_or0;
  wire [0:0] s_csamul_cla12_and1_2;
  wire [0:0] s_csamul_cla12_fa1_2_xor1;
  wire [0:0] s_csamul_cla12_fa1_2_or0;
  wire [0:0] s_csamul_cla12_and2_2;
  wire [0:0] s_csamul_cla12_fa2_2_xor1;
  wire [0:0] s_csamul_cla12_fa2_2_or0;
  wire [0:0] s_csamul_cla12_and3_2;
  wire [0:0] s_csamul_cla12_fa3_2_xor1;
  wire [0:0] s_csamul_cla12_fa3_2_or0;
  wire [0:0] s_csamul_cla12_and4_2;
  wire [0:0] s_csamul_cla12_fa4_2_xor1;
  wire [0:0] s_csamul_cla12_fa4_2_or0;
  wire [0:0] s_csamul_cla12_and5_2;
  wire [0:0] s_csamul_cla12_fa5_2_xor1;
  wire [0:0] s_csamul_cla12_fa5_2_or0;
  wire [0:0] s_csamul_cla12_and6_2;
  wire [0:0] s_csamul_cla12_fa6_2_xor1;
  wire [0:0] s_csamul_cla12_fa6_2_or0;
  wire [0:0] s_csamul_cla12_and7_2;
  wire [0:0] s_csamul_cla12_fa7_2_xor1;
  wire [0:0] s_csamul_cla12_fa7_2_or0;
  wire [0:0] s_csamul_cla12_and8_2;
  wire [0:0] s_csamul_cla12_fa8_2_xor1;
  wire [0:0] s_csamul_cla12_fa8_2_or0;
  wire [0:0] s_csamul_cla12_and9_2;
  wire [0:0] s_csamul_cla12_fa9_2_xor1;
  wire [0:0] s_csamul_cla12_fa9_2_or0;
  wire [0:0] s_csamul_cla12_and10_2;
  wire [0:0] s_csamul_cla12_fa10_2_xor1;
  wire [0:0] s_csamul_cla12_fa10_2_or0;
  wire [0:0] s_csamul_cla12_nand11_2;
  wire [0:0] s_csamul_cla12_ha11_2_xor0;
  wire [0:0] s_csamul_cla12_ha11_2_and0;
  wire [0:0] s_csamul_cla12_and0_3;
  wire [0:0] s_csamul_cla12_fa0_3_xor1;
  wire [0:0] s_csamul_cla12_fa0_3_or0;
  wire [0:0] s_csamul_cla12_and1_3;
  wire [0:0] s_csamul_cla12_fa1_3_xor1;
  wire [0:0] s_csamul_cla12_fa1_3_or0;
  wire [0:0] s_csamul_cla12_and2_3;
  wire [0:0] s_csamul_cla12_fa2_3_xor1;
  wire [0:0] s_csamul_cla12_fa2_3_or0;
  wire [0:0] s_csamul_cla12_and3_3;
  wire [0:0] s_csamul_cla12_fa3_3_xor1;
  wire [0:0] s_csamul_cla12_fa3_3_or0;
  wire [0:0] s_csamul_cla12_and4_3;
  wire [0:0] s_csamul_cla12_fa4_3_xor1;
  wire [0:0] s_csamul_cla12_fa4_3_or0;
  wire [0:0] s_csamul_cla12_and5_3;
  wire [0:0] s_csamul_cla12_fa5_3_xor1;
  wire [0:0] s_csamul_cla12_fa5_3_or0;
  wire [0:0] s_csamul_cla12_and6_3;
  wire [0:0] s_csamul_cla12_fa6_3_xor1;
  wire [0:0] s_csamul_cla12_fa6_3_or0;
  wire [0:0] s_csamul_cla12_and7_3;
  wire [0:0] s_csamul_cla12_fa7_3_xor1;
  wire [0:0] s_csamul_cla12_fa7_3_or0;
  wire [0:0] s_csamul_cla12_and8_3;
  wire [0:0] s_csamul_cla12_fa8_3_xor1;
  wire [0:0] s_csamul_cla12_fa8_3_or0;
  wire [0:0] s_csamul_cla12_and9_3;
  wire [0:0] s_csamul_cla12_fa9_3_xor1;
  wire [0:0] s_csamul_cla12_fa9_3_or0;
  wire [0:0] s_csamul_cla12_and10_3;
  wire [0:0] s_csamul_cla12_fa10_3_xor1;
  wire [0:0] s_csamul_cla12_fa10_3_or0;
  wire [0:0] s_csamul_cla12_nand11_3;
  wire [0:0] s_csamul_cla12_ha11_3_xor0;
  wire [0:0] s_csamul_cla12_ha11_3_and0;
  wire [0:0] s_csamul_cla12_and0_4;
  wire [0:0] s_csamul_cla12_fa0_4_xor1;
  wire [0:0] s_csamul_cla12_fa0_4_or0;
  wire [0:0] s_csamul_cla12_and1_4;
  wire [0:0] s_csamul_cla12_fa1_4_xor1;
  wire [0:0] s_csamul_cla12_fa1_4_or0;
  wire [0:0] s_csamul_cla12_and2_4;
  wire [0:0] s_csamul_cla12_fa2_4_xor1;
  wire [0:0] s_csamul_cla12_fa2_4_or0;
  wire [0:0] s_csamul_cla12_and3_4;
  wire [0:0] s_csamul_cla12_fa3_4_xor1;
  wire [0:0] s_csamul_cla12_fa3_4_or0;
  wire [0:0] s_csamul_cla12_and4_4;
  wire [0:0] s_csamul_cla12_fa4_4_xor1;
  wire [0:0] s_csamul_cla12_fa4_4_or0;
  wire [0:0] s_csamul_cla12_and5_4;
  wire [0:0] s_csamul_cla12_fa5_4_xor1;
  wire [0:0] s_csamul_cla12_fa5_4_or0;
  wire [0:0] s_csamul_cla12_and6_4;
  wire [0:0] s_csamul_cla12_fa6_4_xor1;
  wire [0:0] s_csamul_cla12_fa6_4_or0;
  wire [0:0] s_csamul_cla12_and7_4;
  wire [0:0] s_csamul_cla12_fa7_4_xor1;
  wire [0:0] s_csamul_cla12_fa7_4_or0;
  wire [0:0] s_csamul_cla12_and8_4;
  wire [0:0] s_csamul_cla12_fa8_4_xor1;
  wire [0:0] s_csamul_cla12_fa8_4_or0;
  wire [0:0] s_csamul_cla12_and9_4;
  wire [0:0] s_csamul_cla12_fa9_4_xor1;
  wire [0:0] s_csamul_cla12_fa9_4_or0;
  wire [0:0] s_csamul_cla12_and10_4;
  wire [0:0] s_csamul_cla12_fa10_4_xor1;
  wire [0:0] s_csamul_cla12_fa10_4_or0;
  wire [0:0] s_csamul_cla12_nand11_4;
  wire [0:0] s_csamul_cla12_ha11_4_xor0;
  wire [0:0] s_csamul_cla12_ha11_4_and0;
  wire [0:0] s_csamul_cla12_and0_5;
  wire [0:0] s_csamul_cla12_fa0_5_xor1;
  wire [0:0] s_csamul_cla12_fa0_5_or0;
  wire [0:0] s_csamul_cla12_and1_5;
  wire [0:0] s_csamul_cla12_fa1_5_xor1;
  wire [0:0] s_csamul_cla12_fa1_5_or0;
  wire [0:0] s_csamul_cla12_and2_5;
  wire [0:0] s_csamul_cla12_fa2_5_xor1;
  wire [0:0] s_csamul_cla12_fa2_5_or0;
  wire [0:0] s_csamul_cla12_and3_5;
  wire [0:0] s_csamul_cla12_fa3_5_xor1;
  wire [0:0] s_csamul_cla12_fa3_5_or0;
  wire [0:0] s_csamul_cla12_and4_5;
  wire [0:0] s_csamul_cla12_fa4_5_xor1;
  wire [0:0] s_csamul_cla12_fa4_5_or0;
  wire [0:0] s_csamul_cla12_and5_5;
  wire [0:0] s_csamul_cla12_fa5_5_xor1;
  wire [0:0] s_csamul_cla12_fa5_5_or0;
  wire [0:0] s_csamul_cla12_and6_5;
  wire [0:0] s_csamul_cla12_fa6_5_xor1;
  wire [0:0] s_csamul_cla12_fa6_5_or0;
  wire [0:0] s_csamul_cla12_and7_5;
  wire [0:0] s_csamul_cla12_fa7_5_xor1;
  wire [0:0] s_csamul_cla12_fa7_5_or0;
  wire [0:0] s_csamul_cla12_and8_5;
  wire [0:0] s_csamul_cla12_fa8_5_xor1;
  wire [0:0] s_csamul_cla12_fa8_5_or0;
  wire [0:0] s_csamul_cla12_and9_5;
  wire [0:0] s_csamul_cla12_fa9_5_xor1;
  wire [0:0] s_csamul_cla12_fa9_5_or0;
  wire [0:0] s_csamul_cla12_and10_5;
  wire [0:0] s_csamul_cla12_fa10_5_xor1;
  wire [0:0] s_csamul_cla12_fa10_5_or0;
  wire [0:0] s_csamul_cla12_nand11_5;
  wire [0:0] s_csamul_cla12_ha11_5_xor0;
  wire [0:0] s_csamul_cla12_ha11_5_and0;
  wire [0:0] s_csamul_cla12_and0_6;
  wire [0:0] s_csamul_cla12_fa0_6_xor1;
  wire [0:0] s_csamul_cla12_fa0_6_or0;
  wire [0:0] s_csamul_cla12_and1_6;
  wire [0:0] s_csamul_cla12_fa1_6_xor1;
  wire [0:0] s_csamul_cla12_fa1_6_or0;
  wire [0:0] s_csamul_cla12_and2_6;
  wire [0:0] s_csamul_cla12_fa2_6_xor1;
  wire [0:0] s_csamul_cla12_fa2_6_or0;
  wire [0:0] s_csamul_cla12_and3_6;
  wire [0:0] s_csamul_cla12_fa3_6_xor1;
  wire [0:0] s_csamul_cla12_fa3_6_or0;
  wire [0:0] s_csamul_cla12_and4_6;
  wire [0:0] s_csamul_cla12_fa4_6_xor1;
  wire [0:0] s_csamul_cla12_fa4_6_or0;
  wire [0:0] s_csamul_cla12_and5_6;
  wire [0:0] s_csamul_cla12_fa5_6_xor1;
  wire [0:0] s_csamul_cla12_fa5_6_or0;
  wire [0:0] s_csamul_cla12_and6_6;
  wire [0:0] s_csamul_cla12_fa6_6_xor1;
  wire [0:0] s_csamul_cla12_fa6_6_or0;
  wire [0:0] s_csamul_cla12_and7_6;
  wire [0:0] s_csamul_cla12_fa7_6_xor1;
  wire [0:0] s_csamul_cla12_fa7_6_or0;
  wire [0:0] s_csamul_cla12_and8_6;
  wire [0:0] s_csamul_cla12_fa8_6_xor1;
  wire [0:0] s_csamul_cla12_fa8_6_or0;
  wire [0:0] s_csamul_cla12_and9_6;
  wire [0:0] s_csamul_cla12_fa9_6_xor1;
  wire [0:0] s_csamul_cla12_fa9_6_or0;
  wire [0:0] s_csamul_cla12_and10_6;
  wire [0:0] s_csamul_cla12_fa10_6_xor1;
  wire [0:0] s_csamul_cla12_fa10_6_or0;
  wire [0:0] s_csamul_cla12_nand11_6;
  wire [0:0] s_csamul_cla12_ha11_6_xor0;
  wire [0:0] s_csamul_cla12_ha11_6_and0;
  wire [0:0] s_csamul_cla12_and0_7;
  wire [0:0] s_csamul_cla12_fa0_7_xor1;
  wire [0:0] s_csamul_cla12_fa0_7_or0;
  wire [0:0] s_csamul_cla12_and1_7;
  wire [0:0] s_csamul_cla12_fa1_7_xor1;
  wire [0:0] s_csamul_cla12_fa1_7_or0;
  wire [0:0] s_csamul_cla12_and2_7;
  wire [0:0] s_csamul_cla12_fa2_7_xor1;
  wire [0:0] s_csamul_cla12_fa2_7_or0;
  wire [0:0] s_csamul_cla12_and3_7;
  wire [0:0] s_csamul_cla12_fa3_7_xor1;
  wire [0:0] s_csamul_cla12_fa3_7_or0;
  wire [0:0] s_csamul_cla12_and4_7;
  wire [0:0] s_csamul_cla12_fa4_7_xor1;
  wire [0:0] s_csamul_cla12_fa4_7_or0;
  wire [0:0] s_csamul_cla12_and5_7;
  wire [0:0] s_csamul_cla12_fa5_7_xor1;
  wire [0:0] s_csamul_cla12_fa5_7_or0;
  wire [0:0] s_csamul_cla12_and6_7;
  wire [0:0] s_csamul_cla12_fa6_7_xor1;
  wire [0:0] s_csamul_cla12_fa6_7_or0;
  wire [0:0] s_csamul_cla12_and7_7;
  wire [0:0] s_csamul_cla12_fa7_7_xor1;
  wire [0:0] s_csamul_cla12_fa7_7_or0;
  wire [0:0] s_csamul_cla12_and8_7;
  wire [0:0] s_csamul_cla12_fa8_7_xor1;
  wire [0:0] s_csamul_cla12_fa8_7_or0;
  wire [0:0] s_csamul_cla12_and9_7;
  wire [0:0] s_csamul_cla12_fa9_7_xor1;
  wire [0:0] s_csamul_cla12_fa9_7_or0;
  wire [0:0] s_csamul_cla12_and10_7;
  wire [0:0] s_csamul_cla12_fa10_7_xor1;
  wire [0:0] s_csamul_cla12_fa10_7_or0;
  wire [0:0] s_csamul_cla12_nand11_7;
  wire [0:0] s_csamul_cla12_ha11_7_xor0;
  wire [0:0] s_csamul_cla12_ha11_7_and0;
  wire [0:0] s_csamul_cla12_and0_8;
  wire [0:0] s_csamul_cla12_fa0_8_xor1;
  wire [0:0] s_csamul_cla12_fa0_8_or0;
  wire [0:0] s_csamul_cla12_and1_8;
  wire [0:0] s_csamul_cla12_fa1_8_xor1;
  wire [0:0] s_csamul_cla12_fa1_8_or0;
  wire [0:0] s_csamul_cla12_and2_8;
  wire [0:0] s_csamul_cla12_fa2_8_xor1;
  wire [0:0] s_csamul_cla12_fa2_8_or0;
  wire [0:0] s_csamul_cla12_and3_8;
  wire [0:0] s_csamul_cla12_fa3_8_xor1;
  wire [0:0] s_csamul_cla12_fa3_8_or0;
  wire [0:0] s_csamul_cla12_and4_8;
  wire [0:0] s_csamul_cla12_fa4_8_xor1;
  wire [0:0] s_csamul_cla12_fa4_8_or0;
  wire [0:0] s_csamul_cla12_and5_8;
  wire [0:0] s_csamul_cla12_fa5_8_xor1;
  wire [0:0] s_csamul_cla12_fa5_8_or0;
  wire [0:0] s_csamul_cla12_and6_8;
  wire [0:0] s_csamul_cla12_fa6_8_xor1;
  wire [0:0] s_csamul_cla12_fa6_8_or0;
  wire [0:0] s_csamul_cla12_and7_8;
  wire [0:0] s_csamul_cla12_fa7_8_xor1;
  wire [0:0] s_csamul_cla12_fa7_8_or0;
  wire [0:0] s_csamul_cla12_and8_8;
  wire [0:0] s_csamul_cla12_fa8_8_xor1;
  wire [0:0] s_csamul_cla12_fa8_8_or0;
  wire [0:0] s_csamul_cla12_and9_8;
  wire [0:0] s_csamul_cla12_fa9_8_xor1;
  wire [0:0] s_csamul_cla12_fa9_8_or0;
  wire [0:0] s_csamul_cla12_and10_8;
  wire [0:0] s_csamul_cla12_fa10_8_xor1;
  wire [0:0] s_csamul_cla12_fa10_8_or0;
  wire [0:0] s_csamul_cla12_nand11_8;
  wire [0:0] s_csamul_cla12_ha11_8_xor0;
  wire [0:0] s_csamul_cla12_ha11_8_and0;
  wire [0:0] s_csamul_cla12_and0_9;
  wire [0:0] s_csamul_cla12_fa0_9_xor1;
  wire [0:0] s_csamul_cla12_fa0_9_or0;
  wire [0:0] s_csamul_cla12_and1_9;
  wire [0:0] s_csamul_cla12_fa1_9_xor1;
  wire [0:0] s_csamul_cla12_fa1_9_or0;
  wire [0:0] s_csamul_cla12_and2_9;
  wire [0:0] s_csamul_cla12_fa2_9_xor1;
  wire [0:0] s_csamul_cla12_fa2_9_or0;
  wire [0:0] s_csamul_cla12_and3_9;
  wire [0:0] s_csamul_cla12_fa3_9_xor1;
  wire [0:0] s_csamul_cla12_fa3_9_or0;
  wire [0:0] s_csamul_cla12_and4_9;
  wire [0:0] s_csamul_cla12_fa4_9_xor1;
  wire [0:0] s_csamul_cla12_fa4_9_or0;
  wire [0:0] s_csamul_cla12_and5_9;
  wire [0:0] s_csamul_cla12_fa5_9_xor1;
  wire [0:0] s_csamul_cla12_fa5_9_or0;
  wire [0:0] s_csamul_cla12_and6_9;
  wire [0:0] s_csamul_cla12_fa6_9_xor1;
  wire [0:0] s_csamul_cla12_fa6_9_or0;
  wire [0:0] s_csamul_cla12_and7_9;
  wire [0:0] s_csamul_cla12_fa7_9_xor1;
  wire [0:0] s_csamul_cla12_fa7_9_or0;
  wire [0:0] s_csamul_cla12_and8_9;
  wire [0:0] s_csamul_cla12_fa8_9_xor1;
  wire [0:0] s_csamul_cla12_fa8_9_or0;
  wire [0:0] s_csamul_cla12_and9_9;
  wire [0:0] s_csamul_cla12_fa9_9_xor1;
  wire [0:0] s_csamul_cla12_fa9_9_or0;
  wire [0:0] s_csamul_cla12_and10_9;
  wire [0:0] s_csamul_cla12_fa10_9_xor1;
  wire [0:0] s_csamul_cla12_fa10_9_or0;
  wire [0:0] s_csamul_cla12_nand11_9;
  wire [0:0] s_csamul_cla12_ha11_9_xor0;
  wire [0:0] s_csamul_cla12_ha11_9_and0;
  wire [0:0] s_csamul_cla12_and0_10;
  wire [0:0] s_csamul_cla12_fa0_10_xor1;
  wire [0:0] s_csamul_cla12_fa0_10_or0;
  wire [0:0] s_csamul_cla12_and1_10;
  wire [0:0] s_csamul_cla12_fa1_10_xor1;
  wire [0:0] s_csamul_cla12_fa1_10_or0;
  wire [0:0] s_csamul_cla12_and2_10;
  wire [0:0] s_csamul_cla12_fa2_10_xor1;
  wire [0:0] s_csamul_cla12_fa2_10_or0;
  wire [0:0] s_csamul_cla12_and3_10;
  wire [0:0] s_csamul_cla12_fa3_10_xor1;
  wire [0:0] s_csamul_cla12_fa3_10_or0;
  wire [0:0] s_csamul_cla12_and4_10;
  wire [0:0] s_csamul_cla12_fa4_10_xor1;
  wire [0:0] s_csamul_cla12_fa4_10_or0;
  wire [0:0] s_csamul_cla12_and5_10;
  wire [0:0] s_csamul_cla12_fa5_10_xor1;
  wire [0:0] s_csamul_cla12_fa5_10_or0;
  wire [0:0] s_csamul_cla12_and6_10;
  wire [0:0] s_csamul_cla12_fa6_10_xor1;
  wire [0:0] s_csamul_cla12_fa6_10_or0;
  wire [0:0] s_csamul_cla12_and7_10;
  wire [0:0] s_csamul_cla12_fa7_10_xor1;
  wire [0:0] s_csamul_cla12_fa7_10_or0;
  wire [0:0] s_csamul_cla12_and8_10;
  wire [0:0] s_csamul_cla12_fa8_10_xor1;
  wire [0:0] s_csamul_cla12_fa8_10_or0;
  wire [0:0] s_csamul_cla12_and9_10;
  wire [0:0] s_csamul_cla12_fa9_10_xor1;
  wire [0:0] s_csamul_cla12_fa9_10_or0;
  wire [0:0] s_csamul_cla12_and10_10;
  wire [0:0] s_csamul_cla12_fa10_10_xor1;
  wire [0:0] s_csamul_cla12_fa10_10_or0;
  wire [0:0] s_csamul_cla12_nand11_10;
  wire [0:0] s_csamul_cla12_ha11_10_xor0;
  wire [0:0] s_csamul_cla12_ha11_10_and0;
  wire [0:0] s_csamul_cla12_nand0_11;
  wire [0:0] s_csamul_cla12_fa0_11_xor1;
  wire [0:0] s_csamul_cla12_fa0_11_or0;
  wire [0:0] s_csamul_cla12_nand1_11;
  wire [0:0] s_csamul_cla12_fa1_11_xor1;
  wire [0:0] s_csamul_cla12_fa1_11_or0;
  wire [0:0] s_csamul_cla12_nand2_11;
  wire [0:0] s_csamul_cla12_fa2_11_xor1;
  wire [0:0] s_csamul_cla12_fa2_11_or0;
  wire [0:0] s_csamul_cla12_nand3_11;
  wire [0:0] s_csamul_cla12_fa3_11_xor1;
  wire [0:0] s_csamul_cla12_fa3_11_or0;
  wire [0:0] s_csamul_cla12_nand4_11;
  wire [0:0] s_csamul_cla12_fa4_11_xor1;
  wire [0:0] s_csamul_cla12_fa4_11_or0;
  wire [0:0] s_csamul_cla12_nand5_11;
  wire [0:0] s_csamul_cla12_fa5_11_xor1;
  wire [0:0] s_csamul_cla12_fa5_11_or0;
  wire [0:0] s_csamul_cla12_nand6_11;
  wire [0:0] s_csamul_cla12_fa6_11_xor1;
  wire [0:0] s_csamul_cla12_fa6_11_or0;
  wire [0:0] s_csamul_cla12_nand7_11;
  wire [0:0] s_csamul_cla12_fa7_11_xor1;
  wire [0:0] s_csamul_cla12_fa7_11_or0;
  wire [0:0] s_csamul_cla12_nand8_11;
  wire [0:0] s_csamul_cla12_fa8_11_xor1;
  wire [0:0] s_csamul_cla12_fa8_11_or0;
  wire [0:0] s_csamul_cla12_nand9_11;
  wire [0:0] s_csamul_cla12_fa9_11_xor1;
  wire [0:0] s_csamul_cla12_fa9_11_or0;
  wire [0:0] s_csamul_cla12_nand10_11;
  wire [0:0] s_csamul_cla12_fa10_11_xor1;
  wire [0:0] s_csamul_cla12_fa10_11_or0;
  wire [0:0] s_csamul_cla12_and11_11;
  wire [0:0] s_csamul_cla12_ha11_11_xor0;
  wire [0:0] s_csamul_cla12_ha11_11_and0;
  wire [11:0] s_csamul_cla12_u_cla12_a;
  wire [11:0] s_csamul_cla12_u_cla12_b;
  wire [12:0] s_csamul_cla12_u_cla12_out;

  and_gate and_gate_s_csamul_cla12_and0_0(.a(a[0]), .b(b[0]), .out(s_csamul_cla12_and0_0));
  and_gate and_gate_s_csamul_cla12_and1_0(.a(a[1]), .b(b[0]), .out(s_csamul_cla12_and1_0));
  and_gate and_gate_s_csamul_cla12_and2_0(.a(a[2]), .b(b[0]), .out(s_csamul_cla12_and2_0));
  and_gate and_gate_s_csamul_cla12_and3_0(.a(a[3]), .b(b[0]), .out(s_csamul_cla12_and3_0));
  and_gate and_gate_s_csamul_cla12_and4_0(.a(a[4]), .b(b[0]), .out(s_csamul_cla12_and4_0));
  and_gate and_gate_s_csamul_cla12_and5_0(.a(a[5]), .b(b[0]), .out(s_csamul_cla12_and5_0));
  and_gate and_gate_s_csamul_cla12_and6_0(.a(a[6]), .b(b[0]), .out(s_csamul_cla12_and6_0));
  and_gate and_gate_s_csamul_cla12_and7_0(.a(a[7]), .b(b[0]), .out(s_csamul_cla12_and7_0));
  and_gate and_gate_s_csamul_cla12_and8_0(.a(a[8]), .b(b[0]), .out(s_csamul_cla12_and8_0));
  and_gate and_gate_s_csamul_cla12_and9_0(.a(a[9]), .b(b[0]), .out(s_csamul_cla12_and9_0));
  and_gate and_gate_s_csamul_cla12_and10_0(.a(a[10]), .b(b[0]), .out(s_csamul_cla12_and10_0));
  nand_gate nand_gate_s_csamul_cla12_nand11_0(.a(a[11]), .b(b[0]), .out(s_csamul_cla12_nand11_0));
  and_gate and_gate_s_csamul_cla12_and0_1(.a(a[0]), .b(b[1]), .out(s_csamul_cla12_and0_1));
  ha ha_s_csamul_cla12_ha0_1_out(.a(s_csamul_cla12_and0_1[0]), .b(s_csamul_cla12_and1_0[0]), .ha_xor0(s_csamul_cla12_ha0_1_xor0), .ha_and0(s_csamul_cla12_ha0_1_and0));
  and_gate and_gate_s_csamul_cla12_and1_1(.a(a[1]), .b(b[1]), .out(s_csamul_cla12_and1_1));
  ha ha_s_csamul_cla12_ha1_1_out(.a(s_csamul_cla12_and1_1[0]), .b(s_csamul_cla12_and2_0[0]), .ha_xor0(s_csamul_cla12_ha1_1_xor0), .ha_and0(s_csamul_cla12_ha1_1_and0));
  and_gate and_gate_s_csamul_cla12_and2_1(.a(a[2]), .b(b[1]), .out(s_csamul_cla12_and2_1));
  ha ha_s_csamul_cla12_ha2_1_out(.a(s_csamul_cla12_and2_1[0]), .b(s_csamul_cla12_and3_0[0]), .ha_xor0(s_csamul_cla12_ha2_1_xor0), .ha_and0(s_csamul_cla12_ha2_1_and0));
  and_gate and_gate_s_csamul_cla12_and3_1(.a(a[3]), .b(b[1]), .out(s_csamul_cla12_and3_1));
  ha ha_s_csamul_cla12_ha3_1_out(.a(s_csamul_cla12_and3_1[0]), .b(s_csamul_cla12_and4_0[0]), .ha_xor0(s_csamul_cla12_ha3_1_xor0), .ha_and0(s_csamul_cla12_ha3_1_and0));
  and_gate and_gate_s_csamul_cla12_and4_1(.a(a[4]), .b(b[1]), .out(s_csamul_cla12_and4_1));
  ha ha_s_csamul_cla12_ha4_1_out(.a(s_csamul_cla12_and4_1[0]), .b(s_csamul_cla12_and5_0[0]), .ha_xor0(s_csamul_cla12_ha4_1_xor0), .ha_and0(s_csamul_cla12_ha4_1_and0));
  and_gate and_gate_s_csamul_cla12_and5_1(.a(a[5]), .b(b[1]), .out(s_csamul_cla12_and5_1));
  ha ha_s_csamul_cla12_ha5_1_out(.a(s_csamul_cla12_and5_1[0]), .b(s_csamul_cla12_and6_0[0]), .ha_xor0(s_csamul_cla12_ha5_1_xor0), .ha_and0(s_csamul_cla12_ha5_1_and0));
  and_gate and_gate_s_csamul_cla12_and6_1(.a(a[6]), .b(b[1]), .out(s_csamul_cla12_and6_1));
  ha ha_s_csamul_cla12_ha6_1_out(.a(s_csamul_cla12_and6_1[0]), .b(s_csamul_cla12_and7_0[0]), .ha_xor0(s_csamul_cla12_ha6_1_xor0), .ha_and0(s_csamul_cla12_ha6_1_and0));
  and_gate and_gate_s_csamul_cla12_and7_1(.a(a[7]), .b(b[1]), .out(s_csamul_cla12_and7_1));
  ha ha_s_csamul_cla12_ha7_1_out(.a(s_csamul_cla12_and7_1[0]), .b(s_csamul_cla12_and8_0[0]), .ha_xor0(s_csamul_cla12_ha7_1_xor0), .ha_and0(s_csamul_cla12_ha7_1_and0));
  and_gate and_gate_s_csamul_cla12_and8_1(.a(a[8]), .b(b[1]), .out(s_csamul_cla12_and8_1));
  ha ha_s_csamul_cla12_ha8_1_out(.a(s_csamul_cla12_and8_1[0]), .b(s_csamul_cla12_and9_0[0]), .ha_xor0(s_csamul_cla12_ha8_1_xor0), .ha_and0(s_csamul_cla12_ha8_1_and0));
  and_gate and_gate_s_csamul_cla12_and9_1(.a(a[9]), .b(b[1]), .out(s_csamul_cla12_and9_1));
  ha ha_s_csamul_cla12_ha9_1_out(.a(s_csamul_cla12_and9_1[0]), .b(s_csamul_cla12_and10_0[0]), .ha_xor0(s_csamul_cla12_ha9_1_xor0), .ha_and0(s_csamul_cla12_ha9_1_and0));
  and_gate and_gate_s_csamul_cla12_and10_1(.a(a[10]), .b(b[1]), .out(s_csamul_cla12_and10_1));
  ha ha_s_csamul_cla12_ha10_1_out(.a(s_csamul_cla12_and10_1[0]), .b(s_csamul_cla12_nand11_0[0]), .ha_xor0(s_csamul_cla12_ha10_1_xor0), .ha_and0(s_csamul_cla12_ha10_1_and0));
  nand_gate nand_gate_s_csamul_cla12_nand11_1(.a(a[11]), .b(b[1]), .out(s_csamul_cla12_nand11_1));
  ha ha_s_csamul_cla12_ha11_1_out(.a(s_csamul_cla12_nand11_1[0]), .b(1'b1), .ha_xor0(s_csamul_cla12_ha11_1_xor0), .ha_and0(s_csamul_cla12_nand11_1));
  and_gate and_gate_s_csamul_cla12_and0_2(.a(a[0]), .b(b[2]), .out(s_csamul_cla12_and0_2));
  fa fa_s_csamul_cla12_fa0_2_out(.a(s_csamul_cla12_and0_2[0]), .b(s_csamul_cla12_ha1_1_xor0[0]), .cin(s_csamul_cla12_ha0_1_and0[0]), .fa_xor1(s_csamul_cla12_fa0_2_xor1), .fa_or0(s_csamul_cla12_fa0_2_or0));
  and_gate and_gate_s_csamul_cla12_and1_2(.a(a[1]), .b(b[2]), .out(s_csamul_cla12_and1_2));
  fa fa_s_csamul_cla12_fa1_2_out(.a(s_csamul_cla12_and1_2[0]), .b(s_csamul_cla12_ha2_1_xor0[0]), .cin(s_csamul_cla12_ha1_1_and0[0]), .fa_xor1(s_csamul_cla12_fa1_2_xor1), .fa_or0(s_csamul_cla12_fa1_2_or0));
  and_gate and_gate_s_csamul_cla12_and2_2(.a(a[2]), .b(b[2]), .out(s_csamul_cla12_and2_2));
  fa fa_s_csamul_cla12_fa2_2_out(.a(s_csamul_cla12_and2_2[0]), .b(s_csamul_cla12_ha3_1_xor0[0]), .cin(s_csamul_cla12_ha2_1_and0[0]), .fa_xor1(s_csamul_cla12_fa2_2_xor1), .fa_or0(s_csamul_cla12_fa2_2_or0));
  and_gate and_gate_s_csamul_cla12_and3_2(.a(a[3]), .b(b[2]), .out(s_csamul_cla12_and3_2));
  fa fa_s_csamul_cla12_fa3_2_out(.a(s_csamul_cla12_and3_2[0]), .b(s_csamul_cla12_ha4_1_xor0[0]), .cin(s_csamul_cla12_ha3_1_and0[0]), .fa_xor1(s_csamul_cla12_fa3_2_xor1), .fa_or0(s_csamul_cla12_fa3_2_or0));
  and_gate and_gate_s_csamul_cla12_and4_2(.a(a[4]), .b(b[2]), .out(s_csamul_cla12_and4_2));
  fa fa_s_csamul_cla12_fa4_2_out(.a(s_csamul_cla12_and4_2[0]), .b(s_csamul_cla12_ha5_1_xor0[0]), .cin(s_csamul_cla12_ha4_1_and0[0]), .fa_xor1(s_csamul_cla12_fa4_2_xor1), .fa_or0(s_csamul_cla12_fa4_2_or0));
  and_gate and_gate_s_csamul_cla12_and5_2(.a(a[5]), .b(b[2]), .out(s_csamul_cla12_and5_2));
  fa fa_s_csamul_cla12_fa5_2_out(.a(s_csamul_cla12_and5_2[0]), .b(s_csamul_cla12_ha6_1_xor0[0]), .cin(s_csamul_cla12_ha5_1_and0[0]), .fa_xor1(s_csamul_cla12_fa5_2_xor1), .fa_or0(s_csamul_cla12_fa5_2_or0));
  and_gate and_gate_s_csamul_cla12_and6_2(.a(a[6]), .b(b[2]), .out(s_csamul_cla12_and6_2));
  fa fa_s_csamul_cla12_fa6_2_out(.a(s_csamul_cla12_and6_2[0]), .b(s_csamul_cla12_ha7_1_xor0[0]), .cin(s_csamul_cla12_ha6_1_and0[0]), .fa_xor1(s_csamul_cla12_fa6_2_xor1), .fa_or0(s_csamul_cla12_fa6_2_or0));
  and_gate and_gate_s_csamul_cla12_and7_2(.a(a[7]), .b(b[2]), .out(s_csamul_cla12_and7_2));
  fa fa_s_csamul_cla12_fa7_2_out(.a(s_csamul_cla12_and7_2[0]), .b(s_csamul_cla12_ha8_1_xor0[0]), .cin(s_csamul_cla12_ha7_1_and0[0]), .fa_xor1(s_csamul_cla12_fa7_2_xor1), .fa_or0(s_csamul_cla12_fa7_2_or0));
  and_gate and_gate_s_csamul_cla12_and8_2(.a(a[8]), .b(b[2]), .out(s_csamul_cla12_and8_2));
  fa fa_s_csamul_cla12_fa8_2_out(.a(s_csamul_cla12_and8_2[0]), .b(s_csamul_cla12_ha9_1_xor0[0]), .cin(s_csamul_cla12_ha8_1_and0[0]), .fa_xor1(s_csamul_cla12_fa8_2_xor1), .fa_or0(s_csamul_cla12_fa8_2_or0));
  and_gate and_gate_s_csamul_cla12_and9_2(.a(a[9]), .b(b[2]), .out(s_csamul_cla12_and9_2));
  fa fa_s_csamul_cla12_fa9_2_out(.a(s_csamul_cla12_and9_2[0]), .b(s_csamul_cla12_ha10_1_xor0[0]), .cin(s_csamul_cla12_ha9_1_and0[0]), .fa_xor1(s_csamul_cla12_fa9_2_xor1), .fa_or0(s_csamul_cla12_fa9_2_or0));
  and_gate and_gate_s_csamul_cla12_and10_2(.a(a[10]), .b(b[2]), .out(s_csamul_cla12_and10_2));
  fa fa_s_csamul_cla12_fa10_2_out(.a(s_csamul_cla12_and10_2[0]), .b(s_csamul_cla12_ha11_1_xor0[0]), .cin(s_csamul_cla12_ha10_1_and0[0]), .fa_xor1(s_csamul_cla12_fa10_2_xor1), .fa_or0(s_csamul_cla12_fa10_2_or0));
  nand_gate nand_gate_s_csamul_cla12_nand11_2(.a(a[11]), .b(b[2]), .out(s_csamul_cla12_nand11_2));
  ha ha_s_csamul_cla12_ha11_2_out(.a(s_csamul_cla12_nand11_2[0]), .b(s_csamul_cla12_nand11_1[0]), .ha_xor0(s_csamul_cla12_ha11_2_xor0), .ha_and0(s_csamul_cla12_ha11_2_and0));
  and_gate and_gate_s_csamul_cla12_and0_3(.a(a[0]), .b(b[3]), .out(s_csamul_cla12_and0_3));
  fa fa_s_csamul_cla12_fa0_3_out(.a(s_csamul_cla12_and0_3[0]), .b(s_csamul_cla12_fa1_2_xor1[0]), .cin(s_csamul_cla12_fa0_2_or0[0]), .fa_xor1(s_csamul_cla12_fa0_3_xor1), .fa_or0(s_csamul_cla12_fa0_3_or0));
  and_gate and_gate_s_csamul_cla12_and1_3(.a(a[1]), .b(b[3]), .out(s_csamul_cla12_and1_3));
  fa fa_s_csamul_cla12_fa1_3_out(.a(s_csamul_cla12_and1_3[0]), .b(s_csamul_cla12_fa2_2_xor1[0]), .cin(s_csamul_cla12_fa1_2_or0[0]), .fa_xor1(s_csamul_cla12_fa1_3_xor1), .fa_or0(s_csamul_cla12_fa1_3_or0));
  and_gate and_gate_s_csamul_cla12_and2_3(.a(a[2]), .b(b[3]), .out(s_csamul_cla12_and2_3));
  fa fa_s_csamul_cla12_fa2_3_out(.a(s_csamul_cla12_and2_3[0]), .b(s_csamul_cla12_fa3_2_xor1[0]), .cin(s_csamul_cla12_fa2_2_or0[0]), .fa_xor1(s_csamul_cla12_fa2_3_xor1), .fa_or0(s_csamul_cla12_fa2_3_or0));
  and_gate and_gate_s_csamul_cla12_and3_3(.a(a[3]), .b(b[3]), .out(s_csamul_cla12_and3_3));
  fa fa_s_csamul_cla12_fa3_3_out(.a(s_csamul_cla12_and3_3[0]), .b(s_csamul_cla12_fa4_2_xor1[0]), .cin(s_csamul_cla12_fa3_2_or0[0]), .fa_xor1(s_csamul_cla12_fa3_3_xor1), .fa_or0(s_csamul_cla12_fa3_3_or0));
  and_gate and_gate_s_csamul_cla12_and4_3(.a(a[4]), .b(b[3]), .out(s_csamul_cla12_and4_3));
  fa fa_s_csamul_cla12_fa4_3_out(.a(s_csamul_cla12_and4_3[0]), .b(s_csamul_cla12_fa5_2_xor1[0]), .cin(s_csamul_cla12_fa4_2_or0[0]), .fa_xor1(s_csamul_cla12_fa4_3_xor1), .fa_or0(s_csamul_cla12_fa4_3_or0));
  and_gate and_gate_s_csamul_cla12_and5_3(.a(a[5]), .b(b[3]), .out(s_csamul_cla12_and5_3));
  fa fa_s_csamul_cla12_fa5_3_out(.a(s_csamul_cla12_and5_3[0]), .b(s_csamul_cla12_fa6_2_xor1[0]), .cin(s_csamul_cla12_fa5_2_or0[0]), .fa_xor1(s_csamul_cla12_fa5_3_xor1), .fa_or0(s_csamul_cla12_fa5_3_or0));
  and_gate and_gate_s_csamul_cla12_and6_3(.a(a[6]), .b(b[3]), .out(s_csamul_cla12_and6_3));
  fa fa_s_csamul_cla12_fa6_3_out(.a(s_csamul_cla12_and6_3[0]), .b(s_csamul_cla12_fa7_2_xor1[0]), .cin(s_csamul_cla12_fa6_2_or0[0]), .fa_xor1(s_csamul_cla12_fa6_3_xor1), .fa_or0(s_csamul_cla12_fa6_3_or0));
  and_gate and_gate_s_csamul_cla12_and7_3(.a(a[7]), .b(b[3]), .out(s_csamul_cla12_and7_3));
  fa fa_s_csamul_cla12_fa7_3_out(.a(s_csamul_cla12_and7_3[0]), .b(s_csamul_cla12_fa8_2_xor1[0]), .cin(s_csamul_cla12_fa7_2_or0[0]), .fa_xor1(s_csamul_cla12_fa7_3_xor1), .fa_or0(s_csamul_cla12_fa7_3_or0));
  and_gate and_gate_s_csamul_cla12_and8_3(.a(a[8]), .b(b[3]), .out(s_csamul_cla12_and8_3));
  fa fa_s_csamul_cla12_fa8_3_out(.a(s_csamul_cla12_and8_3[0]), .b(s_csamul_cla12_fa9_2_xor1[0]), .cin(s_csamul_cla12_fa8_2_or0[0]), .fa_xor1(s_csamul_cla12_fa8_3_xor1), .fa_or0(s_csamul_cla12_fa8_3_or0));
  and_gate and_gate_s_csamul_cla12_and9_3(.a(a[9]), .b(b[3]), .out(s_csamul_cla12_and9_3));
  fa fa_s_csamul_cla12_fa9_3_out(.a(s_csamul_cla12_and9_3[0]), .b(s_csamul_cla12_fa10_2_xor1[0]), .cin(s_csamul_cla12_fa9_2_or0[0]), .fa_xor1(s_csamul_cla12_fa9_3_xor1), .fa_or0(s_csamul_cla12_fa9_3_or0));
  and_gate and_gate_s_csamul_cla12_and10_3(.a(a[10]), .b(b[3]), .out(s_csamul_cla12_and10_3));
  fa fa_s_csamul_cla12_fa10_3_out(.a(s_csamul_cla12_and10_3[0]), .b(s_csamul_cla12_ha11_2_xor0[0]), .cin(s_csamul_cla12_fa10_2_or0[0]), .fa_xor1(s_csamul_cla12_fa10_3_xor1), .fa_or0(s_csamul_cla12_fa10_3_or0));
  nand_gate nand_gate_s_csamul_cla12_nand11_3(.a(a[11]), .b(b[3]), .out(s_csamul_cla12_nand11_3));
  ha ha_s_csamul_cla12_ha11_3_out(.a(s_csamul_cla12_nand11_3[0]), .b(s_csamul_cla12_ha11_2_and0[0]), .ha_xor0(s_csamul_cla12_ha11_3_xor0), .ha_and0(s_csamul_cla12_ha11_3_and0));
  and_gate and_gate_s_csamul_cla12_and0_4(.a(a[0]), .b(b[4]), .out(s_csamul_cla12_and0_4));
  fa fa_s_csamul_cla12_fa0_4_out(.a(s_csamul_cla12_and0_4[0]), .b(s_csamul_cla12_fa1_3_xor1[0]), .cin(s_csamul_cla12_fa0_3_or0[0]), .fa_xor1(s_csamul_cla12_fa0_4_xor1), .fa_or0(s_csamul_cla12_fa0_4_or0));
  and_gate and_gate_s_csamul_cla12_and1_4(.a(a[1]), .b(b[4]), .out(s_csamul_cla12_and1_4));
  fa fa_s_csamul_cla12_fa1_4_out(.a(s_csamul_cla12_and1_4[0]), .b(s_csamul_cla12_fa2_3_xor1[0]), .cin(s_csamul_cla12_fa1_3_or0[0]), .fa_xor1(s_csamul_cla12_fa1_4_xor1), .fa_or0(s_csamul_cla12_fa1_4_or0));
  and_gate and_gate_s_csamul_cla12_and2_4(.a(a[2]), .b(b[4]), .out(s_csamul_cla12_and2_4));
  fa fa_s_csamul_cla12_fa2_4_out(.a(s_csamul_cla12_and2_4[0]), .b(s_csamul_cla12_fa3_3_xor1[0]), .cin(s_csamul_cla12_fa2_3_or0[0]), .fa_xor1(s_csamul_cla12_fa2_4_xor1), .fa_or0(s_csamul_cla12_fa2_4_or0));
  and_gate and_gate_s_csamul_cla12_and3_4(.a(a[3]), .b(b[4]), .out(s_csamul_cla12_and3_4));
  fa fa_s_csamul_cla12_fa3_4_out(.a(s_csamul_cla12_and3_4[0]), .b(s_csamul_cla12_fa4_3_xor1[0]), .cin(s_csamul_cla12_fa3_3_or0[0]), .fa_xor1(s_csamul_cla12_fa3_4_xor1), .fa_or0(s_csamul_cla12_fa3_4_or0));
  and_gate and_gate_s_csamul_cla12_and4_4(.a(a[4]), .b(b[4]), .out(s_csamul_cla12_and4_4));
  fa fa_s_csamul_cla12_fa4_4_out(.a(s_csamul_cla12_and4_4[0]), .b(s_csamul_cla12_fa5_3_xor1[0]), .cin(s_csamul_cla12_fa4_3_or0[0]), .fa_xor1(s_csamul_cla12_fa4_4_xor1), .fa_or0(s_csamul_cla12_fa4_4_or0));
  and_gate and_gate_s_csamul_cla12_and5_4(.a(a[5]), .b(b[4]), .out(s_csamul_cla12_and5_4));
  fa fa_s_csamul_cla12_fa5_4_out(.a(s_csamul_cla12_and5_4[0]), .b(s_csamul_cla12_fa6_3_xor1[0]), .cin(s_csamul_cla12_fa5_3_or0[0]), .fa_xor1(s_csamul_cla12_fa5_4_xor1), .fa_or0(s_csamul_cla12_fa5_4_or0));
  and_gate and_gate_s_csamul_cla12_and6_4(.a(a[6]), .b(b[4]), .out(s_csamul_cla12_and6_4));
  fa fa_s_csamul_cla12_fa6_4_out(.a(s_csamul_cla12_and6_4[0]), .b(s_csamul_cla12_fa7_3_xor1[0]), .cin(s_csamul_cla12_fa6_3_or0[0]), .fa_xor1(s_csamul_cla12_fa6_4_xor1), .fa_or0(s_csamul_cla12_fa6_4_or0));
  and_gate and_gate_s_csamul_cla12_and7_4(.a(a[7]), .b(b[4]), .out(s_csamul_cla12_and7_4));
  fa fa_s_csamul_cla12_fa7_4_out(.a(s_csamul_cla12_and7_4[0]), .b(s_csamul_cla12_fa8_3_xor1[0]), .cin(s_csamul_cla12_fa7_3_or0[0]), .fa_xor1(s_csamul_cla12_fa7_4_xor1), .fa_or0(s_csamul_cla12_fa7_4_or0));
  and_gate and_gate_s_csamul_cla12_and8_4(.a(a[8]), .b(b[4]), .out(s_csamul_cla12_and8_4));
  fa fa_s_csamul_cla12_fa8_4_out(.a(s_csamul_cla12_and8_4[0]), .b(s_csamul_cla12_fa9_3_xor1[0]), .cin(s_csamul_cla12_fa8_3_or0[0]), .fa_xor1(s_csamul_cla12_fa8_4_xor1), .fa_or0(s_csamul_cla12_fa8_4_or0));
  and_gate and_gate_s_csamul_cla12_and9_4(.a(a[9]), .b(b[4]), .out(s_csamul_cla12_and9_4));
  fa fa_s_csamul_cla12_fa9_4_out(.a(s_csamul_cla12_and9_4[0]), .b(s_csamul_cla12_fa10_3_xor1[0]), .cin(s_csamul_cla12_fa9_3_or0[0]), .fa_xor1(s_csamul_cla12_fa9_4_xor1), .fa_or0(s_csamul_cla12_fa9_4_or0));
  and_gate and_gate_s_csamul_cla12_and10_4(.a(a[10]), .b(b[4]), .out(s_csamul_cla12_and10_4));
  fa fa_s_csamul_cla12_fa10_4_out(.a(s_csamul_cla12_and10_4[0]), .b(s_csamul_cla12_ha11_3_xor0[0]), .cin(s_csamul_cla12_fa10_3_or0[0]), .fa_xor1(s_csamul_cla12_fa10_4_xor1), .fa_or0(s_csamul_cla12_fa10_4_or0));
  nand_gate nand_gate_s_csamul_cla12_nand11_4(.a(a[11]), .b(b[4]), .out(s_csamul_cla12_nand11_4));
  ha ha_s_csamul_cla12_ha11_4_out(.a(s_csamul_cla12_nand11_4[0]), .b(s_csamul_cla12_ha11_3_and0[0]), .ha_xor0(s_csamul_cla12_ha11_4_xor0), .ha_and0(s_csamul_cla12_ha11_4_and0));
  and_gate and_gate_s_csamul_cla12_and0_5(.a(a[0]), .b(b[5]), .out(s_csamul_cla12_and0_5));
  fa fa_s_csamul_cla12_fa0_5_out(.a(s_csamul_cla12_and0_5[0]), .b(s_csamul_cla12_fa1_4_xor1[0]), .cin(s_csamul_cla12_fa0_4_or0[0]), .fa_xor1(s_csamul_cla12_fa0_5_xor1), .fa_or0(s_csamul_cla12_fa0_5_or0));
  and_gate and_gate_s_csamul_cla12_and1_5(.a(a[1]), .b(b[5]), .out(s_csamul_cla12_and1_5));
  fa fa_s_csamul_cla12_fa1_5_out(.a(s_csamul_cla12_and1_5[0]), .b(s_csamul_cla12_fa2_4_xor1[0]), .cin(s_csamul_cla12_fa1_4_or0[0]), .fa_xor1(s_csamul_cla12_fa1_5_xor1), .fa_or0(s_csamul_cla12_fa1_5_or0));
  and_gate and_gate_s_csamul_cla12_and2_5(.a(a[2]), .b(b[5]), .out(s_csamul_cla12_and2_5));
  fa fa_s_csamul_cla12_fa2_5_out(.a(s_csamul_cla12_and2_5[0]), .b(s_csamul_cla12_fa3_4_xor1[0]), .cin(s_csamul_cla12_fa2_4_or0[0]), .fa_xor1(s_csamul_cla12_fa2_5_xor1), .fa_or0(s_csamul_cla12_fa2_5_or0));
  and_gate and_gate_s_csamul_cla12_and3_5(.a(a[3]), .b(b[5]), .out(s_csamul_cla12_and3_5));
  fa fa_s_csamul_cla12_fa3_5_out(.a(s_csamul_cla12_and3_5[0]), .b(s_csamul_cla12_fa4_4_xor1[0]), .cin(s_csamul_cla12_fa3_4_or0[0]), .fa_xor1(s_csamul_cla12_fa3_5_xor1), .fa_or0(s_csamul_cla12_fa3_5_or0));
  and_gate and_gate_s_csamul_cla12_and4_5(.a(a[4]), .b(b[5]), .out(s_csamul_cla12_and4_5));
  fa fa_s_csamul_cla12_fa4_5_out(.a(s_csamul_cla12_and4_5[0]), .b(s_csamul_cla12_fa5_4_xor1[0]), .cin(s_csamul_cla12_fa4_4_or0[0]), .fa_xor1(s_csamul_cla12_fa4_5_xor1), .fa_or0(s_csamul_cla12_fa4_5_or0));
  and_gate and_gate_s_csamul_cla12_and5_5(.a(a[5]), .b(b[5]), .out(s_csamul_cla12_and5_5));
  fa fa_s_csamul_cla12_fa5_5_out(.a(s_csamul_cla12_and5_5[0]), .b(s_csamul_cla12_fa6_4_xor1[0]), .cin(s_csamul_cla12_fa5_4_or0[0]), .fa_xor1(s_csamul_cla12_fa5_5_xor1), .fa_or0(s_csamul_cla12_fa5_5_or0));
  and_gate and_gate_s_csamul_cla12_and6_5(.a(a[6]), .b(b[5]), .out(s_csamul_cla12_and6_5));
  fa fa_s_csamul_cla12_fa6_5_out(.a(s_csamul_cla12_and6_5[0]), .b(s_csamul_cla12_fa7_4_xor1[0]), .cin(s_csamul_cla12_fa6_4_or0[0]), .fa_xor1(s_csamul_cla12_fa6_5_xor1), .fa_or0(s_csamul_cla12_fa6_5_or0));
  and_gate and_gate_s_csamul_cla12_and7_5(.a(a[7]), .b(b[5]), .out(s_csamul_cla12_and7_5));
  fa fa_s_csamul_cla12_fa7_5_out(.a(s_csamul_cla12_and7_5[0]), .b(s_csamul_cla12_fa8_4_xor1[0]), .cin(s_csamul_cla12_fa7_4_or0[0]), .fa_xor1(s_csamul_cla12_fa7_5_xor1), .fa_or0(s_csamul_cla12_fa7_5_or0));
  and_gate and_gate_s_csamul_cla12_and8_5(.a(a[8]), .b(b[5]), .out(s_csamul_cla12_and8_5));
  fa fa_s_csamul_cla12_fa8_5_out(.a(s_csamul_cla12_and8_5[0]), .b(s_csamul_cla12_fa9_4_xor1[0]), .cin(s_csamul_cla12_fa8_4_or0[0]), .fa_xor1(s_csamul_cla12_fa8_5_xor1), .fa_or0(s_csamul_cla12_fa8_5_or0));
  and_gate and_gate_s_csamul_cla12_and9_5(.a(a[9]), .b(b[5]), .out(s_csamul_cla12_and9_5));
  fa fa_s_csamul_cla12_fa9_5_out(.a(s_csamul_cla12_and9_5[0]), .b(s_csamul_cla12_fa10_4_xor1[0]), .cin(s_csamul_cla12_fa9_4_or0[0]), .fa_xor1(s_csamul_cla12_fa9_5_xor1), .fa_or0(s_csamul_cla12_fa9_5_or0));
  and_gate and_gate_s_csamul_cla12_and10_5(.a(a[10]), .b(b[5]), .out(s_csamul_cla12_and10_5));
  fa fa_s_csamul_cla12_fa10_5_out(.a(s_csamul_cla12_and10_5[0]), .b(s_csamul_cla12_ha11_4_xor0[0]), .cin(s_csamul_cla12_fa10_4_or0[0]), .fa_xor1(s_csamul_cla12_fa10_5_xor1), .fa_or0(s_csamul_cla12_fa10_5_or0));
  nand_gate nand_gate_s_csamul_cla12_nand11_5(.a(a[11]), .b(b[5]), .out(s_csamul_cla12_nand11_5));
  ha ha_s_csamul_cla12_ha11_5_out(.a(s_csamul_cla12_nand11_5[0]), .b(s_csamul_cla12_ha11_4_and0[0]), .ha_xor0(s_csamul_cla12_ha11_5_xor0), .ha_and0(s_csamul_cla12_ha11_5_and0));
  and_gate and_gate_s_csamul_cla12_and0_6(.a(a[0]), .b(b[6]), .out(s_csamul_cla12_and0_6));
  fa fa_s_csamul_cla12_fa0_6_out(.a(s_csamul_cla12_and0_6[0]), .b(s_csamul_cla12_fa1_5_xor1[0]), .cin(s_csamul_cla12_fa0_5_or0[0]), .fa_xor1(s_csamul_cla12_fa0_6_xor1), .fa_or0(s_csamul_cla12_fa0_6_or0));
  and_gate and_gate_s_csamul_cla12_and1_6(.a(a[1]), .b(b[6]), .out(s_csamul_cla12_and1_6));
  fa fa_s_csamul_cla12_fa1_6_out(.a(s_csamul_cla12_and1_6[0]), .b(s_csamul_cla12_fa2_5_xor1[0]), .cin(s_csamul_cla12_fa1_5_or0[0]), .fa_xor1(s_csamul_cla12_fa1_6_xor1), .fa_or0(s_csamul_cla12_fa1_6_or0));
  and_gate and_gate_s_csamul_cla12_and2_6(.a(a[2]), .b(b[6]), .out(s_csamul_cla12_and2_6));
  fa fa_s_csamul_cla12_fa2_6_out(.a(s_csamul_cla12_and2_6[0]), .b(s_csamul_cla12_fa3_5_xor1[0]), .cin(s_csamul_cla12_fa2_5_or0[0]), .fa_xor1(s_csamul_cla12_fa2_6_xor1), .fa_or0(s_csamul_cla12_fa2_6_or0));
  and_gate and_gate_s_csamul_cla12_and3_6(.a(a[3]), .b(b[6]), .out(s_csamul_cla12_and3_6));
  fa fa_s_csamul_cla12_fa3_6_out(.a(s_csamul_cla12_and3_6[0]), .b(s_csamul_cla12_fa4_5_xor1[0]), .cin(s_csamul_cla12_fa3_5_or0[0]), .fa_xor1(s_csamul_cla12_fa3_6_xor1), .fa_or0(s_csamul_cla12_fa3_6_or0));
  and_gate and_gate_s_csamul_cla12_and4_6(.a(a[4]), .b(b[6]), .out(s_csamul_cla12_and4_6));
  fa fa_s_csamul_cla12_fa4_6_out(.a(s_csamul_cla12_and4_6[0]), .b(s_csamul_cla12_fa5_5_xor1[0]), .cin(s_csamul_cla12_fa4_5_or0[0]), .fa_xor1(s_csamul_cla12_fa4_6_xor1), .fa_or0(s_csamul_cla12_fa4_6_or0));
  and_gate and_gate_s_csamul_cla12_and5_6(.a(a[5]), .b(b[6]), .out(s_csamul_cla12_and5_6));
  fa fa_s_csamul_cla12_fa5_6_out(.a(s_csamul_cla12_and5_6[0]), .b(s_csamul_cla12_fa6_5_xor1[0]), .cin(s_csamul_cla12_fa5_5_or0[0]), .fa_xor1(s_csamul_cla12_fa5_6_xor1), .fa_or0(s_csamul_cla12_fa5_6_or0));
  and_gate and_gate_s_csamul_cla12_and6_6(.a(a[6]), .b(b[6]), .out(s_csamul_cla12_and6_6));
  fa fa_s_csamul_cla12_fa6_6_out(.a(s_csamul_cla12_and6_6[0]), .b(s_csamul_cla12_fa7_5_xor1[0]), .cin(s_csamul_cla12_fa6_5_or0[0]), .fa_xor1(s_csamul_cla12_fa6_6_xor1), .fa_or0(s_csamul_cla12_fa6_6_or0));
  and_gate and_gate_s_csamul_cla12_and7_6(.a(a[7]), .b(b[6]), .out(s_csamul_cla12_and7_6));
  fa fa_s_csamul_cla12_fa7_6_out(.a(s_csamul_cla12_and7_6[0]), .b(s_csamul_cla12_fa8_5_xor1[0]), .cin(s_csamul_cla12_fa7_5_or0[0]), .fa_xor1(s_csamul_cla12_fa7_6_xor1), .fa_or0(s_csamul_cla12_fa7_6_or0));
  and_gate and_gate_s_csamul_cla12_and8_6(.a(a[8]), .b(b[6]), .out(s_csamul_cla12_and8_6));
  fa fa_s_csamul_cla12_fa8_6_out(.a(s_csamul_cla12_and8_6[0]), .b(s_csamul_cla12_fa9_5_xor1[0]), .cin(s_csamul_cla12_fa8_5_or0[0]), .fa_xor1(s_csamul_cla12_fa8_6_xor1), .fa_or0(s_csamul_cla12_fa8_6_or0));
  and_gate and_gate_s_csamul_cla12_and9_6(.a(a[9]), .b(b[6]), .out(s_csamul_cla12_and9_6));
  fa fa_s_csamul_cla12_fa9_6_out(.a(s_csamul_cla12_and9_6[0]), .b(s_csamul_cla12_fa10_5_xor1[0]), .cin(s_csamul_cla12_fa9_5_or0[0]), .fa_xor1(s_csamul_cla12_fa9_6_xor1), .fa_or0(s_csamul_cla12_fa9_6_or0));
  and_gate and_gate_s_csamul_cla12_and10_6(.a(a[10]), .b(b[6]), .out(s_csamul_cla12_and10_6));
  fa fa_s_csamul_cla12_fa10_6_out(.a(s_csamul_cla12_and10_6[0]), .b(s_csamul_cla12_ha11_5_xor0[0]), .cin(s_csamul_cla12_fa10_5_or0[0]), .fa_xor1(s_csamul_cla12_fa10_6_xor1), .fa_or0(s_csamul_cla12_fa10_6_or0));
  nand_gate nand_gate_s_csamul_cla12_nand11_6(.a(a[11]), .b(b[6]), .out(s_csamul_cla12_nand11_6));
  ha ha_s_csamul_cla12_ha11_6_out(.a(s_csamul_cla12_nand11_6[0]), .b(s_csamul_cla12_ha11_5_and0[0]), .ha_xor0(s_csamul_cla12_ha11_6_xor0), .ha_and0(s_csamul_cla12_ha11_6_and0));
  and_gate and_gate_s_csamul_cla12_and0_7(.a(a[0]), .b(b[7]), .out(s_csamul_cla12_and0_7));
  fa fa_s_csamul_cla12_fa0_7_out(.a(s_csamul_cla12_and0_7[0]), .b(s_csamul_cla12_fa1_6_xor1[0]), .cin(s_csamul_cla12_fa0_6_or0[0]), .fa_xor1(s_csamul_cla12_fa0_7_xor1), .fa_or0(s_csamul_cla12_fa0_7_or0));
  and_gate and_gate_s_csamul_cla12_and1_7(.a(a[1]), .b(b[7]), .out(s_csamul_cla12_and1_7));
  fa fa_s_csamul_cla12_fa1_7_out(.a(s_csamul_cla12_and1_7[0]), .b(s_csamul_cla12_fa2_6_xor1[0]), .cin(s_csamul_cla12_fa1_6_or0[0]), .fa_xor1(s_csamul_cla12_fa1_7_xor1), .fa_or0(s_csamul_cla12_fa1_7_or0));
  and_gate and_gate_s_csamul_cla12_and2_7(.a(a[2]), .b(b[7]), .out(s_csamul_cla12_and2_7));
  fa fa_s_csamul_cla12_fa2_7_out(.a(s_csamul_cla12_and2_7[0]), .b(s_csamul_cla12_fa3_6_xor1[0]), .cin(s_csamul_cla12_fa2_6_or0[0]), .fa_xor1(s_csamul_cla12_fa2_7_xor1), .fa_or0(s_csamul_cla12_fa2_7_or0));
  and_gate and_gate_s_csamul_cla12_and3_7(.a(a[3]), .b(b[7]), .out(s_csamul_cla12_and3_7));
  fa fa_s_csamul_cla12_fa3_7_out(.a(s_csamul_cla12_and3_7[0]), .b(s_csamul_cla12_fa4_6_xor1[0]), .cin(s_csamul_cla12_fa3_6_or0[0]), .fa_xor1(s_csamul_cla12_fa3_7_xor1), .fa_or0(s_csamul_cla12_fa3_7_or0));
  and_gate and_gate_s_csamul_cla12_and4_7(.a(a[4]), .b(b[7]), .out(s_csamul_cla12_and4_7));
  fa fa_s_csamul_cla12_fa4_7_out(.a(s_csamul_cla12_and4_7[0]), .b(s_csamul_cla12_fa5_6_xor1[0]), .cin(s_csamul_cla12_fa4_6_or0[0]), .fa_xor1(s_csamul_cla12_fa4_7_xor1), .fa_or0(s_csamul_cla12_fa4_7_or0));
  and_gate and_gate_s_csamul_cla12_and5_7(.a(a[5]), .b(b[7]), .out(s_csamul_cla12_and5_7));
  fa fa_s_csamul_cla12_fa5_7_out(.a(s_csamul_cla12_and5_7[0]), .b(s_csamul_cla12_fa6_6_xor1[0]), .cin(s_csamul_cla12_fa5_6_or0[0]), .fa_xor1(s_csamul_cla12_fa5_7_xor1), .fa_or0(s_csamul_cla12_fa5_7_or0));
  and_gate and_gate_s_csamul_cla12_and6_7(.a(a[6]), .b(b[7]), .out(s_csamul_cla12_and6_7));
  fa fa_s_csamul_cla12_fa6_7_out(.a(s_csamul_cla12_and6_7[0]), .b(s_csamul_cla12_fa7_6_xor1[0]), .cin(s_csamul_cla12_fa6_6_or0[0]), .fa_xor1(s_csamul_cla12_fa6_7_xor1), .fa_or0(s_csamul_cla12_fa6_7_or0));
  and_gate and_gate_s_csamul_cla12_and7_7(.a(a[7]), .b(b[7]), .out(s_csamul_cla12_and7_7));
  fa fa_s_csamul_cla12_fa7_7_out(.a(s_csamul_cla12_and7_7[0]), .b(s_csamul_cla12_fa8_6_xor1[0]), .cin(s_csamul_cla12_fa7_6_or0[0]), .fa_xor1(s_csamul_cla12_fa7_7_xor1), .fa_or0(s_csamul_cla12_fa7_7_or0));
  and_gate and_gate_s_csamul_cla12_and8_7(.a(a[8]), .b(b[7]), .out(s_csamul_cla12_and8_7));
  fa fa_s_csamul_cla12_fa8_7_out(.a(s_csamul_cla12_and8_7[0]), .b(s_csamul_cla12_fa9_6_xor1[0]), .cin(s_csamul_cla12_fa8_6_or0[0]), .fa_xor1(s_csamul_cla12_fa8_7_xor1), .fa_or0(s_csamul_cla12_fa8_7_or0));
  and_gate and_gate_s_csamul_cla12_and9_7(.a(a[9]), .b(b[7]), .out(s_csamul_cla12_and9_7));
  fa fa_s_csamul_cla12_fa9_7_out(.a(s_csamul_cla12_and9_7[0]), .b(s_csamul_cla12_fa10_6_xor1[0]), .cin(s_csamul_cla12_fa9_6_or0[0]), .fa_xor1(s_csamul_cla12_fa9_7_xor1), .fa_or0(s_csamul_cla12_fa9_7_or0));
  and_gate and_gate_s_csamul_cla12_and10_7(.a(a[10]), .b(b[7]), .out(s_csamul_cla12_and10_7));
  fa fa_s_csamul_cla12_fa10_7_out(.a(s_csamul_cla12_and10_7[0]), .b(s_csamul_cla12_ha11_6_xor0[0]), .cin(s_csamul_cla12_fa10_6_or0[0]), .fa_xor1(s_csamul_cla12_fa10_7_xor1), .fa_or0(s_csamul_cla12_fa10_7_or0));
  nand_gate nand_gate_s_csamul_cla12_nand11_7(.a(a[11]), .b(b[7]), .out(s_csamul_cla12_nand11_7));
  ha ha_s_csamul_cla12_ha11_7_out(.a(s_csamul_cla12_nand11_7[0]), .b(s_csamul_cla12_ha11_6_and0[0]), .ha_xor0(s_csamul_cla12_ha11_7_xor0), .ha_and0(s_csamul_cla12_ha11_7_and0));
  and_gate and_gate_s_csamul_cla12_and0_8(.a(a[0]), .b(b[8]), .out(s_csamul_cla12_and0_8));
  fa fa_s_csamul_cla12_fa0_8_out(.a(s_csamul_cla12_and0_8[0]), .b(s_csamul_cla12_fa1_7_xor1[0]), .cin(s_csamul_cla12_fa0_7_or0[0]), .fa_xor1(s_csamul_cla12_fa0_8_xor1), .fa_or0(s_csamul_cla12_fa0_8_or0));
  and_gate and_gate_s_csamul_cla12_and1_8(.a(a[1]), .b(b[8]), .out(s_csamul_cla12_and1_8));
  fa fa_s_csamul_cla12_fa1_8_out(.a(s_csamul_cla12_and1_8[0]), .b(s_csamul_cla12_fa2_7_xor1[0]), .cin(s_csamul_cla12_fa1_7_or0[0]), .fa_xor1(s_csamul_cla12_fa1_8_xor1), .fa_or0(s_csamul_cla12_fa1_8_or0));
  and_gate and_gate_s_csamul_cla12_and2_8(.a(a[2]), .b(b[8]), .out(s_csamul_cla12_and2_8));
  fa fa_s_csamul_cla12_fa2_8_out(.a(s_csamul_cla12_and2_8[0]), .b(s_csamul_cla12_fa3_7_xor1[0]), .cin(s_csamul_cla12_fa2_7_or0[0]), .fa_xor1(s_csamul_cla12_fa2_8_xor1), .fa_or0(s_csamul_cla12_fa2_8_or0));
  and_gate and_gate_s_csamul_cla12_and3_8(.a(a[3]), .b(b[8]), .out(s_csamul_cla12_and3_8));
  fa fa_s_csamul_cla12_fa3_8_out(.a(s_csamul_cla12_and3_8[0]), .b(s_csamul_cla12_fa4_7_xor1[0]), .cin(s_csamul_cla12_fa3_7_or0[0]), .fa_xor1(s_csamul_cla12_fa3_8_xor1), .fa_or0(s_csamul_cla12_fa3_8_or0));
  and_gate and_gate_s_csamul_cla12_and4_8(.a(a[4]), .b(b[8]), .out(s_csamul_cla12_and4_8));
  fa fa_s_csamul_cla12_fa4_8_out(.a(s_csamul_cla12_and4_8[0]), .b(s_csamul_cla12_fa5_7_xor1[0]), .cin(s_csamul_cla12_fa4_7_or0[0]), .fa_xor1(s_csamul_cla12_fa4_8_xor1), .fa_or0(s_csamul_cla12_fa4_8_or0));
  and_gate and_gate_s_csamul_cla12_and5_8(.a(a[5]), .b(b[8]), .out(s_csamul_cla12_and5_8));
  fa fa_s_csamul_cla12_fa5_8_out(.a(s_csamul_cla12_and5_8[0]), .b(s_csamul_cla12_fa6_7_xor1[0]), .cin(s_csamul_cla12_fa5_7_or0[0]), .fa_xor1(s_csamul_cla12_fa5_8_xor1), .fa_or0(s_csamul_cla12_fa5_8_or0));
  and_gate and_gate_s_csamul_cla12_and6_8(.a(a[6]), .b(b[8]), .out(s_csamul_cla12_and6_8));
  fa fa_s_csamul_cla12_fa6_8_out(.a(s_csamul_cla12_and6_8[0]), .b(s_csamul_cla12_fa7_7_xor1[0]), .cin(s_csamul_cla12_fa6_7_or0[0]), .fa_xor1(s_csamul_cla12_fa6_8_xor1), .fa_or0(s_csamul_cla12_fa6_8_or0));
  and_gate and_gate_s_csamul_cla12_and7_8(.a(a[7]), .b(b[8]), .out(s_csamul_cla12_and7_8));
  fa fa_s_csamul_cla12_fa7_8_out(.a(s_csamul_cla12_and7_8[0]), .b(s_csamul_cla12_fa8_7_xor1[0]), .cin(s_csamul_cla12_fa7_7_or0[0]), .fa_xor1(s_csamul_cla12_fa7_8_xor1), .fa_or0(s_csamul_cla12_fa7_8_or0));
  and_gate and_gate_s_csamul_cla12_and8_8(.a(a[8]), .b(b[8]), .out(s_csamul_cla12_and8_8));
  fa fa_s_csamul_cla12_fa8_8_out(.a(s_csamul_cla12_and8_8[0]), .b(s_csamul_cla12_fa9_7_xor1[0]), .cin(s_csamul_cla12_fa8_7_or0[0]), .fa_xor1(s_csamul_cla12_fa8_8_xor1), .fa_or0(s_csamul_cla12_fa8_8_or0));
  and_gate and_gate_s_csamul_cla12_and9_8(.a(a[9]), .b(b[8]), .out(s_csamul_cla12_and9_8));
  fa fa_s_csamul_cla12_fa9_8_out(.a(s_csamul_cla12_and9_8[0]), .b(s_csamul_cla12_fa10_7_xor1[0]), .cin(s_csamul_cla12_fa9_7_or0[0]), .fa_xor1(s_csamul_cla12_fa9_8_xor1), .fa_or0(s_csamul_cla12_fa9_8_or0));
  and_gate and_gate_s_csamul_cla12_and10_8(.a(a[10]), .b(b[8]), .out(s_csamul_cla12_and10_8));
  fa fa_s_csamul_cla12_fa10_8_out(.a(s_csamul_cla12_and10_8[0]), .b(s_csamul_cla12_ha11_7_xor0[0]), .cin(s_csamul_cla12_fa10_7_or0[0]), .fa_xor1(s_csamul_cla12_fa10_8_xor1), .fa_or0(s_csamul_cla12_fa10_8_or0));
  nand_gate nand_gate_s_csamul_cla12_nand11_8(.a(a[11]), .b(b[8]), .out(s_csamul_cla12_nand11_8));
  ha ha_s_csamul_cla12_ha11_8_out(.a(s_csamul_cla12_nand11_8[0]), .b(s_csamul_cla12_ha11_7_and0[0]), .ha_xor0(s_csamul_cla12_ha11_8_xor0), .ha_and0(s_csamul_cla12_ha11_8_and0));
  and_gate and_gate_s_csamul_cla12_and0_9(.a(a[0]), .b(b[9]), .out(s_csamul_cla12_and0_9));
  fa fa_s_csamul_cla12_fa0_9_out(.a(s_csamul_cla12_and0_9[0]), .b(s_csamul_cla12_fa1_8_xor1[0]), .cin(s_csamul_cla12_fa0_8_or0[0]), .fa_xor1(s_csamul_cla12_fa0_9_xor1), .fa_or0(s_csamul_cla12_fa0_9_or0));
  and_gate and_gate_s_csamul_cla12_and1_9(.a(a[1]), .b(b[9]), .out(s_csamul_cla12_and1_9));
  fa fa_s_csamul_cla12_fa1_9_out(.a(s_csamul_cla12_and1_9[0]), .b(s_csamul_cla12_fa2_8_xor1[0]), .cin(s_csamul_cla12_fa1_8_or0[0]), .fa_xor1(s_csamul_cla12_fa1_9_xor1), .fa_or0(s_csamul_cla12_fa1_9_or0));
  and_gate and_gate_s_csamul_cla12_and2_9(.a(a[2]), .b(b[9]), .out(s_csamul_cla12_and2_9));
  fa fa_s_csamul_cla12_fa2_9_out(.a(s_csamul_cla12_and2_9[0]), .b(s_csamul_cla12_fa3_8_xor1[0]), .cin(s_csamul_cla12_fa2_8_or0[0]), .fa_xor1(s_csamul_cla12_fa2_9_xor1), .fa_or0(s_csamul_cla12_fa2_9_or0));
  and_gate and_gate_s_csamul_cla12_and3_9(.a(a[3]), .b(b[9]), .out(s_csamul_cla12_and3_9));
  fa fa_s_csamul_cla12_fa3_9_out(.a(s_csamul_cla12_and3_9[0]), .b(s_csamul_cla12_fa4_8_xor1[0]), .cin(s_csamul_cla12_fa3_8_or0[0]), .fa_xor1(s_csamul_cla12_fa3_9_xor1), .fa_or0(s_csamul_cla12_fa3_9_or0));
  and_gate and_gate_s_csamul_cla12_and4_9(.a(a[4]), .b(b[9]), .out(s_csamul_cla12_and4_9));
  fa fa_s_csamul_cla12_fa4_9_out(.a(s_csamul_cla12_and4_9[0]), .b(s_csamul_cla12_fa5_8_xor1[0]), .cin(s_csamul_cla12_fa4_8_or0[0]), .fa_xor1(s_csamul_cla12_fa4_9_xor1), .fa_or0(s_csamul_cla12_fa4_9_or0));
  and_gate and_gate_s_csamul_cla12_and5_9(.a(a[5]), .b(b[9]), .out(s_csamul_cla12_and5_9));
  fa fa_s_csamul_cla12_fa5_9_out(.a(s_csamul_cla12_and5_9[0]), .b(s_csamul_cla12_fa6_8_xor1[0]), .cin(s_csamul_cla12_fa5_8_or0[0]), .fa_xor1(s_csamul_cla12_fa5_9_xor1), .fa_or0(s_csamul_cla12_fa5_9_or0));
  and_gate and_gate_s_csamul_cla12_and6_9(.a(a[6]), .b(b[9]), .out(s_csamul_cla12_and6_9));
  fa fa_s_csamul_cla12_fa6_9_out(.a(s_csamul_cla12_and6_9[0]), .b(s_csamul_cla12_fa7_8_xor1[0]), .cin(s_csamul_cla12_fa6_8_or0[0]), .fa_xor1(s_csamul_cla12_fa6_9_xor1), .fa_or0(s_csamul_cla12_fa6_9_or0));
  and_gate and_gate_s_csamul_cla12_and7_9(.a(a[7]), .b(b[9]), .out(s_csamul_cla12_and7_9));
  fa fa_s_csamul_cla12_fa7_9_out(.a(s_csamul_cla12_and7_9[0]), .b(s_csamul_cla12_fa8_8_xor1[0]), .cin(s_csamul_cla12_fa7_8_or0[0]), .fa_xor1(s_csamul_cla12_fa7_9_xor1), .fa_or0(s_csamul_cla12_fa7_9_or0));
  and_gate and_gate_s_csamul_cla12_and8_9(.a(a[8]), .b(b[9]), .out(s_csamul_cla12_and8_9));
  fa fa_s_csamul_cla12_fa8_9_out(.a(s_csamul_cla12_and8_9[0]), .b(s_csamul_cla12_fa9_8_xor1[0]), .cin(s_csamul_cla12_fa8_8_or0[0]), .fa_xor1(s_csamul_cla12_fa8_9_xor1), .fa_or0(s_csamul_cla12_fa8_9_or0));
  and_gate and_gate_s_csamul_cla12_and9_9(.a(a[9]), .b(b[9]), .out(s_csamul_cla12_and9_9));
  fa fa_s_csamul_cla12_fa9_9_out(.a(s_csamul_cla12_and9_9[0]), .b(s_csamul_cla12_fa10_8_xor1[0]), .cin(s_csamul_cla12_fa9_8_or0[0]), .fa_xor1(s_csamul_cla12_fa9_9_xor1), .fa_or0(s_csamul_cla12_fa9_9_or0));
  and_gate and_gate_s_csamul_cla12_and10_9(.a(a[10]), .b(b[9]), .out(s_csamul_cla12_and10_9));
  fa fa_s_csamul_cla12_fa10_9_out(.a(s_csamul_cla12_and10_9[0]), .b(s_csamul_cla12_ha11_8_xor0[0]), .cin(s_csamul_cla12_fa10_8_or0[0]), .fa_xor1(s_csamul_cla12_fa10_9_xor1), .fa_or0(s_csamul_cla12_fa10_9_or0));
  nand_gate nand_gate_s_csamul_cla12_nand11_9(.a(a[11]), .b(b[9]), .out(s_csamul_cla12_nand11_9));
  ha ha_s_csamul_cla12_ha11_9_out(.a(s_csamul_cla12_nand11_9[0]), .b(s_csamul_cla12_ha11_8_and0[0]), .ha_xor0(s_csamul_cla12_ha11_9_xor0), .ha_and0(s_csamul_cla12_ha11_9_and0));
  and_gate and_gate_s_csamul_cla12_and0_10(.a(a[0]), .b(b[10]), .out(s_csamul_cla12_and0_10));
  fa fa_s_csamul_cla12_fa0_10_out(.a(s_csamul_cla12_and0_10[0]), .b(s_csamul_cla12_fa1_9_xor1[0]), .cin(s_csamul_cla12_fa0_9_or0[0]), .fa_xor1(s_csamul_cla12_fa0_10_xor1), .fa_or0(s_csamul_cla12_fa0_10_or0));
  and_gate and_gate_s_csamul_cla12_and1_10(.a(a[1]), .b(b[10]), .out(s_csamul_cla12_and1_10));
  fa fa_s_csamul_cla12_fa1_10_out(.a(s_csamul_cla12_and1_10[0]), .b(s_csamul_cla12_fa2_9_xor1[0]), .cin(s_csamul_cla12_fa1_9_or0[0]), .fa_xor1(s_csamul_cla12_fa1_10_xor1), .fa_or0(s_csamul_cla12_fa1_10_or0));
  and_gate and_gate_s_csamul_cla12_and2_10(.a(a[2]), .b(b[10]), .out(s_csamul_cla12_and2_10));
  fa fa_s_csamul_cla12_fa2_10_out(.a(s_csamul_cla12_and2_10[0]), .b(s_csamul_cla12_fa3_9_xor1[0]), .cin(s_csamul_cla12_fa2_9_or0[0]), .fa_xor1(s_csamul_cla12_fa2_10_xor1), .fa_or0(s_csamul_cla12_fa2_10_or0));
  and_gate and_gate_s_csamul_cla12_and3_10(.a(a[3]), .b(b[10]), .out(s_csamul_cla12_and3_10));
  fa fa_s_csamul_cla12_fa3_10_out(.a(s_csamul_cla12_and3_10[0]), .b(s_csamul_cla12_fa4_9_xor1[0]), .cin(s_csamul_cla12_fa3_9_or0[0]), .fa_xor1(s_csamul_cla12_fa3_10_xor1), .fa_or0(s_csamul_cla12_fa3_10_or0));
  and_gate and_gate_s_csamul_cla12_and4_10(.a(a[4]), .b(b[10]), .out(s_csamul_cla12_and4_10));
  fa fa_s_csamul_cla12_fa4_10_out(.a(s_csamul_cla12_and4_10[0]), .b(s_csamul_cla12_fa5_9_xor1[0]), .cin(s_csamul_cla12_fa4_9_or0[0]), .fa_xor1(s_csamul_cla12_fa4_10_xor1), .fa_or0(s_csamul_cla12_fa4_10_or0));
  and_gate and_gate_s_csamul_cla12_and5_10(.a(a[5]), .b(b[10]), .out(s_csamul_cla12_and5_10));
  fa fa_s_csamul_cla12_fa5_10_out(.a(s_csamul_cla12_and5_10[0]), .b(s_csamul_cla12_fa6_9_xor1[0]), .cin(s_csamul_cla12_fa5_9_or0[0]), .fa_xor1(s_csamul_cla12_fa5_10_xor1), .fa_or0(s_csamul_cla12_fa5_10_or0));
  and_gate and_gate_s_csamul_cla12_and6_10(.a(a[6]), .b(b[10]), .out(s_csamul_cla12_and6_10));
  fa fa_s_csamul_cla12_fa6_10_out(.a(s_csamul_cla12_and6_10[0]), .b(s_csamul_cla12_fa7_9_xor1[0]), .cin(s_csamul_cla12_fa6_9_or0[0]), .fa_xor1(s_csamul_cla12_fa6_10_xor1), .fa_or0(s_csamul_cla12_fa6_10_or0));
  and_gate and_gate_s_csamul_cla12_and7_10(.a(a[7]), .b(b[10]), .out(s_csamul_cla12_and7_10));
  fa fa_s_csamul_cla12_fa7_10_out(.a(s_csamul_cla12_and7_10[0]), .b(s_csamul_cla12_fa8_9_xor1[0]), .cin(s_csamul_cla12_fa7_9_or0[0]), .fa_xor1(s_csamul_cla12_fa7_10_xor1), .fa_or0(s_csamul_cla12_fa7_10_or0));
  and_gate and_gate_s_csamul_cla12_and8_10(.a(a[8]), .b(b[10]), .out(s_csamul_cla12_and8_10));
  fa fa_s_csamul_cla12_fa8_10_out(.a(s_csamul_cla12_and8_10[0]), .b(s_csamul_cla12_fa9_9_xor1[0]), .cin(s_csamul_cla12_fa8_9_or0[0]), .fa_xor1(s_csamul_cla12_fa8_10_xor1), .fa_or0(s_csamul_cla12_fa8_10_or0));
  and_gate and_gate_s_csamul_cla12_and9_10(.a(a[9]), .b(b[10]), .out(s_csamul_cla12_and9_10));
  fa fa_s_csamul_cla12_fa9_10_out(.a(s_csamul_cla12_and9_10[0]), .b(s_csamul_cla12_fa10_9_xor1[0]), .cin(s_csamul_cla12_fa9_9_or0[0]), .fa_xor1(s_csamul_cla12_fa9_10_xor1), .fa_or0(s_csamul_cla12_fa9_10_or0));
  and_gate and_gate_s_csamul_cla12_and10_10(.a(a[10]), .b(b[10]), .out(s_csamul_cla12_and10_10));
  fa fa_s_csamul_cla12_fa10_10_out(.a(s_csamul_cla12_and10_10[0]), .b(s_csamul_cla12_ha11_9_xor0[0]), .cin(s_csamul_cla12_fa10_9_or0[0]), .fa_xor1(s_csamul_cla12_fa10_10_xor1), .fa_or0(s_csamul_cla12_fa10_10_or0));
  nand_gate nand_gate_s_csamul_cla12_nand11_10(.a(a[11]), .b(b[10]), .out(s_csamul_cla12_nand11_10));
  ha ha_s_csamul_cla12_ha11_10_out(.a(s_csamul_cla12_nand11_10[0]), .b(s_csamul_cla12_ha11_9_and0[0]), .ha_xor0(s_csamul_cla12_ha11_10_xor0), .ha_and0(s_csamul_cla12_ha11_10_and0));
  nand_gate nand_gate_s_csamul_cla12_nand0_11(.a(a[0]), .b(b[11]), .out(s_csamul_cla12_nand0_11));
  fa fa_s_csamul_cla12_fa0_11_out(.a(s_csamul_cla12_nand0_11[0]), .b(s_csamul_cla12_fa1_10_xor1[0]), .cin(s_csamul_cla12_fa0_10_or0[0]), .fa_xor1(s_csamul_cla12_fa0_11_xor1), .fa_or0(s_csamul_cla12_fa0_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand1_11(.a(a[1]), .b(b[11]), .out(s_csamul_cla12_nand1_11));
  fa fa_s_csamul_cla12_fa1_11_out(.a(s_csamul_cla12_nand1_11[0]), .b(s_csamul_cla12_fa2_10_xor1[0]), .cin(s_csamul_cla12_fa1_10_or0[0]), .fa_xor1(s_csamul_cla12_fa1_11_xor1), .fa_or0(s_csamul_cla12_fa1_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand2_11(.a(a[2]), .b(b[11]), .out(s_csamul_cla12_nand2_11));
  fa fa_s_csamul_cla12_fa2_11_out(.a(s_csamul_cla12_nand2_11[0]), .b(s_csamul_cla12_fa3_10_xor1[0]), .cin(s_csamul_cla12_fa2_10_or0[0]), .fa_xor1(s_csamul_cla12_fa2_11_xor1), .fa_or0(s_csamul_cla12_fa2_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand3_11(.a(a[3]), .b(b[11]), .out(s_csamul_cla12_nand3_11));
  fa fa_s_csamul_cla12_fa3_11_out(.a(s_csamul_cla12_nand3_11[0]), .b(s_csamul_cla12_fa4_10_xor1[0]), .cin(s_csamul_cla12_fa3_10_or0[0]), .fa_xor1(s_csamul_cla12_fa3_11_xor1), .fa_or0(s_csamul_cla12_fa3_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand4_11(.a(a[4]), .b(b[11]), .out(s_csamul_cla12_nand4_11));
  fa fa_s_csamul_cla12_fa4_11_out(.a(s_csamul_cla12_nand4_11[0]), .b(s_csamul_cla12_fa5_10_xor1[0]), .cin(s_csamul_cla12_fa4_10_or0[0]), .fa_xor1(s_csamul_cla12_fa4_11_xor1), .fa_or0(s_csamul_cla12_fa4_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand5_11(.a(a[5]), .b(b[11]), .out(s_csamul_cla12_nand5_11));
  fa fa_s_csamul_cla12_fa5_11_out(.a(s_csamul_cla12_nand5_11[0]), .b(s_csamul_cla12_fa6_10_xor1[0]), .cin(s_csamul_cla12_fa5_10_or0[0]), .fa_xor1(s_csamul_cla12_fa5_11_xor1), .fa_or0(s_csamul_cla12_fa5_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand6_11(.a(a[6]), .b(b[11]), .out(s_csamul_cla12_nand6_11));
  fa fa_s_csamul_cla12_fa6_11_out(.a(s_csamul_cla12_nand6_11[0]), .b(s_csamul_cla12_fa7_10_xor1[0]), .cin(s_csamul_cla12_fa6_10_or0[0]), .fa_xor1(s_csamul_cla12_fa6_11_xor1), .fa_or0(s_csamul_cla12_fa6_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand7_11(.a(a[7]), .b(b[11]), .out(s_csamul_cla12_nand7_11));
  fa fa_s_csamul_cla12_fa7_11_out(.a(s_csamul_cla12_nand7_11[0]), .b(s_csamul_cla12_fa8_10_xor1[0]), .cin(s_csamul_cla12_fa7_10_or0[0]), .fa_xor1(s_csamul_cla12_fa7_11_xor1), .fa_or0(s_csamul_cla12_fa7_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand8_11(.a(a[8]), .b(b[11]), .out(s_csamul_cla12_nand8_11));
  fa fa_s_csamul_cla12_fa8_11_out(.a(s_csamul_cla12_nand8_11[0]), .b(s_csamul_cla12_fa9_10_xor1[0]), .cin(s_csamul_cla12_fa8_10_or0[0]), .fa_xor1(s_csamul_cla12_fa8_11_xor1), .fa_or0(s_csamul_cla12_fa8_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand9_11(.a(a[9]), .b(b[11]), .out(s_csamul_cla12_nand9_11));
  fa fa_s_csamul_cla12_fa9_11_out(.a(s_csamul_cla12_nand9_11[0]), .b(s_csamul_cla12_fa10_10_xor1[0]), .cin(s_csamul_cla12_fa9_10_or0[0]), .fa_xor1(s_csamul_cla12_fa9_11_xor1), .fa_or0(s_csamul_cla12_fa9_11_or0));
  nand_gate nand_gate_s_csamul_cla12_nand10_11(.a(a[10]), .b(b[11]), .out(s_csamul_cla12_nand10_11));
  fa fa_s_csamul_cla12_fa10_11_out(.a(s_csamul_cla12_nand10_11[0]), .b(s_csamul_cla12_ha11_10_xor0[0]), .cin(s_csamul_cla12_fa10_10_or0[0]), .fa_xor1(s_csamul_cla12_fa10_11_xor1), .fa_or0(s_csamul_cla12_fa10_11_or0));
  and_gate and_gate_s_csamul_cla12_and11_11(.a(a[11]), .b(b[11]), .out(s_csamul_cla12_and11_11));
  ha ha_s_csamul_cla12_ha11_11_out(.a(s_csamul_cla12_and11_11[0]), .b(s_csamul_cla12_ha11_10_and0[0]), .ha_xor0(s_csamul_cla12_ha11_11_xor0), .ha_and0(s_csamul_cla12_ha11_11_and0));
  assign s_csamul_cla12_u_cla12_a[0] = s_csamul_cla12_fa1_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[1] = s_csamul_cla12_fa2_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[2] = s_csamul_cla12_fa3_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[3] = s_csamul_cla12_fa4_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[4] = s_csamul_cla12_fa5_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[5] = s_csamul_cla12_fa6_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[6] = s_csamul_cla12_fa7_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[7] = s_csamul_cla12_fa8_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[8] = s_csamul_cla12_fa9_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[9] = s_csamul_cla12_fa10_11_xor1[0];
  assign s_csamul_cla12_u_cla12_a[10] = s_csamul_cla12_ha11_11_xor0[0];
  assign s_csamul_cla12_u_cla12_a[11] = 1'b1;
  assign s_csamul_cla12_u_cla12_b[0] = s_csamul_cla12_fa0_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[1] = s_csamul_cla12_fa1_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[2] = s_csamul_cla12_fa2_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[3] = s_csamul_cla12_fa3_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[4] = s_csamul_cla12_fa4_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[5] = s_csamul_cla12_fa5_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[6] = s_csamul_cla12_fa6_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[7] = s_csamul_cla12_fa7_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[8] = s_csamul_cla12_fa8_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[9] = s_csamul_cla12_fa9_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[10] = s_csamul_cla12_fa10_11_or0[0];
  assign s_csamul_cla12_u_cla12_b[11] = s_csamul_cla12_ha11_11_and0[0];
  u_cla12 u_cla12_s_csamul_cla12_u_cla12_out(.a(s_csamul_cla12_u_cla12_a), .b(s_csamul_cla12_u_cla12_b), .u_cla12_out(s_csamul_cla12_u_cla12_out));

  assign s_csamul_cla12_out[0] = s_csamul_cla12_and0_0[0];
  assign s_csamul_cla12_out[1] = s_csamul_cla12_ha0_1_xor0[0];
  assign s_csamul_cla12_out[2] = s_csamul_cla12_fa0_2_xor1[0];
  assign s_csamul_cla12_out[3] = s_csamul_cla12_fa0_3_xor1[0];
  assign s_csamul_cla12_out[4] = s_csamul_cla12_fa0_4_xor1[0];
  assign s_csamul_cla12_out[5] = s_csamul_cla12_fa0_5_xor1[0];
  assign s_csamul_cla12_out[6] = s_csamul_cla12_fa0_6_xor1[0];
  assign s_csamul_cla12_out[7] = s_csamul_cla12_fa0_7_xor1[0];
  assign s_csamul_cla12_out[8] = s_csamul_cla12_fa0_8_xor1[0];
  assign s_csamul_cla12_out[9] = s_csamul_cla12_fa0_9_xor1[0];
  assign s_csamul_cla12_out[10] = s_csamul_cla12_fa0_10_xor1[0];
  assign s_csamul_cla12_out[11] = s_csamul_cla12_fa0_11_xor1[0];
  assign s_csamul_cla12_out[12] = s_csamul_cla12_u_cla12_out[0];
  assign s_csamul_cla12_out[13] = s_csamul_cla12_u_cla12_out[1];
  assign s_csamul_cla12_out[14] = s_csamul_cla12_u_cla12_out[2];
  assign s_csamul_cla12_out[15] = s_csamul_cla12_u_cla12_out[3];
  assign s_csamul_cla12_out[16] = s_csamul_cla12_u_cla12_out[4];
  assign s_csamul_cla12_out[17] = s_csamul_cla12_u_cla12_out[5];
  assign s_csamul_cla12_out[18] = s_csamul_cla12_u_cla12_out[6];
  assign s_csamul_cla12_out[19] = s_csamul_cla12_u_cla12_out[7];
  assign s_csamul_cla12_out[20] = s_csamul_cla12_u_cla12_out[8];
  assign s_csamul_cla12_out[21] = s_csamul_cla12_u_cla12_out[9];
  assign s_csamul_cla12_out[22] = s_csamul_cla12_u_cla12_out[10];
  assign s_csamul_cla12_out[23] = s_csamul_cla12_u_cla12_out[11];
endmodule