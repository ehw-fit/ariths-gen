module u_dadda_cla8(input [7:0] a, input [7:0] b, output [15:0] u_dadda_cla8_out);
  wire u_dadda_cla8_and_6_0;
  wire u_dadda_cla8_and_5_1;
  wire u_dadda_cla8_ha0_xor0;
  wire u_dadda_cla8_ha0_and0;
  wire u_dadda_cla8_and_7_0;
  wire u_dadda_cla8_and_6_1;
  wire u_dadda_cla8_fa0_xor0;
  wire u_dadda_cla8_fa0_and0;
  wire u_dadda_cla8_fa0_xor1;
  wire u_dadda_cla8_fa0_and1;
  wire u_dadda_cla8_fa0_or0;
  wire u_dadda_cla8_and_5_2;
  wire u_dadda_cla8_and_4_3;
  wire u_dadda_cla8_ha1_xor0;
  wire u_dadda_cla8_ha1_and0;
  wire u_dadda_cla8_and_7_1;
  wire u_dadda_cla8_fa1_xor0;
  wire u_dadda_cla8_fa1_and0;
  wire u_dadda_cla8_fa1_xor1;
  wire u_dadda_cla8_fa1_and1;
  wire u_dadda_cla8_fa1_or0;
  wire u_dadda_cla8_and_6_2;
  wire u_dadda_cla8_and_5_3;
  wire u_dadda_cla8_ha2_xor0;
  wire u_dadda_cla8_ha2_and0;
  wire u_dadda_cla8_and_7_2;
  wire u_dadda_cla8_fa2_xor0;
  wire u_dadda_cla8_fa2_and0;
  wire u_dadda_cla8_fa2_xor1;
  wire u_dadda_cla8_fa2_and1;
  wire u_dadda_cla8_fa2_or0;
  wire u_dadda_cla8_and_3_0;
  wire u_dadda_cla8_and_2_1;
  wire u_dadda_cla8_ha3_xor0;
  wire u_dadda_cla8_ha3_and0;
  wire u_dadda_cla8_and_4_0;
  wire u_dadda_cla8_and_3_1;
  wire u_dadda_cla8_fa3_xor0;
  wire u_dadda_cla8_fa3_and0;
  wire u_dadda_cla8_fa3_xor1;
  wire u_dadda_cla8_fa3_and1;
  wire u_dadda_cla8_fa3_or0;
  wire u_dadda_cla8_and_2_2;
  wire u_dadda_cla8_and_1_3;
  wire u_dadda_cla8_ha4_xor0;
  wire u_dadda_cla8_ha4_and0;
  wire u_dadda_cla8_and_5_0;
  wire u_dadda_cla8_fa4_xor0;
  wire u_dadda_cla8_fa4_and0;
  wire u_dadda_cla8_fa4_xor1;
  wire u_dadda_cla8_fa4_and1;
  wire u_dadda_cla8_fa4_or0;
  wire u_dadda_cla8_and_4_1;
  wire u_dadda_cla8_and_3_2;
  wire u_dadda_cla8_and_2_3;
  wire u_dadda_cla8_fa5_xor0;
  wire u_dadda_cla8_fa5_and0;
  wire u_dadda_cla8_fa5_xor1;
  wire u_dadda_cla8_fa5_and1;
  wire u_dadda_cla8_fa5_or0;
  wire u_dadda_cla8_and_1_4;
  wire u_dadda_cla8_and_0_5;
  wire u_dadda_cla8_ha5_xor0;
  wire u_dadda_cla8_ha5_and0;
  wire u_dadda_cla8_fa6_xor0;
  wire u_dadda_cla8_fa6_and0;
  wire u_dadda_cla8_fa6_xor1;
  wire u_dadda_cla8_fa6_and1;
  wire u_dadda_cla8_fa6_or0;
  wire u_dadda_cla8_and_4_2;
  wire u_dadda_cla8_and_3_3;
  wire u_dadda_cla8_and_2_4;
  wire u_dadda_cla8_fa7_xor0;
  wire u_dadda_cla8_fa7_and0;
  wire u_dadda_cla8_fa7_xor1;
  wire u_dadda_cla8_fa7_and1;
  wire u_dadda_cla8_fa7_or0;
  wire u_dadda_cla8_and_1_5;
  wire u_dadda_cla8_and_0_6;
  wire u_dadda_cla8_fa8_xor0;
  wire u_dadda_cla8_fa8_and0;
  wire u_dadda_cla8_fa8_xor1;
  wire u_dadda_cla8_fa8_and1;
  wire u_dadda_cla8_fa8_or0;
  wire u_dadda_cla8_fa9_xor0;
  wire u_dadda_cla8_fa9_and0;
  wire u_dadda_cla8_fa9_xor1;
  wire u_dadda_cla8_fa9_and1;
  wire u_dadda_cla8_fa9_or0;
  wire u_dadda_cla8_and_3_4;
  wire u_dadda_cla8_and_2_5;
  wire u_dadda_cla8_and_1_6;
  wire u_dadda_cla8_fa10_xor0;
  wire u_dadda_cla8_fa10_and0;
  wire u_dadda_cla8_fa10_xor1;
  wire u_dadda_cla8_fa10_and1;
  wire u_dadda_cla8_fa10_or0;
  wire u_dadda_cla8_and_0_7;
  wire u_dadda_cla8_fa11_xor0;
  wire u_dadda_cla8_fa11_and0;
  wire u_dadda_cla8_fa11_xor1;
  wire u_dadda_cla8_fa11_and1;
  wire u_dadda_cla8_fa11_or0;
  wire u_dadda_cla8_fa12_xor0;
  wire u_dadda_cla8_fa12_and0;
  wire u_dadda_cla8_fa12_xor1;
  wire u_dadda_cla8_fa12_and1;
  wire u_dadda_cla8_fa12_or0;
  wire u_dadda_cla8_and_4_4;
  wire u_dadda_cla8_and_3_5;
  wire u_dadda_cla8_and_2_6;
  wire u_dadda_cla8_fa13_xor0;
  wire u_dadda_cla8_fa13_and0;
  wire u_dadda_cla8_fa13_xor1;
  wire u_dadda_cla8_fa13_and1;
  wire u_dadda_cla8_fa13_or0;
  wire u_dadda_cla8_and_1_7;
  wire u_dadda_cla8_fa14_xor0;
  wire u_dadda_cla8_fa14_and0;
  wire u_dadda_cla8_fa14_xor1;
  wire u_dadda_cla8_fa14_and1;
  wire u_dadda_cla8_fa14_or0;
  wire u_dadda_cla8_fa15_xor0;
  wire u_dadda_cla8_fa15_and0;
  wire u_dadda_cla8_fa15_xor1;
  wire u_dadda_cla8_fa15_and1;
  wire u_dadda_cla8_fa15_or0;
  wire u_dadda_cla8_and_6_3;
  wire u_dadda_cla8_and_5_4;
  wire u_dadda_cla8_and_4_5;
  wire u_dadda_cla8_fa16_xor0;
  wire u_dadda_cla8_fa16_and0;
  wire u_dadda_cla8_fa16_xor1;
  wire u_dadda_cla8_fa16_and1;
  wire u_dadda_cla8_fa16_or0;
  wire u_dadda_cla8_and_3_6;
  wire u_dadda_cla8_and_2_7;
  wire u_dadda_cla8_fa17_xor0;
  wire u_dadda_cla8_fa17_and0;
  wire u_dadda_cla8_fa17_xor1;
  wire u_dadda_cla8_fa17_and1;
  wire u_dadda_cla8_fa17_or0;
  wire u_dadda_cla8_fa18_xor0;
  wire u_dadda_cla8_fa18_and0;
  wire u_dadda_cla8_fa18_xor1;
  wire u_dadda_cla8_fa18_and1;
  wire u_dadda_cla8_fa18_or0;
  wire u_dadda_cla8_and_7_3;
  wire u_dadda_cla8_and_6_4;
  wire u_dadda_cla8_fa19_xor0;
  wire u_dadda_cla8_fa19_and0;
  wire u_dadda_cla8_fa19_xor1;
  wire u_dadda_cla8_fa19_and1;
  wire u_dadda_cla8_fa19_or0;
  wire u_dadda_cla8_and_5_5;
  wire u_dadda_cla8_and_4_6;
  wire u_dadda_cla8_and_3_7;
  wire u_dadda_cla8_fa20_xor0;
  wire u_dadda_cla8_fa20_and0;
  wire u_dadda_cla8_fa20_xor1;
  wire u_dadda_cla8_fa20_and1;
  wire u_dadda_cla8_fa20_or0;
  wire u_dadda_cla8_fa21_xor0;
  wire u_dadda_cla8_fa21_and0;
  wire u_dadda_cla8_fa21_xor1;
  wire u_dadda_cla8_fa21_and1;
  wire u_dadda_cla8_fa21_or0;
  wire u_dadda_cla8_and_7_4;
  wire u_dadda_cla8_and_6_5;
  wire u_dadda_cla8_and_5_6;
  wire u_dadda_cla8_fa22_xor0;
  wire u_dadda_cla8_fa22_and0;
  wire u_dadda_cla8_fa22_xor1;
  wire u_dadda_cla8_fa22_and1;
  wire u_dadda_cla8_fa22_or0;
  wire u_dadda_cla8_and_7_5;
  wire u_dadda_cla8_fa23_xor0;
  wire u_dadda_cla8_fa23_and0;
  wire u_dadda_cla8_fa23_xor1;
  wire u_dadda_cla8_fa23_and1;
  wire u_dadda_cla8_fa23_or0;
  wire u_dadda_cla8_and_2_0;
  wire u_dadda_cla8_and_1_1;
  wire u_dadda_cla8_ha6_xor0;
  wire u_dadda_cla8_ha6_and0;
  wire u_dadda_cla8_and_1_2;
  wire u_dadda_cla8_and_0_3;
  wire u_dadda_cla8_fa24_xor0;
  wire u_dadda_cla8_fa24_and0;
  wire u_dadda_cla8_fa24_xor1;
  wire u_dadda_cla8_fa24_and1;
  wire u_dadda_cla8_fa24_or0;
  wire u_dadda_cla8_and_0_4;
  wire u_dadda_cla8_fa25_xor0;
  wire u_dadda_cla8_fa25_and0;
  wire u_dadda_cla8_fa25_xor1;
  wire u_dadda_cla8_fa25_and1;
  wire u_dadda_cla8_fa25_or0;
  wire u_dadda_cla8_fa26_xor0;
  wire u_dadda_cla8_fa26_and0;
  wire u_dadda_cla8_fa26_xor1;
  wire u_dadda_cla8_fa26_and1;
  wire u_dadda_cla8_fa26_or0;
  wire u_dadda_cla8_fa27_xor0;
  wire u_dadda_cla8_fa27_and0;
  wire u_dadda_cla8_fa27_xor1;
  wire u_dadda_cla8_fa27_and1;
  wire u_dadda_cla8_fa27_or0;
  wire u_dadda_cla8_fa28_xor0;
  wire u_dadda_cla8_fa28_and0;
  wire u_dadda_cla8_fa28_xor1;
  wire u_dadda_cla8_fa28_and1;
  wire u_dadda_cla8_fa28_or0;
  wire u_dadda_cla8_fa29_xor0;
  wire u_dadda_cla8_fa29_and0;
  wire u_dadda_cla8_fa29_xor1;
  wire u_dadda_cla8_fa29_and1;
  wire u_dadda_cla8_fa29_or0;
  wire u_dadda_cla8_fa30_xor0;
  wire u_dadda_cla8_fa30_and0;
  wire u_dadda_cla8_fa30_xor1;
  wire u_dadda_cla8_fa30_and1;
  wire u_dadda_cla8_fa30_or0;
  wire u_dadda_cla8_fa31_xor0;
  wire u_dadda_cla8_fa31_and0;
  wire u_dadda_cla8_fa31_xor1;
  wire u_dadda_cla8_fa31_and1;
  wire u_dadda_cla8_fa31_or0;
  wire u_dadda_cla8_and_4_7;
  wire u_dadda_cla8_fa32_xor0;
  wire u_dadda_cla8_fa32_and0;
  wire u_dadda_cla8_fa32_xor1;
  wire u_dadda_cla8_fa32_and1;
  wire u_dadda_cla8_fa32_or0;
  wire u_dadda_cla8_and_6_6;
  wire u_dadda_cla8_and_5_7;
  wire u_dadda_cla8_fa33_xor0;
  wire u_dadda_cla8_fa33_and0;
  wire u_dadda_cla8_fa33_xor1;
  wire u_dadda_cla8_fa33_and1;
  wire u_dadda_cla8_fa33_or0;
  wire u_dadda_cla8_and_7_6;
  wire u_dadda_cla8_fa34_xor0;
  wire u_dadda_cla8_fa34_and0;
  wire u_dadda_cla8_fa34_xor1;
  wire u_dadda_cla8_fa34_and1;
  wire u_dadda_cla8_fa34_or0;
  wire u_dadda_cla8_and_0_0;
  wire u_dadda_cla8_and_1_0;
  wire u_dadda_cla8_and_0_2;
  wire u_dadda_cla8_and_6_7;
  wire u_dadda_cla8_and_0_1;
  wire u_dadda_cla8_and_7_7;
  wire u_dadda_cla8_u_cla14_pg_logic0_or0;
  wire u_dadda_cla8_u_cla14_pg_logic0_and0;
  wire u_dadda_cla8_u_cla14_pg_logic0_xor0;
  wire u_dadda_cla8_u_cla14_pg_logic1_or0;
  wire u_dadda_cla8_u_cla14_pg_logic1_and0;
  wire u_dadda_cla8_u_cla14_pg_logic1_xor0;
  wire u_dadda_cla8_u_cla14_xor1;
  wire u_dadda_cla8_u_cla14_and0;
  wire u_dadda_cla8_u_cla14_or0;
  wire u_dadda_cla8_u_cla14_pg_logic2_or0;
  wire u_dadda_cla8_u_cla14_pg_logic2_and0;
  wire u_dadda_cla8_u_cla14_pg_logic2_xor0;
  wire u_dadda_cla8_u_cla14_xor2;
  wire u_dadda_cla8_u_cla14_and1;
  wire u_dadda_cla8_u_cla14_and2;
  wire u_dadda_cla8_u_cla14_and3;
  wire u_dadda_cla8_u_cla14_and4;
  wire u_dadda_cla8_u_cla14_or1;
  wire u_dadda_cla8_u_cla14_or2;
  wire u_dadda_cla8_u_cla14_pg_logic3_or0;
  wire u_dadda_cla8_u_cla14_pg_logic3_and0;
  wire u_dadda_cla8_u_cla14_pg_logic3_xor0;
  wire u_dadda_cla8_u_cla14_xor3;
  wire u_dadda_cla8_u_cla14_and5;
  wire u_dadda_cla8_u_cla14_and6;
  wire u_dadda_cla8_u_cla14_and7;
  wire u_dadda_cla8_u_cla14_and8;
  wire u_dadda_cla8_u_cla14_and9;
  wire u_dadda_cla8_u_cla14_and10;
  wire u_dadda_cla8_u_cla14_and11;
  wire u_dadda_cla8_u_cla14_or3;
  wire u_dadda_cla8_u_cla14_or4;
  wire u_dadda_cla8_u_cla14_or5;
  wire u_dadda_cla8_u_cla14_pg_logic4_or0;
  wire u_dadda_cla8_u_cla14_pg_logic4_and0;
  wire u_dadda_cla8_u_cla14_pg_logic4_xor0;
  wire u_dadda_cla8_u_cla14_xor4;
  wire u_dadda_cla8_u_cla14_and12;
  wire u_dadda_cla8_u_cla14_or6;
  wire u_dadda_cla8_u_cla14_pg_logic5_or0;
  wire u_dadda_cla8_u_cla14_pg_logic5_and0;
  wire u_dadda_cla8_u_cla14_pg_logic5_xor0;
  wire u_dadda_cla8_u_cla14_xor5;
  wire u_dadda_cla8_u_cla14_and13;
  wire u_dadda_cla8_u_cla14_and14;
  wire u_dadda_cla8_u_cla14_and15;
  wire u_dadda_cla8_u_cla14_or7;
  wire u_dadda_cla8_u_cla14_or8;
  wire u_dadda_cla8_u_cla14_pg_logic6_or0;
  wire u_dadda_cla8_u_cla14_pg_logic6_and0;
  wire u_dadda_cla8_u_cla14_pg_logic6_xor0;
  wire u_dadda_cla8_u_cla14_xor6;
  wire u_dadda_cla8_u_cla14_and16;
  wire u_dadda_cla8_u_cla14_and17;
  wire u_dadda_cla8_u_cla14_and18;
  wire u_dadda_cla8_u_cla14_and19;
  wire u_dadda_cla8_u_cla14_and20;
  wire u_dadda_cla8_u_cla14_and21;
  wire u_dadda_cla8_u_cla14_or9;
  wire u_dadda_cla8_u_cla14_or10;
  wire u_dadda_cla8_u_cla14_or11;
  wire u_dadda_cla8_u_cla14_pg_logic7_or0;
  wire u_dadda_cla8_u_cla14_pg_logic7_and0;
  wire u_dadda_cla8_u_cla14_pg_logic7_xor0;
  wire u_dadda_cla8_u_cla14_xor7;
  wire u_dadda_cla8_u_cla14_and22;
  wire u_dadda_cla8_u_cla14_and23;
  wire u_dadda_cla8_u_cla14_and24;
  wire u_dadda_cla8_u_cla14_and25;
  wire u_dadda_cla8_u_cla14_and26;
  wire u_dadda_cla8_u_cla14_and27;
  wire u_dadda_cla8_u_cla14_and28;
  wire u_dadda_cla8_u_cla14_and29;
  wire u_dadda_cla8_u_cla14_and30;
  wire u_dadda_cla8_u_cla14_and31;
  wire u_dadda_cla8_u_cla14_or12;
  wire u_dadda_cla8_u_cla14_or13;
  wire u_dadda_cla8_u_cla14_or14;
  wire u_dadda_cla8_u_cla14_or15;
  wire u_dadda_cla8_u_cla14_pg_logic8_or0;
  wire u_dadda_cla8_u_cla14_pg_logic8_and0;
  wire u_dadda_cla8_u_cla14_pg_logic8_xor0;
  wire u_dadda_cla8_u_cla14_xor8;
  wire u_dadda_cla8_u_cla14_and32;
  wire u_dadda_cla8_u_cla14_or16;
  wire u_dadda_cla8_u_cla14_pg_logic9_or0;
  wire u_dadda_cla8_u_cla14_pg_logic9_and0;
  wire u_dadda_cla8_u_cla14_pg_logic9_xor0;
  wire u_dadda_cla8_u_cla14_xor9;
  wire u_dadda_cla8_u_cla14_and33;
  wire u_dadda_cla8_u_cla14_and34;
  wire u_dadda_cla8_u_cla14_and35;
  wire u_dadda_cla8_u_cla14_or17;
  wire u_dadda_cla8_u_cla14_or18;
  wire u_dadda_cla8_u_cla14_pg_logic10_or0;
  wire u_dadda_cla8_u_cla14_pg_logic10_and0;
  wire u_dadda_cla8_u_cla14_pg_logic10_xor0;
  wire u_dadda_cla8_u_cla14_xor10;
  wire u_dadda_cla8_u_cla14_and36;
  wire u_dadda_cla8_u_cla14_and37;
  wire u_dadda_cla8_u_cla14_and38;
  wire u_dadda_cla8_u_cla14_and39;
  wire u_dadda_cla8_u_cla14_and40;
  wire u_dadda_cla8_u_cla14_and41;
  wire u_dadda_cla8_u_cla14_or19;
  wire u_dadda_cla8_u_cla14_or20;
  wire u_dadda_cla8_u_cla14_or21;
  wire u_dadda_cla8_u_cla14_pg_logic11_or0;
  wire u_dadda_cla8_u_cla14_pg_logic11_and0;
  wire u_dadda_cla8_u_cla14_pg_logic11_xor0;
  wire u_dadda_cla8_u_cla14_xor11;
  wire u_dadda_cla8_u_cla14_and42;
  wire u_dadda_cla8_u_cla14_and43;
  wire u_dadda_cla8_u_cla14_and44;
  wire u_dadda_cla8_u_cla14_and45;
  wire u_dadda_cla8_u_cla14_and46;
  wire u_dadda_cla8_u_cla14_and47;
  wire u_dadda_cla8_u_cla14_and48;
  wire u_dadda_cla8_u_cla14_and49;
  wire u_dadda_cla8_u_cla14_and50;
  wire u_dadda_cla8_u_cla14_and51;
  wire u_dadda_cla8_u_cla14_or22;
  wire u_dadda_cla8_u_cla14_or23;
  wire u_dadda_cla8_u_cla14_or24;
  wire u_dadda_cla8_u_cla14_or25;
  wire u_dadda_cla8_u_cla14_pg_logic12_or0;
  wire u_dadda_cla8_u_cla14_pg_logic12_and0;
  wire u_dadda_cla8_u_cla14_pg_logic12_xor0;
  wire u_dadda_cla8_u_cla14_xor12;
  wire u_dadda_cla8_u_cla14_and52;
  wire u_dadda_cla8_u_cla14_or26;
  wire u_dadda_cla8_u_cla14_pg_logic13_or0;
  wire u_dadda_cla8_u_cla14_pg_logic13_and0;
  wire u_dadda_cla8_u_cla14_pg_logic13_xor0;
  wire u_dadda_cla8_u_cla14_xor13;
  wire u_dadda_cla8_u_cla14_and53;
  wire u_dadda_cla8_u_cla14_and54;
  wire u_dadda_cla8_u_cla14_and55;
  wire u_dadda_cla8_u_cla14_or27;
  wire u_dadda_cla8_u_cla14_or28;

  assign u_dadda_cla8_and_6_0 = a[6] & b[0];
  assign u_dadda_cla8_and_5_1 = a[5] & b[1];
  assign u_dadda_cla8_ha0_xor0 = u_dadda_cla8_and_6_0 ^ u_dadda_cla8_and_5_1;
  assign u_dadda_cla8_ha0_and0 = u_dadda_cla8_and_6_0 & u_dadda_cla8_and_5_1;
  assign u_dadda_cla8_and_7_0 = a[7] & b[0];
  assign u_dadda_cla8_and_6_1 = a[6] & b[1];
  assign u_dadda_cla8_fa0_xor0 = u_dadda_cla8_ha0_and0 ^ u_dadda_cla8_and_7_0;
  assign u_dadda_cla8_fa0_and0 = u_dadda_cla8_ha0_and0 & u_dadda_cla8_and_7_0;
  assign u_dadda_cla8_fa0_xor1 = u_dadda_cla8_fa0_xor0 ^ u_dadda_cla8_and_6_1;
  assign u_dadda_cla8_fa0_and1 = u_dadda_cla8_fa0_xor0 & u_dadda_cla8_and_6_1;
  assign u_dadda_cla8_fa0_or0 = u_dadda_cla8_fa0_and0 | u_dadda_cla8_fa0_and1;
  assign u_dadda_cla8_and_5_2 = a[5] & b[2];
  assign u_dadda_cla8_and_4_3 = a[4] & b[3];
  assign u_dadda_cla8_ha1_xor0 = u_dadda_cla8_and_5_2 ^ u_dadda_cla8_and_4_3;
  assign u_dadda_cla8_ha1_and0 = u_dadda_cla8_and_5_2 & u_dadda_cla8_and_4_3;
  assign u_dadda_cla8_and_7_1 = a[7] & b[1];
  assign u_dadda_cla8_fa1_xor0 = u_dadda_cla8_ha1_and0 ^ u_dadda_cla8_fa0_or0;
  assign u_dadda_cla8_fa1_and0 = u_dadda_cla8_ha1_and0 & u_dadda_cla8_fa0_or0;
  assign u_dadda_cla8_fa1_xor1 = u_dadda_cla8_fa1_xor0 ^ u_dadda_cla8_and_7_1;
  assign u_dadda_cla8_fa1_and1 = u_dadda_cla8_fa1_xor0 & u_dadda_cla8_and_7_1;
  assign u_dadda_cla8_fa1_or0 = u_dadda_cla8_fa1_and0 | u_dadda_cla8_fa1_and1;
  assign u_dadda_cla8_and_6_2 = a[6] & b[2];
  assign u_dadda_cla8_and_5_3 = a[5] & b[3];
  assign u_dadda_cla8_ha2_xor0 = u_dadda_cla8_and_6_2 ^ u_dadda_cla8_and_5_3;
  assign u_dadda_cla8_ha2_and0 = u_dadda_cla8_and_6_2 & u_dadda_cla8_and_5_3;
  assign u_dadda_cla8_and_7_2 = a[7] & b[2];
  assign u_dadda_cla8_fa2_xor0 = u_dadda_cla8_ha2_and0 ^ u_dadda_cla8_fa1_or0;
  assign u_dadda_cla8_fa2_and0 = u_dadda_cla8_ha2_and0 & u_dadda_cla8_fa1_or0;
  assign u_dadda_cla8_fa2_xor1 = u_dadda_cla8_fa2_xor0 ^ u_dadda_cla8_and_7_2;
  assign u_dadda_cla8_fa2_and1 = u_dadda_cla8_fa2_xor0 & u_dadda_cla8_and_7_2;
  assign u_dadda_cla8_fa2_or0 = u_dadda_cla8_fa2_and0 | u_dadda_cla8_fa2_and1;
  assign u_dadda_cla8_and_3_0 = a[3] & b[0];
  assign u_dadda_cla8_and_2_1 = a[2] & b[1];
  assign u_dadda_cla8_ha3_xor0 = u_dadda_cla8_and_3_0 ^ u_dadda_cla8_and_2_1;
  assign u_dadda_cla8_ha3_and0 = u_dadda_cla8_and_3_0 & u_dadda_cla8_and_2_1;
  assign u_dadda_cla8_and_4_0 = a[4] & b[0];
  assign u_dadda_cla8_and_3_1 = a[3] & b[1];
  assign u_dadda_cla8_fa3_xor0 = u_dadda_cla8_ha3_and0 ^ u_dadda_cla8_and_4_0;
  assign u_dadda_cla8_fa3_and0 = u_dadda_cla8_ha3_and0 & u_dadda_cla8_and_4_0;
  assign u_dadda_cla8_fa3_xor1 = u_dadda_cla8_fa3_xor0 ^ u_dadda_cla8_and_3_1;
  assign u_dadda_cla8_fa3_and1 = u_dadda_cla8_fa3_xor0 & u_dadda_cla8_and_3_1;
  assign u_dadda_cla8_fa3_or0 = u_dadda_cla8_fa3_and0 | u_dadda_cla8_fa3_and1;
  assign u_dadda_cla8_and_2_2 = a[2] & b[2];
  assign u_dadda_cla8_and_1_3 = a[1] & b[3];
  assign u_dadda_cla8_ha4_xor0 = u_dadda_cla8_and_2_2 ^ u_dadda_cla8_and_1_3;
  assign u_dadda_cla8_ha4_and0 = u_dadda_cla8_and_2_2 & u_dadda_cla8_and_1_3;
  assign u_dadda_cla8_and_5_0 = a[5] & b[0];
  assign u_dadda_cla8_fa4_xor0 = u_dadda_cla8_ha4_and0 ^ u_dadda_cla8_fa3_or0;
  assign u_dadda_cla8_fa4_and0 = u_dadda_cla8_ha4_and0 & u_dadda_cla8_fa3_or0;
  assign u_dadda_cla8_fa4_xor1 = u_dadda_cla8_fa4_xor0 ^ u_dadda_cla8_and_5_0;
  assign u_dadda_cla8_fa4_and1 = u_dadda_cla8_fa4_xor0 & u_dadda_cla8_and_5_0;
  assign u_dadda_cla8_fa4_or0 = u_dadda_cla8_fa4_and0 | u_dadda_cla8_fa4_and1;
  assign u_dadda_cla8_and_4_1 = a[4] & b[1];
  assign u_dadda_cla8_and_3_2 = a[3] & b[2];
  assign u_dadda_cla8_and_2_3 = a[2] & b[3];
  assign u_dadda_cla8_fa5_xor0 = u_dadda_cla8_and_4_1 ^ u_dadda_cla8_and_3_2;
  assign u_dadda_cla8_fa5_and0 = u_dadda_cla8_and_4_1 & u_dadda_cla8_and_3_2;
  assign u_dadda_cla8_fa5_xor1 = u_dadda_cla8_fa5_xor0 ^ u_dadda_cla8_and_2_3;
  assign u_dadda_cla8_fa5_and1 = u_dadda_cla8_fa5_xor0 & u_dadda_cla8_and_2_3;
  assign u_dadda_cla8_fa5_or0 = u_dadda_cla8_fa5_and0 | u_dadda_cla8_fa5_and1;
  assign u_dadda_cla8_and_1_4 = a[1] & b[4];
  assign u_dadda_cla8_and_0_5 = a[0] & b[5];
  assign u_dadda_cla8_ha5_xor0 = u_dadda_cla8_and_1_4 ^ u_dadda_cla8_and_0_5;
  assign u_dadda_cla8_ha5_and0 = u_dadda_cla8_and_1_4 & u_dadda_cla8_and_0_5;
  assign u_dadda_cla8_fa6_xor0 = u_dadda_cla8_ha5_and0 ^ u_dadda_cla8_fa5_or0;
  assign u_dadda_cla8_fa6_and0 = u_dadda_cla8_ha5_and0 & u_dadda_cla8_fa5_or0;
  assign u_dadda_cla8_fa6_xor1 = u_dadda_cla8_fa6_xor0 ^ u_dadda_cla8_fa4_or0;
  assign u_dadda_cla8_fa6_and1 = u_dadda_cla8_fa6_xor0 & u_dadda_cla8_fa4_or0;
  assign u_dadda_cla8_fa6_or0 = u_dadda_cla8_fa6_and0 | u_dadda_cla8_fa6_and1;
  assign u_dadda_cla8_and_4_2 = a[4] & b[2];
  assign u_dadda_cla8_and_3_3 = a[3] & b[3];
  assign u_dadda_cla8_and_2_4 = a[2] & b[4];
  assign u_dadda_cla8_fa7_xor0 = u_dadda_cla8_and_4_2 ^ u_dadda_cla8_and_3_3;
  assign u_dadda_cla8_fa7_and0 = u_dadda_cla8_and_4_2 & u_dadda_cla8_and_3_3;
  assign u_dadda_cla8_fa7_xor1 = u_dadda_cla8_fa7_xor0 ^ u_dadda_cla8_and_2_4;
  assign u_dadda_cla8_fa7_and1 = u_dadda_cla8_fa7_xor0 & u_dadda_cla8_and_2_4;
  assign u_dadda_cla8_fa7_or0 = u_dadda_cla8_fa7_and0 | u_dadda_cla8_fa7_and1;
  assign u_dadda_cla8_and_1_5 = a[1] & b[5];
  assign u_dadda_cla8_and_0_6 = a[0] & b[6];
  assign u_dadda_cla8_fa8_xor0 = u_dadda_cla8_and_1_5 ^ u_dadda_cla8_and_0_6;
  assign u_dadda_cla8_fa8_and0 = u_dadda_cla8_and_1_5 & u_dadda_cla8_and_0_6;
  assign u_dadda_cla8_fa8_xor1 = u_dadda_cla8_fa8_xor0 ^ u_dadda_cla8_ha0_xor0;
  assign u_dadda_cla8_fa8_and1 = u_dadda_cla8_fa8_xor0 & u_dadda_cla8_ha0_xor0;
  assign u_dadda_cla8_fa8_or0 = u_dadda_cla8_fa8_and0 | u_dadda_cla8_fa8_and1;
  assign u_dadda_cla8_fa9_xor0 = u_dadda_cla8_fa8_or0 ^ u_dadda_cla8_fa7_or0;
  assign u_dadda_cla8_fa9_and0 = u_dadda_cla8_fa8_or0 & u_dadda_cla8_fa7_or0;
  assign u_dadda_cla8_fa9_xor1 = u_dadda_cla8_fa9_xor0 ^ u_dadda_cla8_fa6_or0;
  assign u_dadda_cla8_fa9_and1 = u_dadda_cla8_fa9_xor0 & u_dadda_cla8_fa6_or0;
  assign u_dadda_cla8_fa9_or0 = u_dadda_cla8_fa9_and0 | u_dadda_cla8_fa9_and1;
  assign u_dadda_cla8_and_3_4 = a[3] & b[4];
  assign u_dadda_cla8_and_2_5 = a[2] & b[5];
  assign u_dadda_cla8_and_1_6 = a[1] & b[6];
  assign u_dadda_cla8_fa10_xor0 = u_dadda_cla8_and_3_4 ^ u_dadda_cla8_and_2_5;
  assign u_dadda_cla8_fa10_and0 = u_dadda_cla8_and_3_4 & u_dadda_cla8_and_2_5;
  assign u_dadda_cla8_fa10_xor1 = u_dadda_cla8_fa10_xor0 ^ u_dadda_cla8_and_1_6;
  assign u_dadda_cla8_fa10_and1 = u_dadda_cla8_fa10_xor0 & u_dadda_cla8_and_1_6;
  assign u_dadda_cla8_fa10_or0 = u_dadda_cla8_fa10_and0 | u_dadda_cla8_fa10_and1;
  assign u_dadda_cla8_and_0_7 = a[0] & b[7];
  assign u_dadda_cla8_fa11_xor0 = u_dadda_cla8_and_0_7 ^ u_dadda_cla8_fa0_xor1;
  assign u_dadda_cla8_fa11_and0 = u_dadda_cla8_and_0_7 & u_dadda_cla8_fa0_xor1;
  assign u_dadda_cla8_fa11_xor1 = u_dadda_cla8_fa11_xor0 ^ u_dadda_cla8_ha1_xor0;
  assign u_dadda_cla8_fa11_and1 = u_dadda_cla8_fa11_xor0 & u_dadda_cla8_ha1_xor0;
  assign u_dadda_cla8_fa11_or0 = u_dadda_cla8_fa11_and0 | u_dadda_cla8_fa11_and1;
  assign u_dadda_cla8_fa12_xor0 = u_dadda_cla8_fa11_or0 ^ u_dadda_cla8_fa10_or0;
  assign u_dadda_cla8_fa12_and0 = u_dadda_cla8_fa11_or0 & u_dadda_cla8_fa10_or0;
  assign u_dadda_cla8_fa12_xor1 = u_dadda_cla8_fa12_xor0 ^ u_dadda_cla8_fa9_or0;
  assign u_dadda_cla8_fa12_and1 = u_dadda_cla8_fa12_xor0 & u_dadda_cla8_fa9_or0;
  assign u_dadda_cla8_fa12_or0 = u_dadda_cla8_fa12_and0 | u_dadda_cla8_fa12_and1;
  assign u_dadda_cla8_and_4_4 = a[4] & b[4];
  assign u_dadda_cla8_and_3_5 = a[3] & b[5];
  assign u_dadda_cla8_and_2_6 = a[2] & b[6];
  assign u_dadda_cla8_fa13_xor0 = u_dadda_cla8_and_4_4 ^ u_dadda_cla8_and_3_5;
  assign u_dadda_cla8_fa13_and0 = u_dadda_cla8_and_4_4 & u_dadda_cla8_and_3_5;
  assign u_dadda_cla8_fa13_xor1 = u_dadda_cla8_fa13_xor0 ^ u_dadda_cla8_and_2_6;
  assign u_dadda_cla8_fa13_and1 = u_dadda_cla8_fa13_xor0 & u_dadda_cla8_and_2_6;
  assign u_dadda_cla8_fa13_or0 = u_dadda_cla8_fa13_and0 | u_dadda_cla8_fa13_and1;
  assign u_dadda_cla8_and_1_7 = a[1] & b[7];
  assign u_dadda_cla8_fa14_xor0 = u_dadda_cla8_and_1_7 ^ u_dadda_cla8_fa1_xor1;
  assign u_dadda_cla8_fa14_and0 = u_dadda_cla8_and_1_7 & u_dadda_cla8_fa1_xor1;
  assign u_dadda_cla8_fa14_xor1 = u_dadda_cla8_fa14_xor0 ^ u_dadda_cla8_ha2_xor0;
  assign u_dadda_cla8_fa14_and1 = u_dadda_cla8_fa14_xor0 & u_dadda_cla8_ha2_xor0;
  assign u_dadda_cla8_fa14_or0 = u_dadda_cla8_fa14_and0 | u_dadda_cla8_fa14_and1;
  assign u_dadda_cla8_fa15_xor0 = u_dadda_cla8_fa14_or0 ^ u_dadda_cla8_fa13_or0;
  assign u_dadda_cla8_fa15_and0 = u_dadda_cla8_fa14_or0 & u_dadda_cla8_fa13_or0;
  assign u_dadda_cla8_fa15_xor1 = u_dadda_cla8_fa15_xor0 ^ u_dadda_cla8_fa12_or0;
  assign u_dadda_cla8_fa15_and1 = u_dadda_cla8_fa15_xor0 & u_dadda_cla8_fa12_or0;
  assign u_dadda_cla8_fa15_or0 = u_dadda_cla8_fa15_and0 | u_dadda_cla8_fa15_and1;
  assign u_dadda_cla8_and_6_3 = a[6] & b[3];
  assign u_dadda_cla8_and_5_4 = a[5] & b[4];
  assign u_dadda_cla8_and_4_5 = a[4] & b[5];
  assign u_dadda_cla8_fa16_xor0 = u_dadda_cla8_and_6_3 ^ u_dadda_cla8_and_5_4;
  assign u_dadda_cla8_fa16_and0 = u_dadda_cla8_and_6_3 & u_dadda_cla8_and_5_4;
  assign u_dadda_cla8_fa16_xor1 = u_dadda_cla8_fa16_xor0 ^ u_dadda_cla8_and_4_5;
  assign u_dadda_cla8_fa16_and1 = u_dadda_cla8_fa16_xor0 & u_dadda_cla8_and_4_5;
  assign u_dadda_cla8_fa16_or0 = u_dadda_cla8_fa16_and0 | u_dadda_cla8_fa16_and1;
  assign u_dadda_cla8_and_3_6 = a[3] & b[6];
  assign u_dadda_cla8_and_2_7 = a[2] & b[7];
  assign u_dadda_cla8_fa17_xor0 = u_dadda_cla8_and_3_6 ^ u_dadda_cla8_and_2_7;
  assign u_dadda_cla8_fa17_and0 = u_dadda_cla8_and_3_6 & u_dadda_cla8_and_2_7;
  assign u_dadda_cla8_fa17_xor1 = u_dadda_cla8_fa17_xor0 ^ u_dadda_cla8_fa2_xor1;
  assign u_dadda_cla8_fa17_and1 = u_dadda_cla8_fa17_xor0 & u_dadda_cla8_fa2_xor1;
  assign u_dadda_cla8_fa17_or0 = u_dadda_cla8_fa17_and0 | u_dadda_cla8_fa17_and1;
  assign u_dadda_cla8_fa18_xor0 = u_dadda_cla8_fa17_or0 ^ u_dadda_cla8_fa16_or0;
  assign u_dadda_cla8_fa18_and0 = u_dadda_cla8_fa17_or0 & u_dadda_cla8_fa16_or0;
  assign u_dadda_cla8_fa18_xor1 = u_dadda_cla8_fa18_xor0 ^ u_dadda_cla8_fa15_or0;
  assign u_dadda_cla8_fa18_and1 = u_dadda_cla8_fa18_xor0 & u_dadda_cla8_fa15_or0;
  assign u_dadda_cla8_fa18_or0 = u_dadda_cla8_fa18_and0 | u_dadda_cla8_fa18_and1;
  assign u_dadda_cla8_and_7_3 = a[7] & b[3];
  assign u_dadda_cla8_and_6_4 = a[6] & b[4];
  assign u_dadda_cla8_fa19_xor0 = u_dadda_cla8_fa2_or0 ^ u_dadda_cla8_and_7_3;
  assign u_dadda_cla8_fa19_and0 = u_dadda_cla8_fa2_or0 & u_dadda_cla8_and_7_3;
  assign u_dadda_cla8_fa19_xor1 = u_dadda_cla8_fa19_xor0 ^ u_dadda_cla8_and_6_4;
  assign u_dadda_cla8_fa19_and1 = u_dadda_cla8_fa19_xor0 & u_dadda_cla8_and_6_4;
  assign u_dadda_cla8_fa19_or0 = u_dadda_cla8_fa19_and0 | u_dadda_cla8_fa19_and1;
  assign u_dadda_cla8_and_5_5 = a[5] & b[5];
  assign u_dadda_cla8_and_4_6 = a[4] & b[6];
  assign u_dadda_cla8_and_3_7 = a[3] & b[7];
  assign u_dadda_cla8_fa20_xor0 = u_dadda_cla8_and_5_5 ^ u_dadda_cla8_and_4_6;
  assign u_dadda_cla8_fa20_and0 = u_dadda_cla8_and_5_5 & u_dadda_cla8_and_4_6;
  assign u_dadda_cla8_fa20_xor1 = u_dadda_cla8_fa20_xor0 ^ u_dadda_cla8_and_3_7;
  assign u_dadda_cla8_fa20_and1 = u_dadda_cla8_fa20_xor0 & u_dadda_cla8_and_3_7;
  assign u_dadda_cla8_fa20_or0 = u_dadda_cla8_fa20_and0 | u_dadda_cla8_fa20_and1;
  assign u_dadda_cla8_fa21_xor0 = u_dadda_cla8_fa20_or0 ^ u_dadda_cla8_fa19_or0;
  assign u_dadda_cla8_fa21_and0 = u_dadda_cla8_fa20_or0 & u_dadda_cla8_fa19_or0;
  assign u_dadda_cla8_fa21_xor1 = u_dadda_cla8_fa21_xor0 ^ u_dadda_cla8_fa18_or0;
  assign u_dadda_cla8_fa21_and1 = u_dadda_cla8_fa21_xor0 & u_dadda_cla8_fa18_or0;
  assign u_dadda_cla8_fa21_or0 = u_dadda_cla8_fa21_and0 | u_dadda_cla8_fa21_and1;
  assign u_dadda_cla8_and_7_4 = a[7] & b[4];
  assign u_dadda_cla8_and_6_5 = a[6] & b[5];
  assign u_dadda_cla8_and_5_6 = a[5] & b[6];
  assign u_dadda_cla8_fa22_xor0 = u_dadda_cla8_and_7_4 ^ u_dadda_cla8_and_6_5;
  assign u_dadda_cla8_fa22_and0 = u_dadda_cla8_and_7_4 & u_dadda_cla8_and_6_5;
  assign u_dadda_cla8_fa22_xor1 = u_dadda_cla8_fa22_xor0 ^ u_dadda_cla8_and_5_6;
  assign u_dadda_cla8_fa22_and1 = u_dadda_cla8_fa22_xor0 & u_dadda_cla8_and_5_6;
  assign u_dadda_cla8_fa22_or0 = u_dadda_cla8_fa22_and0 | u_dadda_cla8_fa22_and1;
  assign u_dadda_cla8_and_7_5 = a[7] & b[5];
  assign u_dadda_cla8_fa23_xor0 = u_dadda_cla8_fa22_or0 ^ u_dadda_cla8_fa21_or0;
  assign u_dadda_cla8_fa23_and0 = u_dadda_cla8_fa22_or0 & u_dadda_cla8_fa21_or0;
  assign u_dadda_cla8_fa23_xor1 = u_dadda_cla8_fa23_xor0 ^ u_dadda_cla8_and_7_5;
  assign u_dadda_cla8_fa23_and1 = u_dadda_cla8_fa23_xor0 & u_dadda_cla8_and_7_5;
  assign u_dadda_cla8_fa23_or0 = u_dadda_cla8_fa23_and0 | u_dadda_cla8_fa23_and1;
  assign u_dadda_cla8_and_2_0 = a[2] & b[0];
  assign u_dadda_cla8_and_1_1 = a[1] & b[1];
  assign u_dadda_cla8_ha6_xor0 = u_dadda_cla8_and_2_0 ^ u_dadda_cla8_and_1_1;
  assign u_dadda_cla8_ha6_and0 = u_dadda_cla8_and_2_0 & u_dadda_cla8_and_1_1;
  assign u_dadda_cla8_and_1_2 = a[1] & b[2];
  assign u_dadda_cla8_and_0_3 = a[0] & b[3];
  assign u_dadda_cla8_fa24_xor0 = u_dadda_cla8_ha6_and0 ^ u_dadda_cla8_and_1_2;
  assign u_dadda_cla8_fa24_and0 = u_dadda_cla8_ha6_and0 & u_dadda_cla8_and_1_2;
  assign u_dadda_cla8_fa24_xor1 = u_dadda_cla8_fa24_xor0 ^ u_dadda_cla8_and_0_3;
  assign u_dadda_cla8_fa24_and1 = u_dadda_cla8_fa24_xor0 & u_dadda_cla8_and_0_3;
  assign u_dadda_cla8_fa24_or0 = u_dadda_cla8_fa24_and0 | u_dadda_cla8_fa24_and1;
  assign u_dadda_cla8_and_0_4 = a[0] & b[4];
  assign u_dadda_cla8_fa25_xor0 = u_dadda_cla8_fa24_or0 ^ u_dadda_cla8_and_0_4;
  assign u_dadda_cla8_fa25_and0 = u_dadda_cla8_fa24_or0 & u_dadda_cla8_and_0_4;
  assign u_dadda_cla8_fa25_xor1 = u_dadda_cla8_fa25_xor0 ^ u_dadda_cla8_fa3_xor1;
  assign u_dadda_cla8_fa25_and1 = u_dadda_cla8_fa25_xor0 & u_dadda_cla8_fa3_xor1;
  assign u_dadda_cla8_fa25_or0 = u_dadda_cla8_fa25_and0 | u_dadda_cla8_fa25_and1;
  assign u_dadda_cla8_fa26_xor0 = u_dadda_cla8_fa25_or0 ^ u_dadda_cla8_fa4_xor1;
  assign u_dadda_cla8_fa26_and0 = u_dadda_cla8_fa25_or0 & u_dadda_cla8_fa4_xor1;
  assign u_dadda_cla8_fa26_xor1 = u_dadda_cla8_fa26_xor0 ^ u_dadda_cla8_fa5_xor1;
  assign u_dadda_cla8_fa26_and1 = u_dadda_cla8_fa26_xor0 & u_dadda_cla8_fa5_xor1;
  assign u_dadda_cla8_fa26_or0 = u_dadda_cla8_fa26_and0 | u_dadda_cla8_fa26_and1;
  assign u_dadda_cla8_fa27_xor0 = u_dadda_cla8_fa26_or0 ^ u_dadda_cla8_fa6_xor1;
  assign u_dadda_cla8_fa27_and0 = u_dadda_cla8_fa26_or0 & u_dadda_cla8_fa6_xor1;
  assign u_dadda_cla8_fa27_xor1 = u_dadda_cla8_fa27_xor0 ^ u_dadda_cla8_fa7_xor1;
  assign u_dadda_cla8_fa27_and1 = u_dadda_cla8_fa27_xor0 & u_dadda_cla8_fa7_xor1;
  assign u_dadda_cla8_fa27_or0 = u_dadda_cla8_fa27_and0 | u_dadda_cla8_fa27_and1;
  assign u_dadda_cla8_fa28_xor0 = u_dadda_cla8_fa27_or0 ^ u_dadda_cla8_fa9_xor1;
  assign u_dadda_cla8_fa28_and0 = u_dadda_cla8_fa27_or0 & u_dadda_cla8_fa9_xor1;
  assign u_dadda_cla8_fa28_xor1 = u_dadda_cla8_fa28_xor0 ^ u_dadda_cla8_fa10_xor1;
  assign u_dadda_cla8_fa28_and1 = u_dadda_cla8_fa28_xor0 & u_dadda_cla8_fa10_xor1;
  assign u_dadda_cla8_fa28_or0 = u_dadda_cla8_fa28_and0 | u_dadda_cla8_fa28_and1;
  assign u_dadda_cla8_fa29_xor0 = u_dadda_cla8_fa28_or0 ^ u_dadda_cla8_fa12_xor1;
  assign u_dadda_cla8_fa29_and0 = u_dadda_cla8_fa28_or0 & u_dadda_cla8_fa12_xor1;
  assign u_dadda_cla8_fa29_xor1 = u_dadda_cla8_fa29_xor0 ^ u_dadda_cla8_fa13_xor1;
  assign u_dadda_cla8_fa29_and1 = u_dadda_cla8_fa29_xor0 & u_dadda_cla8_fa13_xor1;
  assign u_dadda_cla8_fa29_or0 = u_dadda_cla8_fa29_and0 | u_dadda_cla8_fa29_and1;
  assign u_dadda_cla8_fa30_xor0 = u_dadda_cla8_fa29_or0 ^ u_dadda_cla8_fa15_xor1;
  assign u_dadda_cla8_fa30_and0 = u_dadda_cla8_fa29_or0 & u_dadda_cla8_fa15_xor1;
  assign u_dadda_cla8_fa30_xor1 = u_dadda_cla8_fa30_xor0 ^ u_dadda_cla8_fa16_xor1;
  assign u_dadda_cla8_fa30_and1 = u_dadda_cla8_fa30_xor0 & u_dadda_cla8_fa16_xor1;
  assign u_dadda_cla8_fa30_or0 = u_dadda_cla8_fa30_and0 | u_dadda_cla8_fa30_and1;
  assign u_dadda_cla8_fa31_xor0 = u_dadda_cla8_fa30_or0 ^ u_dadda_cla8_fa18_xor1;
  assign u_dadda_cla8_fa31_and0 = u_dadda_cla8_fa30_or0 & u_dadda_cla8_fa18_xor1;
  assign u_dadda_cla8_fa31_xor1 = u_dadda_cla8_fa31_xor0 ^ u_dadda_cla8_fa19_xor1;
  assign u_dadda_cla8_fa31_and1 = u_dadda_cla8_fa31_xor0 & u_dadda_cla8_fa19_xor1;
  assign u_dadda_cla8_fa31_or0 = u_dadda_cla8_fa31_and0 | u_dadda_cla8_fa31_and1;
  assign u_dadda_cla8_and_4_7 = a[4] & b[7];
  assign u_dadda_cla8_fa32_xor0 = u_dadda_cla8_fa31_or0 ^ u_dadda_cla8_and_4_7;
  assign u_dadda_cla8_fa32_and0 = u_dadda_cla8_fa31_or0 & u_dadda_cla8_and_4_7;
  assign u_dadda_cla8_fa32_xor1 = u_dadda_cla8_fa32_xor0 ^ u_dadda_cla8_fa21_xor1;
  assign u_dadda_cla8_fa32_and1 = u_dadda_cla8_fa32_xor0 & u_dadda_cla8_fa21_xor1;
  assign u_dadda_cla8_fa32_or0 = u_dadda_cla8_fa32_and0 | u_dadda_cla8_fa32_and1;
  assign u_dadda_cla8_and_6_6 = a[6] & b[6];
  assign u_dadda_cla8_and_5_7 = a[5] & b[7];
  assign u_dadda_cla8_fa33_xor0 = u_dadda_cla8_fa32_or0 ^ u_dadda_cla8_and_6_6;
  assign u_dadda_cla8_fa33_and0 = u_dadda_cla8_fa32_or0 & u_dadda_cla8_and_6_6;
  assign u_dadda_cla8_fa33_xor1 = u_dadda_cla8_fa33_xor0 ^ u_dadda_cla8_and_5_7;
  assign u_dadda_cla8_fa33_and1 = u_dadda_cla8_fa33_xor0 & u_dadda_cla8_and_5_7;
  assign u_dadda_cla8_fa33_or0 = u_dadda_cla8_fa33_and0 | u_dadda_cla8_fa33_and1;
  assign u_dadda_cla8_and_7_6 = a[7] & b[6];
  assign u_dadda_cla8_fa34_xor0 = u_dadda_cla8_fa33_or0 ^ u_dadda_cla8_fa23_or0;
  assign u_dadda_cla8_fa34_and0 = u_dadda_cla8_fa33_or0 & u_dadda_cla8_fa23_or0;
  assign u_dadda_cla8_fa34_xor1 = u_dadda_cla8_fa34_xor0 ^ u_dadda_cla8_and_7_6;
  assign u_dadda_cla8_fa34_and1 = u_dadda_cla8_fa34_xor0 & u_dadda_cla8_and_7_6;
  assign u_dadda_cla8_fa34_or0 = u_dadda_cla8_fa34_and0 | u_dadda_cla8_fa34_and1;
  assign u_dadda_cla8_and_0_0 = a[0] & b[0];
  assign u_dadda_cla8_and_1_0 = a[1] & b[0];
  assign u_dadda_cla8_and_0_2 = a[0] & b[2];
  assign u_dadda_cla8_and_6_7 = a[6] & b[7];
  assign u_dadda_cla8_and_0_1 = a[0] & b[1];
  assign u_dadda_cla8_and_7_7 = a[7] & b[7];
  assign u_dadda_cla8_u_cla14_pg_logic0_or0 = u_dadda_cla8_and_1_0 | u_dadda_cla8_and_0_1;
  assign u_dadda_cla8_u_cla14_pg_logic0_and0 = u_dadda_cla8_and_1_0 & u_dadda_cla8_and_0_1;
  assign u_dadda_cla8_u_cla14_pg_logic0_xor0 = u_dadda_cla8_and_1_0 ^ u_dadda_cla8_and_0_1;
  assign u_dadda_cla8_u_cla14_pg_logic1_or0 = u_dadda_cla8_and_0_2 | u_dadda_cla8_ha6_xor0;
  assign u_dadda_cla8_u_cla14_pg_logic1_and0 = u_dadda_cla8_and_0_2 & u_dadda_cla8_ha6_xor0;
  assign u_dadda_cla8_u_cla14_pg_logic1_xor0 = u_dadda_cla8_and_0_2 ^ u_dadda_cla8_ha6_xor0;
  assign u_dadda_cla8_u_cla14_xor1 = u_dadda_cla8_u_cla14_pg_logic1_xor0 ^ u_dadda_cla8_u_cla14_pg_logic0_and0;
  assign u_dadda_cla8_u_cla14_and0 = u_dadda_cla8_u_cla14_pg_logic0_and0 & u_dadda_cla8_u_cla14_pg_logic1_or0;
  assign u_dadda_cla8_u_cla14_or0 = u_dadda_cla8_u_cla14_pg_logic1_and0 | u_dadda_cla8_u_cla14_and0;
  assign u_dadda_cla8_u_cla14_pg_logic2_or0 = u_dadda_cla8_ha3_xor0 | u_dadda_cla8_fa24_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic2_and0 = u_dadda_cla8_ha3_xor0 & u_dadda_cla8_fa24_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic2_xor0 = u_dadda_cla8_ha3_xor0 ^ u_dadda_cla8_fa24_xor1;
  assign u_dadda_cla8_u_cla14_xor2 = u_dadda_cla8_u_cla14_pg_logic2_xor0 ^ u_dadda_cla8_u_cla14_or0;
  assign u_dadda_cla8_u_cla14_and1 = u_dadda_cla8_u_cla14_pg_logic2_or0 & u_dadda_cla8_u_cla14_pg_logic0_or0;
  assign u_dadda_cla8_u_cla14_and2 = u_dadda_cla8_u_cla14_pg_logic0_and0 & u_dadda_cla8_u_cla14_pg_logic2_or0;
  assign u_dadda_cla8_u_cla14_and3 = u_dadda_cla8_u_cla14_and2 & u_dadda_cla8_u_cla14_pg_logic1_or0;
  assign u_dadda_cla8_u_cla14_and4 = u_dadda_cla8_u_cla14_pg_logic1_and0 & u_dadda_cla8_u_cla14_pg_logic2_or0;
  assign u_dadda_cla8_u_cla14_or1 = u_dadda_cla8_u_cla14_and3 | u_dadda_cla8_u_cla14_and4;
  assign u_dadda_cla8_u_cla14_or2 = u_dadda_cla8_u_cla14_pg_logic2_and0 | u_dadda_cla8_u_cla14_or1;
  assign u_dadda_cla8_u_cla14_pg_logic3_or0 = u_dadda_cla8_ha4_xor0 | u_dadda_cla8_fa25_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic3_and0 = u_dadda_cla8_ha4_xor0 & u_dadda_cla8_fa25_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic3_xor0 = u_dadda_cla8_ha4_xor0 ^ u_dadda_cla8_fa25_xor1;
  assign u_dadda_cla8_u_cla14_xor3 = u_dadda_cla8_u_cla14_pg_logic3_xor0 ^ u_dadda_cla8_u_cla14_or2;
  assign u_dadda_cla8_u_cla14_and5 = u_dadda_cla8_u_cla14_pg_logic3_or0 & u_dadda_cla8_u_cla14_pg_logic1_or0;
  assign u_dadda_cla8_u_cla14_and6 = u_dadda_cla8_u_cla14_pg_logic0_and0 & u_dadda_cla8_u_cla14_pg_logic2_or0;
  assign u_dadda_cla8_u_cla14_and7 = u_dadda_cla8_u_cla14_pg_logic3_or0 & u_dadda_cla8_u_cla14_pg_logic1_or0;
  assign u_dadda_cla8_u_cla14_and8 = u_dadda_cla8_u_cla14_and6 & u_dadda_cla8_u_cla14_and7;
  assign u_dadda_cla8_u_cla14_and9 = u_dadda_cla8_u_cla14_pg_logic1_and0 & u_dadda_cla8_u_cla14_pg_logic3_or0;
  assign u_dadda_cla8_u_cla14_and10 = u_dadda_cla8_u_cla14_and9 & u_dadda_cla8_u_cla14_pg_logic2_or0;
  assign u_dadda_cla8_u_cla14_and11 = u_dadda_cla8_u_cla14_pg_logic2_and0 & u_dadda_cla8_u_cla14_pg_logic3_or0;
  assign u_dadda_cla8_u_cla14_or3 = u_dadda_cla8_u_cla14_and8 | u_dadda_cla8_u_cla14_and11;
  assign u_dadda_cla8_u_cla14_or4 = u_dadda_cla8_u_cla14_and10 | u_dadda_cla8_u_cla14_or3;
  assign u_dadda_cla8_u_cla14_or5 = u_dadda_cla8_u_cla14_pg_logic3_and0 | u_dadda_cla8_u_cla14_or4;
  assign u_dadda_cla8_u_cla14_pg_logic4_or0 = u_dadda_cla8_ha5_xor0 | u_dadda_cla8_fa26_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic4_and0 = u_dadda_cla8_ha5_xor0 & u_dadda_cla8_fa26_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic4_xor0 = u_dadda_cla8_ha5_xor0 ^ u_dadda_cla8_fa26_xor1;
  assign u_dadda_cla8_u_cla14_xor4 = u_dadda_cla8_u_cla14_pg_logic4_xor0 ^ u_dadda_cla8_u_cla14_or5;
  assign u_dadda_cla8_u_cla14_and12 = u_dadda_cla8_u_cla14_or5 & u_dadda_cla8_u_cla14_pg_logic4_or0;
  assign u_dadda_cla8_u_cla14_or6 = u_dadda_cla8_u_cla14_pg_logic4_and0 | u_dadda_cla8_u_cla14_and12;
  assign u_dadda_cla8_u_cla14_pg_logic5_or0 = u_dadda_cla8_fa8_xor1 | u_dadda_cla8_fa27_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic5_and0 = u_dadda_cla8_fa8_xor1 & u_dadda_cla8_fa27_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic5_xor0 = u_dadda_cla8_fa8_xor1 ^ u_dadda_cla8_fa27_xor1;
  assign u_dadda_cla8_u_cla14_xor5 = u_dadda_cla8_u_cla14_pg_logic5_xor0 ^ u_dadda_cla8_u_cla14_or6;
  assign u_dadda_cla8_u_cla14_and13 = u_dadda_cla8_u_cla14_or5 & u_dadda_cla8_u_cla14_pg_logic5_or0;
  assign u_dadda_cla8_u_cla14_and14 = u_dadda_cla8_u_cla14_and13 & u_dadda_cla8_u_cla14_pg_logic4_or0;
  assign u_dadda_cla8_u_cla14_and15 = u_dadda_cla8_u_cla14_pg_logic4_and0 & u_dadda_cla8_u_cla14_pg_logic5_or0;
  assign u_dadda_cla8_u_cla14_or7 = u_dadda_cla8_u_cla14_and14 | u_dadda_cla8_u_cla14_and15;
  assign u_dadda_cla8_u_cla14_or8 = u_dadda_cla8_u_cla14_pg_logic5_and0 | u_dadda_cla8_u_cla14_or7;
  assign u_dadda_cla8_u_cla14_pg_logic6_or0 = u_dadda_cla8_fa11_xor1 | u_dadda_cla8_fa28_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic6_and0 = u_dadda_cla8_fa11_xor1 & u_dadda_cla8_fa28_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic6_xor0 = u_dadda_cla8_fa11_xor1 ^ u_dadda_cla8_fa28_xor1;
  assign u_dadda_cla8_u_cla14_xor6 = u_dadda_cla8_u_cla14_pg_logic6_xor0 ^ u_dadda_cla8_u_cla14_or8;
  assign u_dadda_cla8_u_cla14_and16 = u_dadda_cla8_u_cla14_or5 & u_dadda_cla8_u_cla14_pg_logic5_or0;
  assign u_dadda_cla8_u_cla14_and17 = u_dadda_cla8_u_cla14_pg_logic6_or0 & u_dadda_cla8_u_cla14_pg_logic4_or0;
  assign u_dadda_cla8_u_cla14_and18 = u_dadda_cla8_u_cla14_and16 & u_dadda_cla8_u_cla14_and17;
  assign u_dadda_cla8_u_cla14_and19 = u_dadda_cla8_u_cla14_pg_logic4_and0 & u_dadda_cla8_u_cla14_pg_logic6_or0;
  assign u_dadda_cla8_u_cla14_and20 = u_dadda_cla8_u_cla14_and19 & u_dadda_cla8_u_cla14_pg_logic5_or0;
  assign u_dadda_cla8_u_cla14_and21 = u_dadda_cla8_u_cla14_pg_logic5_and0 & u_dadda_cla8_u_cla14_pg_logic6_or0;
  assign u_dadda_cla8_u_cla14_or9 = u_dadda_cla8_u_cla14_and18 | u_dadda_cla8_u_cla14_and20;
  assign u_dadda_cla8_u_cla14_or10 = u_dadda_cla8_u_cla14_or9 | u_dadda_cla8_u_cla14_and21;
  assign u_dadda_cla8_u_cla14_or11 = u_dadda_cla8_u_cla14_pg_logic6_and0 | u_dadda_cla8_u_cla14_or10;
  assign u_dadda_cla8_u_cla14_pg_logic7_or0 = u_dadda_cla8_fa14_xor1 | u_dadda_cla8_fa29_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic7_and0 = u_dadda_cla8_fa14_xor1 & u_dadda_cla8_fa29_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic7_xor0 = u_dadda_cla8_fa14_xor1 ^ u_dadda_cla8_fa29_xor1;
  assign u_dadda_cla8_u_cla14_xor7 = u_dadda_cla8_u_cla14_pg_logic7_xor0 ^ u_dadda_cla8_u_cla14_or11;
  assign u_dadda_cla8_u_cla14_and22 = u_dadda_cla8_u_cla14_or5 & u_dadda_cla8_u_cla14_pg_logic6_or0;
  assign u_dadda_cla8_u_cla14_and23 = u_dadda_cla8_u_cla14_pg_logic7_or0 & u_dadda_cla8_u_cla14_pg_logic5_or0;
  assign u_dadda_cla8_u_cla14_and24 = u_dadda_cla8_u_cla14_and22 & u_dadda_cla8_u_cla14_and23;
  assign u_dadda_cla8_u_cla14_and25 = u_dadda_cla8_u_cla14_and24 & u_dadda_cla8_u_cla14_pg_logic4_or0;
  assign u_dadda_cla8_u_cla14_and26 = u_dadda_cla8_u_cla14_pg_logic4_and0 & u_dadda_cla8_u_cla14_pg_logic6_or0;
  assign u_dadda_cla8_u_cla14_and27 = u_dadda_cla8_u_cla14_pg_logic7_or0 & u_dadda_cla8_u_cla14_pg_logic5_or0;
  assign u_dadda_cla8_u_cla14_and28 = u_dadda_cla8_u_cla14_and26 & u_dadda_cla8_u_cla14_and27;
  assign u_dadda_cla8_u_cla14_and29 = u_dadda_cla8_u_cla14_pg_logic5_and0 & u_dadda_cla8_u_cla14_pg_logic7_or0;
  assign u_dadda_cla8_u_cla14_and30 = u_dadda_cla8_u_cla14_and29 & u_dadda_cla8_u_cla14_pg_logic6_or0;
  assign u_dadda_cla8_u_cla14_and31 = u_dadda_cla8_u_cla14_pg_logic6_and0 & u_dadda_cla8_u_cla14_pg_logic7_or0;
  assign u_dadda_cla8_u_cla14_or12 = u_dadda_cla8_u_cla14_and25 | u_dadda_cla8_u_cla14_and30;
  assign u_dadda_cla8_u_cla14_or13 = u_dadda_cla8_u_cla14_and28 | u_dadda_cla8_u_cla14_and31;
  assign u_dadda_cla8_u_cla14_or14 = u_dadda_cla8_u_cla14_or12 | u_dadda_cla8_u_cla14_or13;
  assign u_dadda_cla8_u_cla14_or15 = u_dadda_cla8_u_cla14_pg_logic7_and0 | u_dadda_cla8_u_cla14_or14;
  assign u_dadda_cla8_u_cla14_pg_logic8_or0 = u_dadda_cla8_fa17_xor1 | u_dadda_cla8_fa30_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic8_and0 = u_dadda_cla8_fa17_xor1 & u_dadda_cla8_fa30_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic8_xor0 = u_dadda_cla8_fa17_xor1 ^ u_dadda_cla8_fa30_xor1;
  assign u_dadda_cla8_u_cla14_xor8 = u_dadda_cla8_u_cla14_pg_logic8_xor0 ^ u_dadda_cla8_u_cla14_or15;
  assign u_dadda_cla8_u_cla14_and32 = u_dadda_cla8_u_cla14_or15 & u_dadda_cla8_u_cla14_pg_logic8_or0;
  assign u_dadda_cla8_u_cla14_or16 = u_dadda_cla8_u_cla14_pg_logic8_and0 | u_dadda_cla8_u_cla14_and32;
  assign u_dadda_cla8_u_cla14_pg_logic9_or0 = u_dadda_cla8_fa20_xor1 | u_dadda_cla8_fa31_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic9_and0 = u_dadda_cla8_fa20_xor1 & u_dadda_cla8_fa31_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic9_xor0 = u_dadda_cla8_fa20_xor1 ^ u_dadda_cla8_fa31_xor1;
  assign u_dadda_cla8_u_cla14_xor9 = u_dadda_cla8_u_cla14_pg_logic9_xor0 ^ u_dadda_cla8_u_cla14_or16;
  assign u_dadda_cla8_u_cla14_and33 = u_dadda_cla8_u_cla14_or15 & u_dadda_cla8_u_cla14_pg_logic9_or0;
  assign u_dadda_cla8_u_cla14_and34 = u_dadda_cla8_u_cla14_and33 & u_dadda_cla8_u_cla14_pg_logic8_or0;
  assign u_dadda_cla8_u_cla14_and35 = u_dadda_cla8_u_cla14_pg_logic8_and0 & u_dadda_cla8_u_cla14_pg_logic9_or0;
  assign u_dadda_cla8_u_cla14_or17 = u_dadda_cla8_u_cla14_and34 | u_dadda_cla8_u_cla14_and35;
  assign u_dadda_cla8_u_cla14_or18 = u_dadda_cla8_u_cla14_pg_logic9_and0 | u_dadda_cla8_u_cla14_or17;
  assign u_dadda_cla8_u_cla14_pg_logic10_or0 = u_dadda_cla8_fa22_xor1 | u_dadda_cla8_fa32_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic10_and0 = u_dadda_cla8_fa22_xor1 & u_dadda_cla8_fa32_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic10_xor0 = u_dadda_cla8_fa22_xor1 ^ u_dadda_cla8_fa32_xor1;
  assign u_dadda_cla8_u_cla14_xor10 = u_dadda_cla8_u_cla14_pg_logic10_xor0 ^ u_dadda_cla8_u_cla14_or18;
  assign u_dadda_cla8_u_cla14_and36 = u_dadda_cla8_u_cla14_or15 & u_dadda_cla8_u_cla14_pg_logic9_or0;
  assign u_dadda_cla8_u_cla14_and37 = u_dadda_cla8_u_cla14_pg_logic10_or0 & u_dadda_cla8_u_cla14_pg_logic8_or0;
  assign u_dadda_cla8_u_cla14_and38 = u_dadda_cla8_u_cla14_and36 & u_dadda_cla8_u_cla14_and37;
  assign u_dadda_cla8_u_cla14_and39 = u_dadda_cla8_u_cla14_pg_logic8_and0 & u_dadda_cla8_u_cla14_pg_logic10_or0;
  assign u_dadda_cla8_u_cla14_and40 = u_dadda_cla8_u_cla14_and39 & u_dadda_cla8_u_cla14_pg_logic9_or0;
  assign u_dadda_cla8_u_cla14_and41 = u_dadda_cla8_u_cla14_pg_logic9_and0 & u_dadda_cla8_u_cla14_pg_logic10_or0;
  assign u_dadda_cla8_u_cla14_or19 = u_dadda_cla8_u_cla14_and38 | u_dadda_cla8_u_cla14_and40;
  assign u_dadda_cla8_u_cla14_or20 = u_dadda_cla8_u_cla14_or19 | u_dadda_cla8_u_cla14_and41;
  assign u_dadda_cla8_u_cla14_or21 = u_dadda_cla8_u_cla14_pg_logic10_and0 | u_dadda_cla8_u_cla14_or20;
  assign u_dadda_cla8_u_cla14_pg_logic11_or0 = u_dadda_cla8_fa23_xor1 | u_dadda_cla8_fa33_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic11_and0 = u_dadda_cla8_fa23_xor1 & u_dadda_cla8_fa33_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic11_xor0 = u_dadda_cla8_fa23_xor1 ^ u_dadda_cla8_fa33_xor1;
  assign u_dadda_cla8_u_cla14_xor11 = u_dadda_cla8_u_cla14_pg_logic11_xor0 ^ u_dadda_cla8_u_cla14_or21;
  assign u_dadda_cla8_u_cla14_and42 = u_dadda_cla8_u_cla14_or15 & u_dadda_cla8_u_cla14_pg_logic10_or0;
  assign u_dadda_cla8_u_cla14_and43 = u_dadda_cla8_u_cla14_pg_logic11_or0 & u_dadda_cla8_u_cla14_pg_logic9_or0;
  assign u_dadda_cla8_u_cla14_and44 = u_dadda_cla8_u_cla14_and42 & u_dadda_cla8_u_cla14_and43;
  assign u_dadda_cla8_u_cla14_and45 = u_dadda_cla8_u_cla14_and44 & u_dadda_cla8_u_cla14_pg_logic8_or0;
  assign u_dadda_cla8_u_cla14_and46 = u_dadda_cla8_u_cla14_pg_logic8_and0 & u_dadda_cla8_u_cla14_pg_logic10_or0;
  assign u_dadda_cla8_u_cla14_and47 = u_dadda_cla8_u_cla14_pg_logic11_or0 & u_dadda_cla8_u_cla14_pg_logic9_or0;
  assign u_dadda_cla8_u_cla14_and48 = u_dadda_cla8_u_cla14_and46 & u_dadda_cla8_u_cla14_and47;
  assign u_dadda_cla8_u_cla14_and49 = u_dadda_cla8_u_cla14_pg_logic9_and0 & u_dadda_cla8_u_cla14_pg_logic11_or0;
  assign u_dadda_cla8_u_cla14_and50 = u_dadda_cla8_u_cla14_and49 & u_dadda_cla8_u_cla14_pg_logic10_or0;
  assign u_dadda_cla8_u_cla14_and51 = u_dadda_cla8_u_cla14_pg_logic10_and0 & u_dadda_cla8_u_cla14_pg_logic11_or0;
  assign u_dadda_cla8_u_cla14_or22 = u_dadda_cla8_u_cla14_and45 | u_dadda_cla8_u_cla14_and50;
  assign u_dadda_cla8_u_cla14_or23 = u_dadda_cla8_u_cla14_and48 | u_dadda_cla8_u_cla14_and51;
  assign u_dadda_cla8_u_cla14_or24 = u_dadda_cla8_u_cla14_or22 | u_dadda_cla8_u_cla14_or23;
  assign u_dadda_cla8_u_cla14_or25 = u_dadda_cla8_u_cla14_pg_logic11_and0 | u_dadda_cla8_u_cla14_or24;
  assign u_dadda_cla8_u_cla14_pg_logic12_or0 = u_dadda_cla8_and_6_7 | u_dadda_cla8_fa34_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic12_and0 = u_dadda_cla8_and_6_7 & u_dadda_cla8_fa34_xor1;
  assign u_dadda_cla8_u_cla14_pg_logic12_xor0 = u_dadda_cla8_and_6_7 ^ u_dadda_cla8_fa34_xor1;
  assign u_dadda_cla8_u_cla14_xor12 = u_dadda_cla8_u_cla14_pg_logic12_xor0 ^ u_dadda_cla8_u_cla14_or25;
  assign u_dadda_cla8_u_cla14_and52 = u_dadda_cla8_u_cla14_or25 & u_dadda_cla8_u_cla14_pg_logic12_or0;
  assign u_dadda_cla8_u_cla14_or26 = u_dadda_cla8_u_cla14_pg_logic12_and0 | u_dadda_cla8_u_cla14_and52;
  assign u_dadda_cla8_u_cla14_pg_logic13_or0 = u_dadda_cla8_fa34_or0 | u_dadda_cla8_and_7_7;
  assign u_dadda_cla8_u_cla14_pg_logic13_and0 = u_dadda_cla8_fa34_or0 & u_dadda_cla8_and_7_7;
  assign u_dadda_cla8_u_cla14_pg_logic13_xor0 = u_dadda_cla8_fa34_or0 ^ u_dadda_cla8_and_7_7;
  assign u_dadda_cla8_u_cla14_xor13 = u_dadda_cla8_u_cla14_pg_logic13_xor0 ^ u_dadda_cla8_u_cla14_or26;
  assign u_dadda_cla8_u_cla14_and53 = u_dadda_cla8_u_cla14_or25 & u_dadda_cla8_u_cla14_pg_logic13_or0;
  assign u_dadda_cla8_u_cla14_and54 = u_dadda_cla8_u_cla14_and53 & u_dadda_cla8_u_cla14_pg_logic12_or0;
  assign u_dadda_cla8_u_cla14_and55 = u_dadda_cla8_u_cla14_pg_logic12_and0 & u_dadda_cla8_u_cla14_pg_logic13_or0;
  assign u_dadda_cla8_u_cla14_or27 = u_dadda_cla8_u_cla14_and54 | u_dadda_cla8_u_cla14_and55;
  assign u_dadda_cla8_u_cla14_or28 = u_dadda_cla8_u_cla14_pg_logic13_and0 | u_dadda_cla8_u_cla14_or27;

  assign u_dadda_cla8_out[0] = u_dadda_cla8_and_0_0;
  assign u_dadda_cla8_out[1] = u_dadda_cla8_u_cla14_pg_logic0_xor0;
  assign u_dadda_cla8_out[2] = u_dadda_cla8_u_cla14_xor1;
  assign u_dadda_cla8_out[3] = u_dadda_cla8_u_cla14_xor2;
  assign u_dadda_cla8_out[4] = u_dadda_cla8_u_cla14_xor3;
  assign u_dadda_cla8_out[5] = u_dadda_cla8_u_cla14_xor4;
  assign u_dadda_cla8_out[6] = u_dadda_cla8_u_cla14_xor5;
  assign u_dadda_cla8_out[7] = u_dadda_cla8_u_cla14_xor6;
  assign u_dadda_cla8_out[8] = u_dadda_cla8_u_cla14_xor7;
  assign u_dadda_cla8_out[9] = u_dadda_cla8_u_cla14_xor8;
  assign u_dadda_cla8_out[10] = u_dadda_cla8_u_cla14_xor9;
  assign u_dadda_cla8_out[11] = u_dadda_cla8_u_cla14_xor10;
  assign u_dadda_cla8_out[12] = u_dadda_cla8_u_cla14_xor11;
  assign u_dadda_cla8_out[13] = u_dadda_cla8_u_cla14_xor12;
  assign u_dadda_cla8_out[14] = u_dadda_cla8_u_cla14_xor13;
  assign u_dadda_cla8_out[15] = u_dadda_cla8_u_cla14_or28;
endmodule