module u_cla12(input [11:0] a, input [11:0] b, output [12:0] u_cla12_out);
  wire u_cla12_pg_logic0_or0;
  wire u_cla12_pg_logic0_and0;
  wire u_cla12_pg_logic0_xor0;
  wire u_cla12_pg_logic1_or0;
  wire u_cla12_pg_logic1_and0;
  wire u_cla12_pg_logic1_xor0;
  wire u_cla12_xor1;
  wire u_cla12_and0;
  wire u_cla12_or0;
  wire u_cla12_pg_logic2_or0;
  wire u_cla12_pg_logic2_and0;
  wire u_cla12_pg_logic2_xor0;
  wire u_cla12_xor2;
  wire u_cla12_and1;
  wire u_cla12_and2;
  wire u_cla12_and3;
  wire u_cla12_and4;
  wire u_cla12_or1;
  wire u_cla12_or2;
  wire u_cla12_pg_logic3_or0;
  wire u_cla12_pg_logic3_and0;
  wire u_cla12_pg_logic3_xor0;
  wire u_cla12_xor3;
  wire u_cla12_and5;
  wire u_cla12_and6;
  wire u_cla12_and7;
  wire u_cla12_and8;
  wire u_cla12_and9;
  wire u_cla12_and10;
  wire u_cla12_and11;
  wire u_cla12_or3;
  wire u_cla12_or4;
  wire u_cla12_or5;
  wire u_cla12_pg_logic4_or0;
  wire u_cla12_pg_logic4_and0;
  wire u_cla12_pg_logic4_xor0;
  wire u_cla12_xor4;
  wire u_cla12_and12;
  wire u_cla12_or6;
  wire u_cla12_pg_logic5_or0;
  wire u_cla12_pg_logic5_and0;
  wire u_cla12_pg_logic5_xor0;
  wire u_cla12_xor5;
  wire u_cla12_and13;
  wire u_cla12_and14;
  wire u_cla12_and15;
  wire u_cla12_or7;
  wire u_cla12_or8;
  wire u_cla12_pg_logic6_or0;
  wire u_cla12_pg_logic6_and0;
  wire u_cla12_pg_logic6_xor0;
  wire u_cla12_xor6;
  wire u_cla12_and16;
  wire u_cla12_and17;
  wire u_cla12_and18;
  wire u_cla12_and19;
  wire u_cla12_and20;
  wire u_cla12_and21;
  wire u_cla12_or9;
  wire u_cla12_or10;
  wire u_cla12_or11;
  wire u_cla12_pg_logic7_or0;
  wire u_cla12_pg_logic7_and0;
  wire u_cla12_pg_logic7_xor0;
  wire u_cla12_xor7;
  wire u_cla12_and22;
  wire u_cla12_and23;
  wire u_cla12_and24;
  wire u_cla12_and25;
  wire u_cla12_and26;
  wire u_cla12_and27;
  wire u_cla12_and28;
  wire u_cla12_and29;
  wire u_cla12_and30;
  wire u_cla12_and31;
  wire u_cla12_or12;
  wire u_cla12_or13;
  wire u_cla12_or14;
  wire u_cla12_or15;
  wire u_cla12_pg_logic8_or0;
  wire u_cla12_pg_logic8_and0;
  wire u_cla12_pg_logic8_xor0;
  wire u_cla12_xor8;
  wire u_cla12_and32;
  wire u_cla12_or16;
  wire u_cla12_pg_logic9_or0;
  wire u_cla12_pg_logic9_and0;
  wire u_cla12_pg_logic9_xor0;
  wire u_cla12_xor9;
  wire u_cla12_and33;
  wire u_cla12_and34;
  wire u_cla12_and35;
  wire u_cla12_or17;
  wire u_cla12_or18;
  wire u_cla12_pg_logic10_or0;
  wire u_cla12_pg_logic10_and0;
  wire u_cla12_pg_logic10_xor0;
  wire u_cla12_xor10;
  wire u_cla12_and36;
  wire u_cla12_and37;
  wire u_cla12_and38;
  wire u_cla12_and39;
  wire u_cla12_and40;
  wire u_cla12_and41;
  wire u_cla12_or19;
  wire u_cla12_or20;
  wire u_cla12_or21;
  wire u_cla12_pg_logic11_or0;
  wire u_cla12_pg_logic11_and0;
  wire u_cla12_pg_logic11_xor0;
  wire u_cla12_xor11;
  wire u_cla12_and42;
  wire u_cla12_and43;
  wire u_cla12_and44;
  wire u_cla12_and45;
  wire u_cla12_and46;
  wire u_cla12_and47;
  wire u_cla12_and48;
  wire u_cla12_and49;
  wire u_cla12_and50;
  wire u_cla12_and51;
  wire u_cla12_or22;
  wire u_cla12_or23;
  wire u_cla12_or24;
  wire u_cla12_or25;

  assign u_cla12_pg_logic0_or0 = a[0] | b[0];
  assign u_cla12_pg_logic0_and0 = a[0] & b[0];
  assign u_cla12_pg_logic0_xor0 = a[0] ^ b[0];
  assign u_cla12_pg_logic1_or0 = a[1] | b[1];
  assign u_cla12_pg_logic1_and0 = a[1] & b[1];
  assign u_cla12_pg_logic1_xor0 = a[1] ^ b[1];
  assign u_cla12_xor1 = u_cla12_pg_logic1_xor0 ^ u_cla12_pg_logic0_and0;
  assign u_cla12_and0 = u_cla12_pg_logic0_and0 & u_cla12_pg_logic1_or0;
  assign u_cla12_or0 = u_cla12_pg_logic1_and0 | u_cla12_and0;
  assign u_cla12_pg_logic2_or0 = a[2] | b[2];
  assign u_cla12_pg_logic2_and0 = a[2] & b[2];
  assign u_cla12_pg_logic2_xor0 = a[2] ^ b[2];
  assign u_cla12_xor2 = u_cla12_pg_logic2_xor0 ^ u_cla12_or0;
  assign u_cla12_and1 = u_cla12_pg_logic2_or0 & u_cla12_pg_logic0_or0;
  assign u_cla12_and2 = u_cla12_pg_logic0_and0 & u_cla12_pg_logic2_or0;
  assign u_cla12_and3 = u_cla12_and2 & u_cla12_pg_logic1_or0;
  assign u_cla12_and4 = u_cla12_pg_logic1_and0 & u_cla12_pg_logic2_or0;
  assign u_cla12_or1 = u_cla12_and3 | u_cla12_and4;
  assign u_cla12_or2 = u_cla12_pg_logic2_and0 | u_cla12_or1;
  assign u_cla12_pg_logic3_or0 = a[3] | b[3];
  assign u_cla12_pg_logic3_and0 = a[3] & b[3];
  assign u_cla12_pg_logic3_xor0 = a[3] ^ b[3];
  assign u_cla12_xor3 = u_cla12_pg_logic3_xor0 ^ u_cla12_or2;
  assign u_cla12_and5 = u_cla12_pg_logic3_or0 & u_cla12_pg_logic1_or0;
  assign u_cla12_and6 = u_cla12_pg_logic0_and0 & u_cla12_pg_logic2_or0;
  assign u_cla12_and7 = u_cla12_pg_logic3_or0 & u_cla12_pg_logic1_or0;
  assign u_cla12_and8 = u_cla12_and6 & u_cla12_and7;
  assign u_cla12_and9 = u_cla12_pg_logic1_and0 & u_cla12_pg_logic3_or0;
  assign u_cla12_and10 = u_cla12_and9 & u_cla12_pg_logic2_or0;
  assign u_cla12_and11 = u_cla12_pg_logic2_and0 & u_cla12_pg_logic3_or0;
  assign u_cla12_or3 = u_cla12_and8 | u_cla12_and11;
  assign u_cla12_or4 = u_cla12_and10 | u_cla12_or3;
  assign u_cla12_or5 = u_cla12_pg_logic3_and0 | u_cla12_or4;
  assign u_cla12_pg_logic4_or0 = a[4] | b[4];
  assign u_cla12_pg_logic4_and0 = a[4] & b[4];
  assign u_cla12_pg_logic4_xor0 = a[4] ^ b[4];
  assign u_cla12_xor4 = u_cla12_pg_logic4_xor0 ^ u_cla12_or5;
  assign u_cla12_and12 = u_cla12_or5 & u_cla12_pg_logic4_or0;
  assign u_cla12_or6 = u_cla12_pg_logic4_and0 | u_cla12_and12;
  assign u_cla12_pg_logic5_or0 = a[5] | b[5];
  assign u_cla12_pg_logic5_and0 = a[5] & b[5];
  assign u_cla12_pg_logic5_xor0 = a[5] ^ b[5];
  assign u_cla12_xor5 = u_cla12_pg_logic5_xor0 ^ u_cla12_or6;
  assign u_cla12_and13 = u_cla12_or5 & u_cla12_pg_logic5_or0;
  assign u_cla12_and14 = u_cla12_and13 & u_cla12_pg_logic4_or0;
  assign u_cla12_and15 = u_cla12_pg_logic4_and0 & u_cla12_pg_logic5_or0;
  assign u_cla12_or7 = u_cla12_and14 | u_cla12_and15;
  assign u_cla12_or8 = u_cla12_pg_logic5_and0 | u_cla12_or7;
  assign u_cla12_pg_logic6_or0 = a[6] | b[6];
  assign u_cla12_pg_logic6_and0 = a[6] & b[6];
  assign u_cla12_pg_logic6_xor0 = a[6] ^ b[6];
  assign u_cla12_xor6 = u_cla12_pg_logic6_xor0 ^ u_cla12_or8;
  assign u_cla12_and16 = u_cla12_or5 & u_cla12_pg_logic5_or0;
  assign u_cla12_and17 = u_cla12_pg_logic6_or0 & u_cla12_pg_logic4_or0;
  assign u_cla12_and18 = u_cla12_and16 & u_cla12_and17;
  assign u_cla12_and19 = u_cla12_pg_logic4_and0 & u_cla12_pg_logic6_or0;
  assign u_cla12_and20 = u_cla12_and19 & u_cla12_pg_logic5_or0;
  assign u_cla12_and21 = u_cla12_pg_logic5_and0 & u_cla12_pg_logic6_or0;
  assign u_cla12_or9 = u_cla12_and18 | u_cla12_and20;
  assign u_cla12_or10 = u_cla12_or9 | u_cla12_and21;
  assign u_cla12_or11 = u_cla12_pg_logic6_and0 | u_cla12_or10;
  assign u_cla12_pg_logic7_or0 = a[7] | b[7];
  assign u_cla12_pg_logic7_and0 = a[7] & b[7];
  assign u_cla12_pg_logic7_xor0 = a[7] ^ b[7];
  assign u_cla12_xor7 = u_cla12_pg_logic7_xor0 ^ u_cla12_or11;
  assign u_cla12_and22 = u_cla12_or5 & u_cla12_pg_logic6_or0;
  assign u_cla12_and23 = u_cla12_pg_logic7_or0 & u_cla12_pg_logic5_or0;
  assign u_cla12_and24 = u_cla12_and22 & u_cla12_and23;
  assign u_cla12_and25 = u_cla12_and24 & u_cla12_pg_logic4_or0;
  assign u_cla12_and26 = u_cla12_pg_logic4_and0 & u_cla12_pg_logic6_or0;
  assign u_cla12_and27 = u_cla12_pg_logic7_or0 & u_cla12_pg_logic5_or0;
  assign u_cla12_and28 = u_cla12_and26 & u_cla12_and27;
  assign u_cla12_and29 = u_cla12_pg_logic5_and0 & u_cla12_pg_logic7_or0;
  assign u_cla12_and30 = u_cla12_and29 & u_cla12_pg_logic6_or0;
  assign u_cla12_and31 = u_cla12_pg_logic6_and0 & u_cla12_pg_logic7_or0;
  assign u_cla12_or12 = u_cla12_and25 | u_cla12_and30;
  assign u_cla12_or13 = u_cla12_and28 | u_cla12_and31;
  assign u_cla12_or14 = u_cla12_or12 | u_cla12_or13;
  assign u_cla12_or15 = u_cla12_pg_logic7_and0 | u_cla12_or14;
  assign u_cla12_pg_logic8_or0 = a[8] | b[8];
  assign u_cla12_pg_logic8_and0 = a[8] & b[8];
  assign u_cla12_pg_logic8_xor0 = a[8] ^ b[8];
  assign u_cla12_xor8 = u_cla12_pg_logic8_xor0 ^ u_cla12_or15;
  assign u_cla12_and32 = u_cla12_or15 & u_cla12_pg_logic8_or0;
  assign u_cla12_or16 = u_cla12_pg_logic8_and0 | u_cla12_and32;
  assign u_cla12_pg_logic9_or0 = a[9] | b[9];
  assign u_cla12_pg_logic9_and0 = a[9] & b[9];
  assign u_cla12_pg_logic9_xor0 = a[9] ^ b[9];
  assign u_cla12_xor9 = u_cla12_pg_logic9_xor0 ^ u_cla12_or16;
  assign u_cla12_and33 = u_cla12_or15 & u_cla12_pg_logic9_or0;
  assign u_cla12_and34 = u_cla12_and33 & u_cla12_pg_logic8_or0;
  assign u_cla12_and35 = u_cla12_pg_logic8_and0 & u_cla12_pg_logic9_or0;
  assign u_cla12_or17 = u_cla12_and34 | u_cla12_and35;
  assign u_cla12_or18 = u_cla12_pg_logic9_and0 | u_cla12_or17;
  assign u_cla12_pg_logic10_or0 = a[10] | b[10];
  assign u_cla12_pg_logic10_and0 = a[10] & b[10];
  assign u_cla12_pg_logic10_xor0 = a[10] ^ b[10];
  assign u_cla12_xor10 = u_cla12_pg_logic10_xor0 ^ u_cla12_or18;
  assign u_cla12_and36 = u_cla12_or15 & u_cla12_pg_logic9_or0;
  assign u_cla12_and37 = u_cla12_pg_logic10_or0 & u_cla12_pg_logic8_or0;
  assign u_cla12_and38 = u_cla12_and36 & u_cla12_and37;
  assign u_cla12_and39 = u_cla12_pg_logic8_and0 & u_cla12_pg_logic10_or0;
  assign u_cla12_and40 = u_cla12_and39 & u_cla12_pg_logic9_or0;
  assign u_cla12_and41 = u_cla12_pg_logic9_and0 & u_cla12_pg_logic10_or0;
  assign u_cla12_or19 = u_cla12_and38 | u_cla12_and40;
  assign u_cla12_or20 = u_cla12_or19 | u_cla12_and41;
  assign u_cla12_or21 = u_cla12_pg_logic10_and0 | u_cla12_or20;
  assign u_cla12_pg_logic11_or0 = a[11] | b[11];
  assign u_cla12_pg_logic11_and0 = a[11] & b[11];
  assign u_cla12_pg_logic11_xor0 = a[11] ^ b[11];
  assign u_cla12_xor11 = u_cla12_pg_logic11_xor0 ^ u_cla12_or21;
  assign u_cla12_and42 = u_cla12_or15 & u_cla12_pg_logic10_or0;
  assign u_cla12_and43 = u_cla12_pg_logic11_or0 & u_cla12_pg_logic9_or0;
  assign u_cla12_and44 = u_cla12_and42 & u_cla12_and43;
  assign u_cla12_and45 = u_cla12_and44 & u_cla12_pg_logic8_or0;
  assign u_cla12_and46 = u_cla12_pg_logic8_and0 & u_cla12_pg_logic10_or0;
  assign u_cla12_and47 = u_cla12_pg_logic11_or0 & u_cla12_pg_logic9_or0;
  assign u_cla12_and48 = u_cla12_and46 & u_cla12_and47;
  assign u_cla12_and49 = u_cla12_pg_logic9_and0 & u_cla12_pg_logic11_or0;
  assign u_cla12_and50 = u_cla12_and49 & u_cla12_pg_logic10_or0;
  assign u_cla12_and51 = u_cla12_pg_logic10_and0 & u_cla12_pg_logic11_or0;
  assign u_cla12_or22 = u_cla12_and45 | u_cla12_and50;
  assign u_cla12_or23 = u_cla12_and48 | u_cla12_and51;
  assign u_cla12_or24 = u_cla12_or22 | u_cla12_or23;
  assign u_cla12_or25 = u_cla12_pg_logic11_and0 | u_cla12_or24;

  assign u_cla12_out[0] = u_cla12_pg_logic0_xor0;
  assign u_cla12_out[1] = u_cla12_xor1;
  assign u_cla12_out[2] = u_cla12_xor2;
  assign u_cla12_out[3] = u_cla12_xor3;
  assign u_cla12_out[4] = u_cla12_xor4;
  assign u_cla12_out[5] = u_cla12_xor5;
  assign u_cla12_out[6] = u_cla12_xor6;
  assign u_cla12_out[7] = u_cla12_xor7;
  assign u_cla12_out[8] = u_cla12_xor8;
  assign u_cla12_out[9] = u_cla12_xor9;
  assign u_cla12_out[10] = u_cla12_xor10;
  assign u_cla12_out[11] = u_cla12_xor11;
  assign u_cla12_out[12] = u_cla12_or25;
endmodule