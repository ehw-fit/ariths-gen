module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module h_s_arrmul16(input [15:0] a, input [15:0] b, output [31:0] h_s_arrmul16_out);
  wire [0:0] h_s_arrmul16_and0_0;
  wire [0:0] h_s_arrmul16_and1_0;
  wire [0:0] h_s_arrmul16_and2_0;
  wire [0:0] h_s_arrmul16_and3_0;
  wire [0:0] h_s_arrmul16_and4_0;
  wire [0:0] h_s_arrmul16_and5_0;
  wire [0:0] h_s_arrmul16_and6_0;
  wire [0:0] h_s_arrmul16_and7_0;
  wire [0:0] h_s_arrmul16_and8_0;
  wire [0:0] h_s_arrmul16_and9_0;
  wire [0:0] h_s_arrmul16_and10_0;
  wire [0:0] h_s_arrmul16_and11_0;
  wire [0:0] h_s_arrmul16_and12_0;
  wire [0:0] h_s_arrmul16_and13_0;
  wire [0:0] h_s_arrmul16_and14_0;
  wire [0:0] h_s_arrmul16_nand15_0;
  wire [0:0] h_s_arrmul16_and0_1;
  wire [0:0] h_s_arrmul16_ha0_1_xor0;
  wire [0:0] h_s_arrmul16_ha0_1_and0;
  wire [0:0] h_s_arrmul16_and1_1;
  wire [0:0] h_s_arrmul16_fa1_1_xor1;
  wire [0:0] h_s_arrmul16_fa1_1_or0;
  wire [0:0] h_s_arrmul16_and2_1;
  wire [0:0] h_s_arrmul16_fa2_1_xor1;
  wire [0:0] h_s_arrmul16_fa2_1_or0;
  wire [0:0] h_s_arrmul16_and3_1;
  wire [0:0] h_s_arrmul16_fa3_1_xor1;
  wire [0:0] h_s_arrmul16_fa3_1_or0;
  wire [0:0] h_s_arrmul16_and4_1;
  wire [0:0] h_s_arrmul16_fa4_1_xor1;
  wire [0:0] h_s_arrmul16_fa4_1_or0;
  wire [0:0] h_s_arrmul16_and5_1;
  wire [0:0] h_s_arrmul16_fa5_1_xor1;
  wire [0:0] h_s_arrmul16_fa5_1_or0;
  wire [0:0] h_s_arrmul16_and6_1;
  wire [0:0] h_s_arrmul16_fa6_1_xor1;
  wire [0:0] h_s_arrmul16_fa6_1_or0;
  wire [0:0] h_s_arrmul16_and7_1;
  wire [0:0] h_s_arrmul16_fa7_1_xor1;
  wire [0:0] h_s_arrmul16_fa7_1_or0;
  wire [0:0] h_s_arrmul16_and8_1;
  wire [0:0] h_s_arrmul16_fa8_1_xor1;
  wire [0:0] h_s_arrmul16_fa8_1_or0;
  wire [0:0] h_s_arrmul16_and9_1;
  wire [0:0] h_s_arrmul16_fa9_1_xor1;
  wire [0:0] h_s_arrmul16_fa9_1_or0;
  wire [0:0] h_s_arrmul16_and10_1;
  wire [0:0] h_s_arrmul16_fa10_1_xor1;
  wire [0:0] h_s_arrmul16_fa10_1_or0;
  wire [0:0] h_s_arrmul16_and11_1;
  wire [0:0] h_s_arrmul16_fa11_1_xor1;
  wire [0:0] h_s_arrmul16_fa11_1_or0;
  wire [0:0] h_s_arrmul16_and12_1;
  wire [0:0] h_s_arrmul16_fa12_1_xor1;
  wire [0:0] h_s_arrmul16_fa12_1_or0;
  wire [0:0] h_s_arrmul16_and13_1;
  wire [0:0] h_s_arrmul16_fa13_1_xor1;
  wire [0:0] h_s_arrmul16_fa13_1_or0;
  wire [0:0] h_s_arrmul16_and14_1;
  wire [0:0] h_s_arrmul16_fa14_1_xor1;
  wire [0:0] h_s_arrmul16_fa14_1_or0;
  wire [0:0] h_s_arrmul16_nand15_1;
  wire [0:0] h_s_arrmul16_fa15_1_xor1;
  wire [0:0] h_s_arrmul16_fa15_1_or0;
  wire [0:0] h_s_arrmul16_and0_2;
  wire [0:0] h_s_arrmul16_ha0_2_xor0;
  wire [0:0] h_s_arrmul16_ha0_2_and0;
  wire [0:0] h_s_arrmul16_and1_2;
  wire [0:0] h_s_arrmul16_fa1_2_xor1;
  wire [0:0] h_s_arrmul16_fa1_2_or0;
  wire [0:0] h_s_arrmul16_and2_2;
  wire [0:0] h_s_arrmul16_fa2_2_xor1;
  wire [0:0] h_s_arrmul16_fa2_2_or0;
  wire [0:0] h_s_arrmul16_and3_2;
  wire [0:0] h_s_arrmul16_fa3_2_xor1;
  wire [0:0] h_s_arrmul16_fa3_2_or0;
  wire [0:0] h_s_arrmul16_and4_2;
  wire [0:0] h_s_arrmul16_fa4_2_xor1;
  wire [0:0] h_s_arrmul16_fa4_2_or0;
  wire [0:0] h_s_arrmul16_and5_2;
  wire [0:0] h_s_arrmul16_fa5_2_xor1;
  wire [0:0] h_s_arrmul16_fa5_2_or0;
  wire [0:0] h_s_arrmul16_and6_2;
  wire [0:0] h_s_arrmul16_fa6_2_xor1;
  wire [0:0] h_s_arrmul16_fa6_2_or0;
  wire [0:0] h_s_arrmul16_and7_2;
  wire [0:0] h_s_arrmul16_fa7_2_xor1;
  wire [0:0] h_s_arrmul16_fa7_2_or0;
  wire [0:0] h_s_arrmul16_and8_2;
  wire [0:0] h_s_arrmul16_fa8_2_xor1;
  wire [0:0] h_s_arrmul16_fa8_2_or0;
  wire [0:0] h_s_arrmul16_and9_2;
  wire [0:0] h_s_arrmul16_fa9_2_xor1;
  wire [0:0] h_s_arrmul16_fa9_2_or0;
  wire [0:0] h_s_arrmul16_and10_2;
  wire [0:0] h_s_arrmul16_fa10_2_xor1;
  wire [0:0] h_s_arrmul16_fa10_2_or0;
  wire [0:0] h_s_arrmul16_and11_2;
  wire [0:0] h_s_arrmul16_fa11_2_xor1;
  wire [0:0] h_s_arrmul16_fa11_2_or0;
  wire [0:0] h_s_arrmul16_and12_2;
  wire [0:0] h_s_arrmul16_fa12_2_xor1;
  wire [0:0] h_s_arrmul16_fa12_2_or0;
  wire [0:0] h_s_arrmul16_and13_2;
  wire [0:0] h_s_arrmul16_fa13_2_xor1;
  wire [0:0] h_s_arrmul16_fa13_2_or0;
  wire [0:0] h_s_arrmul16_and14_2;
  wire [0:0] h_s_arrmul16_fa14_2_xor1;
  wire [0:0] h_s_arrmul16_fa14_2_or0;
  wire [0:0] h_s_arrmul16_nand15_2;
  wire [0:0] h_s_arrmul16_fa15_2_xor1;
  wire [0:0] h_s_arrmul16_fa15_2_or0;
  wire [0:0] h_s_arrmul16_and0_3;
  wire [0:0] h_s_arrmul16_ha0_3_xor0;
  wire [0:0] h_s_arrmul16_ha0_3_and0;
  wire [0:0] h_s_arrmul16_and1_3;
  wire [0:0] h_s_arrmul16_fa1_3_xor1;
  wire [0:0] h_s_arrmul16_fa1_3_or0;
  wire [0:0] h_s_arrmul16_and2_3;
  wire [0:0] h_s_arrmul16_fa2_3_xor1;
  wire [0:0] h_s_arrmul16_fa2_3_or0;
  wire [0:0] h_s_arrmul16_and3_3;
  wire [0:0] h_s_arrmul16_fa3_3_xor1;
  wire [0:0] h_s_arrmul16_fa3_3_or0;
  wire [0:0] h_s_arrmul16_and4_3;
  wire [0:0] h_s_arrmul16_fa4_3_xor1;
  wire [0:0] h_s_arrmul16_fa4_3_or0;
  wire [0:0] h_s_arrmul16_and5_3;
  wire [0:0] h_s_arrmul16_fa5_3_xor1;
  wire [0:0] h_s_arrmul16_fa5_3_or0;
  wire [0:0] h_s_arrmul16_and6_3;
  wire [0:0] h_s_arrmul16_fa6_3_xor1;
  wire [0:0] h_s_arrmul16_fa6_3_or0;
  wire [0:0] h_s_arrmul16_and7_3;
  wire [0:0] h_s_arrmul16_fa7_3_xor1;
  wire [0:0] h_s_arrmul16_fa7_3_or0;
  wire [0:0] h_s_arrmul16_and8_3;
  wire [0:0] h_s_arrmul16_fa8_3_xor1;
  wire [0:0] h_s_arrmul16_fa8_3_or0;
  wire [0:0] h_s_arrmul16_and9_3;
  wire [0:0] h_s_arrmul16_fa9_3_xor1;
  wire [0:0] h_s_arrmul16_fa9_3_or0;
  wire [0:0] h_s_arrmul16_and10_3;
  wire [0:0] h_s_arrmul16_fa10_3_xor1;
  wire [0:0] h_s_arrmul16_fa10_3_or0;
  wire [0:0] h_s_arrmul16_and11_3;
  wire [0:0] h_s_arrmul16_fa11_3_xor1;
  wire [0:0] h_s_arrmul16_fa11_3_or0;
  wire [0:0] h_s_arrmul16_and12_3;
  wire [0:0] h_s_arrmul16_fa12_3_xor1;
  wire [0:0] h_s_arrmul16_fa12_3_or0;
  wire [0:0] h_s_arrmul16_and13_3;
  wire [0:0] h_s_arrmul16_fa13_3_xor1;
  wire [0:0] h_s_arrmul16_fa13_3_or0;
  wire [0:0] h_s_arrmul16_and14_3;
  wire [0:0] h_s_arrmul16_fa14_3_xor1;
  wire [0:0] h_s_arrmul16_fa14_3_or0;
  wire [0:0] h_s_arrmul16_nand15_3;
  wire [0:0] h_s_arrmul16_fa15_3_xor1;
  wire [0:0] h_s_arrmul16_fa15_3_or0;
  wire [0:0] h_s_arrmul16_and0_4;
  wire [0:0] h_s_arrmul16_ha0_4_xor0;
  wire [0:0] h_s_arrmul16_ha0_4_and0;
  wire [0:0] h_s_arrmul16_and1_4;
  wire [0:0] h_s_arrmul16_fa1_4_xor1;
  wire [0:0] h_s_arrmul16_fa1_4_or0;
  wire [0:0] h_s_arrmul16_and2_4;
  wire [0:0] h_s_arrmul16_fa2_4_xor1;
  wire [0:0] h_s_arrmul16_fa2_4_or0;
  wire [0:0] h_s_arrmul16_and3_4;
  wire [0:0] h_s_arrmul16_fa3_4_xor1;
  wire [0:0] h_s_arrmul16_fa3_4_or0;
  wire [0:0] h_s_arrmul16_and4_4;
  wire [0:0] h_s_arrmul16_fa4_4_xor1;
  wire [0:0] h_s_arrmul16_fa4_4_or0;
  wire [0:0] h_s_arrmul16_and5_4;
  wire [0:0] h_s_arrmul16_fa5_4_xor1;
  wire [0:0] h_s_arrmul16_fa5_4_or0;
  wire [0:0] h_s_arrmul16_and6_4;
  wire [0:0] h_s_arrmul16_fa6_4_xor1;
  wire [0:0] h_s_arrmul16_fa6_4_or0;
  wire [0:0] h_s_arrmul16_and7_4;
  wire [0:0] h_s_arrmul16_fa7_4_xor1;
  wire [0:0] h_s_arrmul16_fa7_4_or0;
  wire [0:0] h_s_arrmul16_and8_4;
  wire [0:0] h_s_arrmul16_fa8_4_xor1;
  wire [0:0] h_s_arrmul16_fa8_4_or0;
  wire [0:0] h_s_arrmul16_and9_4;
  wire [0:0] h_s_arrmul16_fa9_4_xor1;
  wire [0:0] h_s_arrmul16_fa9_4_or0;
  wire [0:0] h_s_arrmul16_and10_4;
  wire [0:0] h_s_arrmul16_fa10_4_xor1;
  wire [0:0] h_s_arrmul16_fa10_4_or0;
  wire [0:0] h_s_arrmul16_and11_4;
  wire [0:0] h_s_arrmul16_fa11_4_xor1;
  wire [0:0] h_s_arrmul16_fa11_4_or0;
  wire [0:0] h_s_arrmul16_and12_4;
  wire [0:0] h_s_arrmul16_fa12_4_xor1;
  wire [0:0] h_s_arrmul16_fa12_4_or0;
  wire [0:0] h_s_arrmul16_and13_4;
  wire [0:0] h_s_arrmul16_fa13_4_xor1;
  wire [0:0] h_s_arrmul16_fa13_4_or0;
  wire [0:0] h_s_arrmul16_and14_4;
  wire [0:0] h_s_arrmul16_fa14_4_xor1;
  wire [0:0] h_s_arrmul16_fa14_4_or0;
  wire [0:0] h_s_arrmul16_nand15_4;
  wire [0:0] h_s_arrmul16_fa15_4_xor1;
  wire [0:0] h_s_arrmul16_fa15_4_or0;
  wire [0:0] h_s_arrmul16_and0_5;
  wire [0:0] h_s_arrmul16_ha0_5_xor0;
  wire [0:0] h_s_arrmul16_ha0_5_and0;
  wire [0:0] h_s_arrmul16_and1_5;
  wire [0:0] h_s_arrmul16_fa1_5_xor1;
  wire [0:0] h_s_arrmul16_fa1_5_or0;
  wire [0:0] h_s_arrmul16_and2_5;
  wire [0:0] h_s_arrmul16_fa2_5_xor1;
  wire [0:0] h_s_arrmul16_fa2_5_or0;
  wire [0:0] h_s_arrmul16_and3_5;
  wire [0:0] h_s_arrmul16_fa3_5_xor1;
  wire [0:0] h_s_arrmul16_fa3_5_or0;
  wire [0:0] h_s_arrmul16_and4_5;
  wire [0:0] h_s_arrmul16_fa4_5_xor1;
  wire [0:0] h_s_arrmul16_fa4_5_or0;
  wire [0:0] h_s_arrmul16_and5_5;
  wire [0:0] h_s_arrmul16_fa5_5_xor1;
  wire [0:0] h_s_arrmul16_fa5_5_or0;
  wire [0:0] h_s_arrmul16_and6_5;
  wire [0:0] h_s_arrmul16_fa6_5_xor1;
  wire [0:0] h_s_arrmul16_fa6_5_or0;
  wire [0:0] h_s_arrmul16_and7_5;
  wire [0:0] h_s_arrmul16_fa7_5_xor1;
  wire [0:0] h_s_arrmul16_fa7_5_or0;
  wire [0:0] h_s_arrmul16_and8_5;
  wire [0:0] h_s_arrmul16_fa8_5_xor1;
  wire [0:0] h_s_arrmul16_fa8_5_or0;
  wire [0:0] h_s_arrmul16_and9_5;
  wire [0:0] h_s_arrmul16_fa9_5_xor1;
  wire [0:0] h_s_arrmul16_fa9_5_or0;
  wire [0:0] h_s_arrmul16_and10_5;
  wire [0:0] h_s_arrmul16_fa10_5_xor1;
  wire [0:0] h_s_arrmul16_fa10_5_or0;
  wire [0:0] h_s_arrmul16_and11_5;
  wire [0:0] h_s_arrmul16_fa11_5_xor1;
  wire [0:0] h_s_arrmul16_fa11_5_or0;
  wire [0:0] h_s_arrmul16_and12_5;
  wire [0:0] h_s_arrmul16_fa12_5_xor1;
  wire [0:0] h_s_arrmul16_fa12_5_or0;
  wire [0:0] h_s_arrmul16_and13_5;
  wire [0:0] h_s_arrmul16_fa13_5_xor1;
  wire [0:0] h_s_arrmul16_fa13_5_or0;
  wire [0:0] h_s_arrmul16_and14_5;
  wire [0:0] h_s_arrmul16_fa14_5_xor1;
  wire [0:0] h_s_arrmul16_fa14_5_or0;
  wire [0:0] h_s_arrmul16_nand15_5;
  wire [0:0] h_s_arrmul16_fa15_5_xor1;
  wire [0:0] h_s_arrmul16_fa15_5_or0;
  wire [0:0] h_s_arrmul16_and0_6;
  wire [0:0] h_s_arrmul16_ha0_6_xor0;
  wire [0:0] h_s_arrmul16_ha0_6_and0;
  wire [0:0] h_s_arrmul16_and1_6;
  wire [0:0] h_s_arrmul16_fa1_6_xor1;
  wire [0:0] h_s_arrmul16_fa1_6_or0;
  wire [0:0] h_s_arrmul16_and2_6;
  wire [0:0] h_s_arrmul16_fa2_6_xor1;
  wire [0:0] h_s_arrmul16_fa2_6_or0;
  wire [0:0] h_s_arrmul16_and3_6;
  wire [0:0] h_s_arrmul16_fa3_6_xor1;
  wire [0:0] h_s_arrmul16_fa3_6_or0;
  wire [0:0] h_s_arrmul16_and4_6;
  wire [0:0] h_s_arrmul16_fa4_6_xor1;
  wire [0:0] h_s_arrmul16_fa4_6_or0;
  wire [0:0] h_s_arrmul16_and5_6;
  wire [0:0] h_s_arrmul16_fa5_6_xor1;
  wire [0:0] h_s_arrmul16_fa5_6_or0;
  wire [0:0] h_s_arrmul16_and6_6;
  wire [0:0] h_s_arrmul16_fa6_6_xor1;
  wire [0:0] h_s_arrmul16_fa6_6_or0;
  wire [0:0] h_s_arrmul16_and7_6;
  wire [0:0] h_s_arrmul16_fa7_6_xor1;
  wire [0:0] h_s_arrmul16_fa7_6_or0;
  wire [0:0] h_s_arrmul16_and8_6;
  wire [0:0] h_s_arrmul16_fa8_6_xor1;
  wire [0:0] h_s_arrmul16_fa8_6_or0;
  wire [0:0] h_s_arrmul16_and9_6;
  wire [0:0] h_s_arrmul16_fa9_6_xor1;
  wire [0:0] h_s_arrmul16_fa9_6_or0;
  wire [0:0] h_s_arrmul16_and10_6;
  wire [0:0] h_s_arrmul16_fa10_6_xor1;
  wire [0:0] h_s_arrmul16_fa10_6_or0;
  wire [0:0] h_s_arrmul16_and11_6;
  wire [0:0] h_s_arrmul16_fa11_6_xor1;
  wire [0:0] h_s_arrmul16_fa11_6_or0;
  wire [0:0] h_s_arrmul16_and12_6;
  wire [0:0] h_s_arrmul16_fa12_6_xor1;
  wire [0:0] h_s_arrmul16_fa12_6_or0;
  wire [0:0] h_s_arrmul16_and13_6;
  wire [0:0] h_s_arrmul16_fa13_6_xor1;
  wire [0:0] h_s_arrmul16_fa13_6_or0;
  wire [0:0] h_s_arrmul16_and14_6;
  wire [0:0] h_s_arrmul16_fa14_6_xor1;
  wire [0:0] h_s_arrmul16_fa14_6_or0;
  wire [0:0] h_s_arrmul16_nand15_6;
  wire [0:0] h_s_arrmul16_fa15_6_xor1;
  wire [0:0] h_s_arrmul16_fa15_6_or0;
  wire [0:0] h_s_arrmul16_and0_7;
  wire [0:0] h_s_arrmul16_ha0_7_xor0;
  wire [0:0] h_s_arrmul16_ha0_7_and0;
  wire [0:0] h_s_arrmul16_and1_7;
  wire [0:0] h_s_arrmul16_fa1_7_xor1;
  wire [0:0] h_s_arrmul16_fa1_7_or0;
  wire [0:0] h_s_arrmul16_and2_7;
  wire [0:0] h_s_arrmul16_fa2_7_xor1;
  wire [0:0] h_s_arrmul16_fa2_7_or0;
  wire [0:0] h_s_arrmul16_and3_7;
  wire [0:0] h_s_arrmul16_fa3_7_xor1;
  wire [0:0] h_s_arrmul16_fa3_7_or0;
  wire [0:0] h_s_arrmul16_and4_7;
  wire [0:0] h_s_arrmul16_fa4_7_xor1;
  wire [0:0] h_s_arrmul16_fa4_7_or0;
  wire [0:0] h_s_arrmul16_and5_7;
  wire [0:0] h_s_arrmul16_fa5_7_xor1;
  wire [0:0] h_s_arrmul16_fa5_7_or0;
  wire [0:0] h_s_arrmul16_and6_7;
  wire [0:0] h_s_arrmul16_fa6_7_xor1;
  wire [0:0] h_s_arrmul16_fa6_7_or0;
  wire [0:0] h_s_arrmul16_and7_7;
  wire [0:0] h_s_arrmul16_fa7_7_xor1;
  wire [0:0] h_s_arrmul16_fa7_7_or0;
  wire [0:0] h_s_arrmul16_and8_7;
  wire [0:0] h_s_arrmul16_fa8_7_xor1;
  wire [0:0] h_s_arrmul16_fa8_7_or0;
  wire [0:0] h_s_arrmul16_and9_7;
  wire [0:0] h_s_arrmul16_fa9_7_xor1;
  wire [0:0] h_s_arrmul16_fa9_7_or0;
  wire [0:0] h_s_arrmul16_and10_7;
  wire [0:0] h_s_arrmul16_fa10_7_xor1;
  wire [0:0] h_s_arrmul16_fa10_7_or0;
  wire [0:0] h_s_arrmul16_and11_7;
  wire [0:0] h_s_arrmul16_fa11_7_xor1;
  wire [0:0] h_s_arrmul16_fa11_7_or0;
  wire [0:0] h_s_arrmul16_and12_7;
  wire [0:0] h_s_arrmul16_fa12_7_xor1;
  wire [0:0] h_s_arrmul16_fa12_7_or0;
  wire [0:0] h_s_arrmul16_and13_7;
  wire [0:0] h_s_arrmul16_fa13_7_xor1;
  wire [0:0] h_s_arrmul16_fa13_7_or0;
  wire [0:0] h_s_arrmul16_and14_7;
  wire [0:0] h_s_arrmul16_fa14_7_xor1;
  wire [0:0] h_s_arrmul16_fa14_7_or0;
  wire [0:0] h_s_arrmul16_nand15_7;
  wire [0:0] h_s_arrmul16_fa15_7_xor1;
  wire [0:0] h_s_arrmul16_fa15_7_or0;
  wire [0:0] h_s_arrmul16_and0_8;
  wire [0:0] h_s_arrmul16_ha0_8_xor0;
  wire [0:0] h_s_arrmul16_ha0_8_and0;
  wire [0:0] h_s_arrmul16_and1_8;
  wire [0:0] h_s_arrmul16_fa1_8_xor1;
  wire [0:0] h_s_arrmul16_fa1_8_or0;
  wire [0:0] h_s_arrmul16_and2_8;
  wire [0:0] h_s_arrmul16_fa2_8_xor1;
  wire [0:0] h_s_arrmul16_fa2_8_or0;
  wire [0:0] h_s_arrmul16_and3_8;
  wire [0:0] h_s_arrmul16_fa3_8_xor1;
  wire [0:0] h_s_arrmul16_fa3_8_or0;
  wire [0:0] h_s_arrmul16_and4_8;
  wire [0:0] h_s_arrmul16_fa4_8_xor1;
  wire [0:0] h_s_arrmul16_fa4_8_or0;
  wire [0:0] h_s_arrmul16_and5_8;
  wire [0:0] h_s_arrmul16_fa5_8_xor1;
  wire [0:0] h_s_arrmul16_fa5_8_or0;
  wire [0:0] h_s_arrmul16_and6_8;
  wire [0:0] h_s_arrmul16_fa6_8_xor1;
  wire [0:0] h_s_arrmul16_fa6_8_or0;
  wire [0:0] h_s_arrmul16_and7_8;
  wire [0:0] h_s_arrmul16_fa7_8_xor1;
  wire [0:0] h_s_arrmul16_fa7_8_or0;
  wire [0:0] h_s_arrmul16_and8_8;
  wire [0:0] h_s_arrmul16_fa8_8_xor1;
  wire [0:0] h_s_arrmul16_fa8_8_or0;
  wire [0:0] h_s_arrmul16_and9_8;
  wire [0:0] h_s_arrmul16_fa9_8_xor1;
  wire [0:0] h_s_arrmul16_fa9_8_or0;
  wire [0:0] h_s_arrmul16_and10_8;
  wire [0:0] h_s_arrmul16_fa10_8_xor1;
  wire [0:0] h_s_arrmul16_fa10_8_or0;
  wire [0:0] h_s_arrmul16_and11_8;
  wire [0:0] h_s_arrmul16_fa11_8_xor1;
  wire [0:0] h_s_arrmul16_fa11_8_or0;
  wire [0:0] h_s_arrmul16_and12_8;
  wire [0:0] h_s_arrmul16_fa12_8_xor1;
  wire [0:0] h_s_arrmul16_fa12_8_or0;
  wire [0:0] h_s_arrmul16_and13_8;
  wire [0:0] h_s_arrmul16_fa13_8_xor1;
  wire [0:0] h_s_arrmul16_fa13_8_or0;
  wire [0:0] h_s_arrmul16_and14_8;
  wire [0:0] h_s_arrmul16_fa14_8_xor1;
  wire [0:0] h_s_arrmul16_fa14_8_or0;
  wire [0:0] h_s_arrmul16_nand15_8;
  wire [0:0] h_s_arrmul16_fa15_8_xor1;
  wire [0:0] h_s_arrmul16_fa15_8_or0;
  wire [0:0] h_s_arrmul16_and0_9;
  wire [0:0] h_s_arrmul16_ha0_9_xor0;
  wire [0:0] h_s_arrmul16_ha0_9_and0;
  wire [0:0] h_s_arrmul16_and1_9;
  wire [0:0] h_s_arrmul16_fa1_9_xor1;
  wire [0:0] h_s_arrmul16_fa1_9_or0;
  wire [0:0] h_s_arrmul16_and2_9;
  wire [0:0] h_s_arrmul16_fa2_9_xor1;
  wire [0:0] h_s_arrmul16_fa2_9_or0;
  wire [0:0] h_s_arrmul16_and3_9;
  wire [0:0] h_s_arrmul16_fa3_9_xor1;
  wire [0:0] h_s_arrmul16_fa3_9_or0;
  wire [0:0] h_s_arrmul16_and4_9;
  wire [0:0] h_s_arrmul16_fa4_9_xor1;
  wire [0:0] h_s_arrmul16_fa4_9_or0;
  wire [0:0] h_s_arrmul16_and5_9;
  wire [0:0] h_s_arrmul16_fa5_9_xor1;
  wire [0:0] h_s_arrmul16_fa5_9_or0;
  wire [0:0] h_s_arrmul16_and6_9;
  wire [0:0] h_s_arrmul16_fa6_9_xor1;
  wire [0:0] h_s_arrmul16_fa6_9_or0;
  wire [0:0] h_s_arrmul16_and7_9;
  wire [0:0] h_s_arrmul16_fa7_9_xor1;
  wire [0:0] h_s_arrmul16_fa7_9_or0;
  wire [0:0] h_s_arrmul16_and8_9;
  wire [0:0] h_s_arrmul16_fa8_9_xor1;
  wire [0:0] h_s_arrmul16_fa8_9_or0;
  wire [0:0] h_s_arrmul16_and9_9;
  wire [0:0] h_s_arrmul16_fa9_9_xor1;
  wire [0:0] h_s_arrmul16_fa9_9_or0;
  wire [0:0] h_s_arrmul16_and10_9;
  wire [0:0] h_s_arrmul16_fa10_9_xor1;
  wire [0:0] h_s_arrmul16_fa10_9_or0;
  wire [0:0] h_s_arrmul16_and11_9;
  wire [0:0] h_s_arrmul16_fa11_9_xor1;
  wire [0:0] h_s_arrmul16_fa11_9_or0;
  wire [0:0] h_s_arrmul16_and12_9;
  wire [0:0] h_s_arrmul16_fa12_9_xor1;
  wire [0:0] h_s_arrmul16_fa12_9_or0;
  wire [0:0] h_s_arrmul16_and13_9;
  wire [0:0] h_s_arrmul16_fa13_9_xor1;
  wire [0:0] h_s_arrmul16_fa13_9_or0;
  wire [0:0] h_s_arrmul16_and14_9;
  wire [0:0] h_s_arrmul16_fa14_9_xor1;
  wire [0:0] h_s_arrmul16_fa14_9_or0;
  wire [0:0] h_s_arrmul16_nand15_9;
  wire [0:0] h_s_arrmul16_fa15_9_xor1;
  wire [0:0] h_s_arrmul16_fa15_9_or0;
  wire [0:0] h_s_arrmul16_and0_10;
  wire [0:0] h_s_arrmul16_ha0_10_xor0;
  wire [0:0] h_s_arrmul16_ha0_10_and0;
  wire [0:0] h_s_arrmul16_and1_10;
  wire [0:0] h_s_arrmul16_fa1_10_xor1;
  wire [0:0] h_s_arrmul16_fa1_10_or0;
  wire [0:0] h_s_arrmul16_and2_10;
  wire [0:0] h_s_arrmul16_fa2_10_xor1;
  wire [0:0] h_s_arrmul16_fa2_10_or0;
  wire [0:0] h_s_arrmul16_and3_10;
  wire [0:0] h_s_arrmul16_fa3_10_xor1;
  wire [0:0] h_s_arrmul16_fa3_10_or0;
  wire [0:0] h_s_arrmul16_and4_10;
  wire [0:0] h_s_arrmul16_fa4_10_xor1;
  wire [0:0] h_s_arrmul16_fa4_10_or0;
  wire [0:0] h_s_arrmul16_and5_10;
  wire [0:0] h_s_arrmul16_fa5_10_xor1;
  wire [0:0] h_s_arrmul16_fa5_10_or0;
  wire [0:0] h_s_arrmul16_and6_10;
  wire [0:0] h_s_arrmul16_fa6_10_xor1;
  wire [0:0] h_s_arrmul16_fa6_10_or0;
  wire [0:0] h_s_arrmul16_and7_10;
  wire [0:0] h_s_arrmul16_fa7_10_xor1;
  wire [0:0] h_s_arrmul16_fa7_10_or0;
  wire [0:0] h_s_arrmul16_and8_10;
  wire [0:0] h_s_arrmul16_fa8_10_xor1;
  wire [0:0] h_s_arrmul16_fa8_10_or0;
  wire [0:0] h_s_arrmul16_and9_10;
  wire [0:0] h_s_arrmul16_fa9_10_xor1;
  wire [0:0] h_s_arrmul16_fa9_10_or0;
  wire [0:0] h_s_arrmul16_and10_10;
  wire [0:0] h_s_arrmul16_fa10_10_xor1;
  wire [0:0] h_s_arrmul16_fa10_10_or0;
  wire [0:0] h_s_arrmul16_and11_10;
  wire [0:0] h_s_arrmul16_fa11_10_xor1;
  wire [0:0] h_s_arrmul16_fa11_10_or0;
  wire [0:0] h_s_arrmul16_and12_10;
  wire [0:0] h_s_arrmul16_fa12_10_xor1;
  wire [0:0] h_s_arrmul16_fa12_10_or0;
  wire [0:0] h_s_arrmul16_and13_10;
  wire [0:0] h_s_arrmul16_fa13_10_xor1;
  wire [0:0] h_s_arrmul16_fa13_10_or0;
  wire [0:0] h_s_arrmul16_and14_10;
  wire [0:0] h_s_arrmul16_fa14_10_xor1;
  wire [0:0] h_s_arrmul16_fa14_10_or0;
  wire [0:0] h_s_arrmul16_nand15_10;
  wire [0:0] h_s_arrmul16_fa15_10_xor1;
  wire [0:0] h_s_arrmul16_fa15_10_or0;
  wire [0:0] h_s_arrmul16_and0_11;
  wire [0:0] h_s_arrmul16_ha0_11_xor0;
  wire [0:0] h_s_arrmul16_ha0_11_and0;
  wire [0:0] h_s_arrmul16_and1_11;
  wire [0:0] h_s_arrmul16_fa1_11_xor1;
  wire [0:0] h_s_arrmul16_fa1_11_or0;
  wire [0:0] h_s_arrmul16_and2_11;
  wire [0:0] h_s_arrmul16_fa2_11_xor1;
  wire [0:0] h_s_arrmul16_fa2_11_or0;
  wire [0:0] h_s_arrmul16_and3_11;
  wire [0:0] h_s_arrmul16_fa3_11_xor1;
  wire [0:0] h_s_arrmul16_fa3_11_or0;
  wire [0:0] h_s_arrmul16_and4_11;
  wire [0:0] h_s_arrmul16_fa4_11_xor1;
  wire [0:0] h_s_arrmul16_fa4_11_or0;
  wire [0:0] h_s_arrmul16_and5_11;
  wire [0:0] h_s_arrmul16_fa5_11_xor1;
  wire [0:0] h_s_arrmul16_fa5_11_or0;
  wire [0:0] h_s_arrmul16_and6_11;
  wire [0:0] h_s_arrmul16_fa6_11_xor1;
  wire [0:0] h_s_arrmul16_fa6_11_or0;
  wire [0:0] h_s_arrmul16_and7_11;
  wire [0:0] h_s_arrmul16_fa7_11_xor1;
  wire [0:0] h_s_arrmul16_fa7_11_or0;
  wire [0:0] h_s_arrmul16_and8_11;
  wire [0:0] h_s_arrmul16_fa8_11_xor1;
  wire [0:0] h_s_arrmul16_fa8_11_or0;
  wire [0:0] h_s_arrmul16_and9_11;
  wire [0:0] h_s_arrmul16_fa9_11_xor1;
  wire [0:0] h_s_arrmul16_fa9_11_or0;
  wire [0:0] h_s_arrmul16_and10_11;
  wire [0:0] h_s_arrmul16_fa10_11_xor1;
  wire [0:0] h_s_arrmul16_fa10_11_or0;
  wire [0:0] h_s_arrmul16_and11_11;
  wire [0:0] h_s_arrmul16_fa11_11_xor1;
  wire [0:0] h_s_arrmul16_fa11_11_or0;
  wire [0:0] h_s_arrmul16_and12_11;
  wire [0:0] h_s_arrmul16_fa12_11_xor1;
  wire [0:0] h_s_arrmul16_fa12_11_or0;
  wire [0:0] h_s_arrmul16_and13_11;
  wire [0:0] h_s_arrmul16_fa13_11_xor1;
  wire [0:0] h_s_arrmul16_fa13_11_or0;
  wire [0:0] h_s_arrmul16_and14_11;
  wire [0:0] h_s_arrmul16_fa14_11_xor1;
  wire [0:0] h_s_arrmul16_fa14_11_or0;
  wire [0:0] h_s_arrmul16_nand15_11;
  wire [0:0] h_s_arrmul16_fa15_11_xor1;
  wire [0:0] h_s_arrmul16_fa15_11_or0;
  wire [0:0] h_s_arrmul16_and0_12;
  wire [0:0] h_s_arrmul16_ha0_12_xor0;
  wire [0:0] h_s_arrmul16_ha0_12_and0;
  wire [0:0] h_s_arrmul16_and1_12;
  wire [0:0] h_s_arrmul16_fa1_12_xor1;
  wire [0:0] h_s_arrmul16_fa1_12_or0;
  wire [0:0] h_s_arrmul16_and2_12;
  wire [0:0] h_s_arrmul16_fa2_12_xor1;
  wire [0:0] h_s_arrmul16_fa2_12_or0;
  wire [0:0] h_s_arrmul16_and3_12;
  wire [0:0] h_s_arrmul16_fa3_12_xor1;
  wire [0:0] h_s_arrmul16_fa3_12_or0;
  wire [0:0] h_s_arrmul16_and4_12;
  wire [0:0] h_s_arrmul16_fa4_12_xor1;
  wire [0:0] h_s_arrmul16_fa4_12_or0;
  wire [0:0] h_s_arrmul16_and5_12;
  wire [0:0] h_s_arrmul16_fa5_12_xor1;
  wire [0:0] h_s_arrmul16_fa5_12_or0;
  wire [0:0] h_s_arrmul16_and6_12;
  wire [0:0] h_s_arrmul16_fa6_12_xor1;
  wire [0:0] h_s_arrmul16_fa6_12_or0;
  wire [0:0] h_s_arrmul16_and7_12;
  wire [0:0] h_s_arrmul16_fa7_12_xor1;
  wire [0:0] h_s_arrmul16_fa7_12_or0;
  wire [0:0] h_s_arrmul16_and8_12;
  wire [0:0] h_s_arrmul16_fa8_12_xor1;
  wire [0:0] h_s_arrmul16_fa8_12_or0;
  wire [0:0] h_s_arrmul16_and9_12;
  wire [0:0] h_s_arrmul16_fa9_12_xor1;
  wire [0:0] h_s_arrmul16_fa9_12_or0;
  wire [0:0] h_s_arrmul16_and10_12;
  wire [0:0] h_s_arrmul16_fa10_12_xor1;
  wire [0:0] h_s_arrmul16_fa10_12_or0;
  wire [0:0] h_s_arrmul16_and11_12;
  wire [0:0] h_s_arrmul16_fa11_12_xor1;
  wire [0:0] h_s_arrmul16_fa11_12_or0;
  wire [0:0] h_s_arrmul16_and12_12;
  wire [0:0] h_s_arrmul16_fa12_12_xor1;
  wire [0:0] h_s_arrmul16_fa12_12_or0;
  wire [0:0] h_s_arrmul16_and13_12;
  wire [0:0] h_s_arrmul16_fa13_12_xor1;
  wire [0:0] h_s_arrmul16_fa13_12_or0;
  wire [0:0] h_s_arrmul16_and14_12;
  wire [0:0] h_s_arrmul16_fa14_12_xor1;
  wire [0:0] h_s_arrmul16_fa14_12_or0;
  wire [0:0] h_s_arrmul16_nand15_12;
  wire [0:0] h_s_arrmul16_fa15_12_xor1;
  wire [0:0] h_s_arrmul16_fa15_12_or0;
  wire [0:0] h_s_arrmul16_and0_13;
  wire [0:0] h_s_arrmul16_ha0_13_xor0;
  wire [0:0] h_s_arrmul16_ha0_13_and0;
  wire [0:0] h_s_arrmul16_and1_13;
  wire [0:0] h_s_arrmul16_fa1_13_xor1;
  wire [0:0] h_s_arrmul16_fa1_13_or0;
  wire [0:0] h_s_arrmul16_and2_13;
  wire [0:0] h_s_arrmul16_fa2_13_xor1;
  wire [0:0] h_s_arrmul16_fa2_13_or0;
  wire [0:0] h_s_arrmul16_and3_13;
  wire [0:0] h_s_arrmul16_fa3_13_xor1;
  wire [0:0] h_s_arrmul16_fa3_13_or0;
  wire [0:0] h_s_arrmul16_and4_13;
  wire [0:0] h_s_arrmul16_fa4_13_xor1;
  wire [0:0] h_s_arrmul16_fa4_13_or0;
  wire [0:0] h_s_arrmul16_and5_13;
  wire [0:0] h_s_arrmul16_fa5_13_xor1;
  wire [0:0] h_s_arrmul16_fa5_13_or0;
  wire [0:0] h_s_arrmul16_and6_13;
  wire [0:0] h_s_arrmul16_fa6_13_xor1;
  wire [0:0] h_s_arrmul16_fa6_13_or0;
  wire [0:0] h_s_arrmul16_and7_13;
  wire [0:0] h_s_arrmul16_fa7_13_xor1;
  wire [0:0] h_s_arrmul16_fa7_13_or0;
  wire [0:0] h_s_arrmul16_and8_13;
  wire [0:0] h_s_arrmul16_fa8_13_xor1;
  wire [0:0] h_s_arrmul16_fa8_13_or0;
  wire [0:0] h_s_arrmul16_and9_13;
  wire [0:0] h_s_arrmul16_fa9_13_xor1;
  wire [0:0] h_s_arrmul16_fa9_13_or0;
  wire [0:0] h_s_arrmul16_and10_13;
  wire [0:0] h_s_arrmul16_fa10_13_xor1;
  wire [0:0] h_s_arrmul16_fa10_13_or0;
  wire [0:0] h_s_arrmul16_and11_13;
  wire [0:0] h_s_arrmul16_fa11_13_xor1;
  wire [0:0] h_s_arrmul16_fa11_13_or0;
  wire [0:0] h_s_arrmul16_and12_13;
  wire [0:0] h_s_arrmul16_fa12_13_xor1;
  wire [0:0] h_s_arrmul16_fa12_13_or0;
  wire [0:0] h_s_arrmul16_and13_13;
  wire [0:0] h_s_arrmul16_fa13_13_xor1;
  wire [0:0] h_s_arrmul16_fa13_13_or0;
  wire [0:0] h_s_arrmul16_and14_13;
  wire [0:0] h_s_arrmul16_fa14_13_xor1;
  wire [0:0] h_s_arrmul16_fa14_13_or0;
  wire [0:0] h_s_arrmul16_nand15_13;
  wire [0:0] h_s_arrmul16_fa15_13_xor1;
  wire [0:0] h_s_arrmul16_fa15_13_or0;
  wire [0:0] h_s_arrmul16_and0_14;
  wire [0:0] h_s_arrmul16_ha0_14_xor0;
  wire [0:0] h_s_arrmul16_ha0_14_and0;
  wire [0:0] h_s_arrmul16_and1_14;
  wire [0:0] h_s_arrmul16_fa1_14_xor1;
  wire [0:0] h_s_arrmul16_fa1_14_or0;
  wire [0:0] h_s_arrmul16_and2_14;
  wire [0:0] h_s_arrmul16_fa2_14_xor1;
  wire [0:0] h_s_arrmul16_fa2_14_or0;
  wire [0:0] h_s_arrmul16_and3_14;
  wire [0:0] h_s_arrmul16_fa3_14_xor1;
  wire [0:0] h_s_arrmul16_fa3_14_or0;
  wire [0:0] h_s_arrmul16_and4_14;
  wire [0:0] h_s_arrmul16_fa4_14_xor1;
  wire [0:0] h_s_arrmul16_fa4_14_or0;
  wire [0:0] h_s_arrmul16_and5_14;
  wire [0:0] h_s_arrmul16_fa5_14_xor1;
  wire [0:0] h_s_arrmul16_fa5_14_or0;
  wire [0:0] h_s_arrmul16_and6_14;
  wire [0:0] h_s_arrmul16_fa6_14_xor1;
  wire [0:0] h_s_arrmul16_fa6_14_or0;
  wire [0:0] h_s_arrmul16_and7_14;
  wire [0:0] h_s_arrmul16_fa7_14_xor1;
  wire [0:0] h_s_arrmul16_fa7_14_or0;
  wire [0:0] h_s_arrmul16_and8_14;
  wire [0:0] h_s_arrmul16_fa8_14_xor1;
  wire [0:0] h_s_arrmul16_fa8_14_or0;
  wire [0:0] h_s_arrmul16_and9_14;
  wire [0:0] h_s_arrmul16_fa9_14_xor1;
  wire [0:0] h_s_arrmul16_fa9_14_or0;
  wire [0:0] h_s_arrmul16_and10_14;
  wire [0:0] h_s_arrmul16_fa10_14_xor1;
  wire [0:0] h_s_arrmul16_fa10_14_or0;
  wire [0:0] h_s_arrmul16_and11_14;
  wire [0:0] h_s_arrmul16_fa11_14_xor1;
  wire [0:0] h_s_arrmul16_fa11_14_or0;
  wire [0:0] h_s_arrmul16_and12_14;
  wire [0:0] h_s_arrmul16_fa12_14_xor1;
  wire [0:0] h_s_arrmul16_fa12_14_or0;
  wire [0:0] h_s_arrmul16_and13_14;
  wire [0:0] h_s_arrmul16_fa13_14_xor1;
  wire [0:0] h_s_arrmul16_fa13_14_or0;
  wire [0:0] h_s_arrmul16_and14_14;
  wire [0:0] h_s_arrmul16_fa14_14_xor1;
  wire [0:0] h_s_arrmul16_fa14_14_or0;
  wire [0:0] h_s_arrmul16_nand15_14;
  wire [0:0] h_s_arrmul16_fa15_14_xor1;
  wire [0:0] h_s_arrmul16_fa15_14_or0;
  wire [0:0] h_s_arrmul16_nand0_15;
  wire [0:0] h_s_arrmul16_ha0_15_xor0;
  wire [0:0] h_s_arrmul16_ha0_15_and0;
  wire [0:0] h_s_arrmul16_nand1_15;
  wire [0:0] h_s_arrmul16_fa1_15_xor1;
  wire [0:0] h_s_arrmul16_fa1_15_or0;
  wire [0:0] h_s_arrmul16_nand2_15;
  wire [0:0] h_s_arrmul16_fa2_15_xor1;
  wire [0:0] h_s_arrmul16_fa2_15_or0;
  wire [0:0] h_s_arrmul16_nand3_15;
  wire [0:0] h_s_arrmul16_fa3_15_xor1;
  wire [0:0] h_s_arrmul16_fa3_15_or0;
  wire [0:0] h_s_arrmul16_nand4_15;
  wire [0:0] h_s_arrmul16_fa4_15_xor1;
  wire [0:0] h_s_arrmul16_fa4_15_or0;
  wire [0:0] h_s_arrmul16_nand5_15;
  wire [0:0] h_s_arrmul16_fa5_15_xor1;
  wire [0:0] h_s_arrmul16_fa5_15_or0;
  wire [0:0] h_s_arrmul16_nand6_15;
  wire [0:0] h_s_arrmul16_fa6_15_xor1;
  wire [0:0] h_s_arrmul16_fa6_15_or0;
  wire [0:0] h_s_arrmul16_nand7_15;
  wire [0:0] h_s_arrmul16_fa7_15_xor1;
  wire [0:0] h_s_arrmul16_fa7_15_or0;
  wire [0:0] h_s_arrmul16_nand8_15;
  wire [0:0] h_s_arrmul16_fa8_15_xor1;
  wire [0:0] h_s_arrmul16_fa8_15_or0;
  wire [0:0] h_s_arrmul16_nand9_15;
  wire [0:0] h_s_arrmul16_fa9_15_xor1;
  wire [0:0] h_s_arrmul16_fa9_15_or0;
  wire [0:0] h_s_arrmul16_nand10_15;
  wire [0:0] h_s_arrmul16_fa10_15_xor1;
  wire [0:0] h_s_arrmul16_fa10_15_or0;
  wire [0:0] h_s_arrmul16_nand11_15;
  wire [0:0] h_s_arrmul16_fa11_15_xor1;
  wire [0:0] h_s_arrmul16_fa11_15_or0;
  wire [0:0] h_s_arrmul16_nand12_15;
  wire [0:0] h_s_arrmul16_fa12_15_xor1;
  wire [0:0] h_s_arrmul16_fa12_15_or0;
  wire [0:0] h_s_arrmul16_nand13_15;
  wire [0:0] h_s_arrmul16_fa13_15_xor1;
  wire [0:0] h_s_arrmul16_fa13_15_or0;
  wire [0:0] h_s_arrmul16_nand14_15;
  wire [0:0] h_s_arrmul16_fa14_15_xor1;
  wire [0:0] h_s_arrmul16_fa14_15_or0;
  wire [0:0] h_s_arrmul16_and15_15;
  wire [0:0] h_s_arrmul16_fa15_15_xor1;
  wire [0:0] h_s_arrmul16_fa15_15_or0;
  wire [0:0] h_s_arrmul16_xor16_15;

  and_gate and_gate_h_s_arrmul16_and0_0(.a(a[0]), .b(b[0]), .out(h_s_arrmul16_and0_0));
  and_gate and_gate_h_s_arrmul16_and1_0(.a(a[1]), .b(b[0]), .out(h_s_arrmul16_and1_0));
  and_gate and_gate_h_s_arrmul16_and2_0(.a(a[2]), .b(b[0]), .out(h_s_arrmul16_and2_0));
  and_gate and_gate_h_s_arrmul16_and3_0(.a(a[3]), .b(b[0]), .out(h_s_arrmul16_and3_0));
  and_gate and_gate_h_s_arrmul16_and4_0(.a(a[4]), .b(b[0]), .out(h_s_arrmul16_and4_0));
  and_gate and_gate_h_s_arrmul16_and5_0(.a(a[5]), .b(b[0]), .out(h_s_arrmul16_and5_0));
  and_gate and_gate_h_s_arrmul16_and6_0(.a(a[6]), .b(b[0]), .out(h_s_arrmul16_and6_0));
  and_gate and_gate_h_s_arrmul16_and7_0(.a(a[7]), .b(b[0]), .out(h_s_arrmul16_and7_0));
  and_gate and_gate_h_s_arrmul16_and8_0(.a(a[8]), .b(b[0]), .out(h_s_arrmul16_and8_0));
  and_gate and_gate_h_s_arrmul16_and9_0(.a(a[9]), .b(b[0]), .out(h_s_arrmul16_and9_0));
  and_gate and_gate_h_s_arrmul16_and10_0(.a(a[10]), .b(b[0]), .out(h_s_arrmul16_and10_0));
  and_gate and_gate_h_s_arrmul16_and11_0(.a(a[11]), .b(b[0]), .out(h_s_arrmul16_and11_0));
  and_gate and_gate_h_s_arrmul16_and12_0(.a(a[12]), .b(b[0]), .out(h_s_arrmul16_and12_0));
  and_gate and_gate_h_s_arrmul16_and13_0(.a(a[13]), .b(b[0]), .out(h_s_arrmul16_and13_0));
  and_gate and_gate_h_s_arrmul16_and14_0(.a(a[14]), .b(b[0]), .out(h_s_arrmul16_and14_0));
  nand_gate nand_gate_h_s_arrmul16_nand15_0(.a(a[15]), .b(b[0]), .out(h_s_arrmul16_nand15_0));
  and_gate and_gate_h_s_arrmul16_and0_1(.a(a[0]), .b(b[1]), .out(h_s_arrmul16_and0_1));
  ha ha_h_s_arrmul16_ha0_1_out(.a(h_s_arrmul16_and0_1[0]), .b(h_s_arrmul16_and1_0[0]), .ha_xor0(h_s_arrmul16_ha0_1_xor0), .ha_and0(h_s_arrmul16_ha0_1_and0));
  and_gate and_gate_h_s_arrmul16_and1_1(.a(a[1]), .b(b[1]), .out(h_s_arrmul16_and1_1));
  fa fa_h_s_arrmul16_fa1_1_out(.a(h_s_arrmul16_and1_1[0]), .b(h_s_arrmul16_and2_0[0]), .cin(h_s_arrmul16_ha0_1_and0[0]), .fa_xor1(h_s_arrmul16_fa1_1_xor1), .fa_or0(h_s_arrmul16_fa1_1_or0));
  and_gate and_gate_h_s_arrmul16_and2_1(.a(a[2]), .b(b[1]), .out(h_s_arrmul16_and2_1));
  fa fa_h_s_arrmul16_fa2_1_out(.a(h_s_arrmul16_and2_1[0]), .b(h_s_arrmul16_and3_0[0]), .cin(h_s_arrmul16_fa1_1_or0[0]), .fa_xor1(h_s_arrmul16_fa2_1_xor1), .fa_or0(h_s_arrmul16_fa2_1_or0));
  and_gate and_gate_h_s_arrmul16_and3_1(.a(a[3]), .b(b[1]), .out(h_s_arrmul16_and3_1));
  fa fa_h_s_arrmul16_fa3_1_out(.a(h_s_arrmul16_and3_1[0]), .b(h_s_arrmul16_and4_0[0]), .cin(h_s_arrmul16_fa2_1_or0[0]), .fa_xor1(h_s_arrmul16_fa3_1_xor1), .fa_or0(h_s_arrmul16_fa3_1_or0));
  and_gate and_gate_h_s_arrmul16_and4_1(.a(a[4]), .b(b[1]), .out(h_s_arrmul16_and4_1));
  fa fa_h_s_arrmul16_fa4_1_out(.a(h_s_arrmul16_and4_1[0]), .b(h_s_arrmul16_and5_0[0]), .cin(h_s_arrmul16_fa3_1_or0[0]), .fa_xor1(h_s_arrmul16_fa4_1_xor1), .fa_or0(h_s_arrmul16_fa4_1_or0));
  and_gate and_gate_h_s_arrmul16_and5_1(.a(a[5]), .b(b[1]), .out(h_s_arrmul16_and5_1));
  fa fa_h_s_arrmul16_fa5_1_out(.a(h_s_arrmul16_and5_1[0]), .b(h_s_arrmul16_and6_0[0]), .cin(h_s_arrmul16_fa4_1_or0[0]), .fa_xor1(h_s_arrmul16_fa5_1_xor1), .fa_or0(h_s_arrmul16_fa5_1_or0));
  and_gate and_gate_h_s_arrmul16_and6_1(.a(a[6]), .b(b[1]), .out(h_s_arrmul16_and6_1));
  fa fa_h_s_arrmul16_fa6_1_out(.a(h_s_arrmul16_and6_1[0]), .b(h_s_arrmul16_and7_0[0]), .cin(h_s_arrmul16_fa5_1_or0[0]), .fa_xor1(h_s_arrmul16_fa6_1_xor1), .fa_or0(h_s_arrmul16_fa6_1_or0));
  and_gate and_gate_h_s_arrmul16_and7_1(.a(a[7]), .b(b[1]), .out(h_s_arrmul16_and7_1));
  fa fa_h_s_arrmul16_fa7_1_out(.a(h_s_arrmul16_and7_1[0]), .b(h_s_arrmul16_and8_0[0]), .cin(h_s_arrmul16_fa6_1_or0[0]), .fa_xor1(h_s_arrmul16_fa7_1_xor1), .fa_or0(h_s_arrmul16_fa7_1_or0));
  and_gate and_gate_h_s_arrmul16_and8_1(.a(a[8]), .b(b[1]), .out(h_s_arrmul16_and8_1));
  fa fa_h_s_arrmul16_fa8_1_out(.a(h_s_arrmul16_and8_1[0]), .b(h_s_arrmul16_and9_0[0]), .cin(h_s_arrmul16_fa7_1_or0[0]), .fa_xor1(h_s_arrmul16_fa8_1_xor1), .fa_or0(h_s_arrmul16_fa8_1_or0));
  and_gate and_gate_h_s_arrmul16_and9_1(.a(a[9]), .b(b[1]), .out(h_s_arrmul16_and9_1));
  fa fa_h_s_arrmul16_fa9_1_out(.a(h_s_arrmul16_and9_1[0]), .b(h_s_arrmul16_and10_0[0]), .cin(h_s_arrmul16_fa8_1_or0[0]), .fa_xor1(h_s_arrmul16_fa9_1_xor1), .fa_or0(h_s_arrmul16_fa9_1_or0));
  and_gate and_gate_h_s_arrmul16_and10_1(.a(a[10]), .b(b[1]), .out(h_s_arrmul16_and10_1));
  fa fa_h_s_arrmul16_fa10_1_out(.a(h_s_arrmul16_and10_1[0]), .b(h_s_arrmul16_and11_0[0]), .cin(h_s_arrmul16_fa9_1_or0[0]), .fa_xor1(h_s_arrmul16_fa10_1_xor1), .fa_or0(h_s_arrmul16_fa10_1_or0));
  and_gate and_gate_h_s_arrmul16_and11_1(.a(a[11]), .b(b[1]), .out(h_s_arrmul16_and11_1));
  fa fa_h_s_arrmul16_fa11_1_out(.a(h_s_arrmul16_and11_1[0]), .b(h_s_arrmul16_and12_0[0]), .cin(h_s_arrmul16_fa10_1_or0[0]), .fa_xor1(h_s_arrmul16_fa11_1_xor1), .fa_or0(h_s_arrmul16_fa11_1_or0));
  and_gate and_gate_h_s_arrmul16_and12_1(.a(a[12]), .b(b[1]), .out(h_s_arrmul16_and12_1));
  fa fa_h_s_arrmul16_fa12_1_out(.a(h_s_arrmul16_and12_1[0]), .b(h_s_arrmul16_and13_0[0]), .cin(h_s_arrmul16_fa11_1_or0[0]), .fa_xor1(h_s_arrmul16_fa12_1_xor1), .fa_or0(h_s_arrmul16_fa12_1_or0));
  and_gate and_gate_h_s_arrmul16_and13_1(.a(a[13]), .b(b[1]), .out(h_s_arrmul16_and13_1));
  fa fa_h_s_arrmul16_fa13_1_out(.a(h_s_arrmul16_and13_1[0]), .b(h_s_arrmul16_and14_0[0]), .cin(h_s_arrmul16_fa12_1_or0[0]), .fa_xor1(h_s_arrmul16_fa13_1_xor1), .fa_or0(h_s_arrmul16_fa13_1_or0));
  and_gate and_gate_h_s_arrmul16_and14_1(.a(a[14]), .b(b[1]), .out(h_s_arrmul16_and14_1));
  fa fa_h_s_arrmul16_fa14_1_out(.a(h_s_arrmul16_and14_1[0]), .b(h_s_arrmul16_nand15_0[0]), .cin(h_s_arrmul16_fa13_1_or0[0]), .fa_xor1(h_s_arrmul16_fa14_1_xor1), .fa_or0(h_s_arrmul16_fa14_1_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_1(.a(a[15]), .b(b[1]), .out(h_s_arrmul16_nand15_1));
  fa fa_h_s_arrmul16_fa15_1_out(.a(h_s_arrmul16_nand15_1[0]), .b(1'b1), .cin(h_s_arrmul16_fa14_1_or0[0]), .fa_xor1(h_s_arrmul16_fa15_1_xor1), .fa_or0(h_s_arrmul16_fa15_1_or0));
  and_gate and_gate_h_s_arrmul16_and0_2(.a(a[0]), .b(b[2]), .out(h_s_arrmul16_and0_2));
  ha ha_h_s_arrmul16_ha0_2_out(.a(h_s_arrmul16_and0_2[0]), .b(h_s_arrmul16_fa1_1_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_2_xor0), .ha_and0(h_s_arrmul16_ha0_2_and0));
  and_gate and_gate_h_s_arrmul16_and1_2(.a(a[1]), .b(b[2]), .out(h_s_arrmul16_and1_2));
  fa fa_h_s_arrmul16_fa1_2_out(.a(h_s_arrmul16_and1_2[0]), .b(h_s_arrmul16_fa2_1_xor1[0]), .cin(h_s_arrmul16_ha0_2_and0[0]), .fa_xor1(h_s_arrmul16_fa1_2_xor1), .fa_or0(h_s_arrmul16_fa1_2_or0));
  and_gate and_gate_h_s_arrmul16_and2_2(.a(a[2]), .b(b[2]), .out(h_s_arrmul16_and2_2));
  fa fa_h_s_arrmul16_fa2_2_out(.a(h_s_arrmul16_and2_2[0]), .b(h_s_arrmul16_fa3_1_xor1[0]), .cin(h_s_arrmul16_fa1_2_or0[0]), .fa_xor1(h_s_arrmul16_fa2_2_xor1), .fa_or0(h_s_arrmul16_fa2_2_or0));
  and_gate and_gate_h_s_arrmul16_and3_2(.a(a[3]), .b(b[2]), .out(h_s_arrmul16_and3_2));
  fa fa_h_s_arrmul16_fa3_2_out(.a(h_s_arrmul16_and3_2[0]), .b(h_s_arrmul16_fa4_1_xor1[0]), .cin(h_s_arrmul16_fa2_2_or0[0]), .fa_xor1(h_s_arrmul16_fa3_2_xor1), .fa_or0(h_s_arrmul16_fa3_2_or0));
  and_gate and_gate_h_s_arrmul16_and4_2(.a(a[4]), .b(b[2]), .out(h_s_arrmul16_and4_2));
  fa fa_h_s_arrmul16_fa4_2_out(.a(h_s_arrmul16_and4_2[0]), .b(h_s_arrmul16_fa5_1_xor1[0]), .cin(h_s_arrmul16_fa3_2_or0[0]), .fa_xor1(h_s_arrmul16_fa4_2_xor1), .fa_or0(h_s_arrmul16_fa4_2_or0));
  and_gate and_gate_h_s_arrmul16_and5_2(.a(a[5]), .b(b[2]), .out(h_s_arrmul16_and5_2));
  fa fa_h_s_arrmul16_fa5_2_out(.a(h_s_arrmul16_and5_2[0]), .b(h_s_arrmul16_fa6_1_xor1[0]), .cin(h_s_arrmul16_fa4_2_or0[0]), .fa_xor1(h_s_arrmul16_fa5_2_xor1), .fa_or0(h_s_arrmul16_fa5_2_or0));
  and_gate and_gate_h_s_arrmul16_and6_2(.a(a[6]), .b(b[2]), .out(h_s_arrmul16_and6_2));
  fa fa_h_s_arrmul16_fa6_2_out(.a(h_s_arrmul16_and6_2[0]), .b(h_s_arrmul16_fa7_1_xor1[0]), .cin(h_s_arrmul16_fa5_2_or0[0]), .fa_xor1(h_s_arrmul16_fa6_2_xor1), .fa_or0(h_s_arrmul16_fa6_2_or0));
  and_gate and_gate_h_s_arrmul16_and7_2(.a(a[7]), .b(b[2]), .out(h_s_arrmul16_and7_2));
  fa fa_h_s_arrmul16_fa7_2_out(.a(h_s_arrmul16_and7_2[0]), .b(h_s_arrmul16_fa8_1_xor1[0]), .cin(h_s_arrmul16_fa6_2_or0[0]), .fa_xor1(h_s_arrmul16_fa7_2_xor1), .fa_or0(h_s_arrmul16_fa7_2_or0));
  and_gate and_gate_h_s_arrmul16_and8_2(.a(a[8]), .b(b[2]), .out(h_s_arrmul16_and8_2));
  fa fa_h_s_arrmul16_fa8_2_out(.a(h_s_arrmul16_and8_2[0]), .b(h_s_arrmul16_fa9_1_xor1[0]), .cin(h_s_arrmul16_fa7_2_or0[0]), .fa_xor1(h_s_arrmul16_fa8_2_xor1), .fa_or0(h_s_arrmul16_fa8_2_or0));
  and_gate and_gate_h_s_arrmul16_and9_2(.a(a[9]), .b(b[2]), .out(h_s_arrmul16_and9_2));
  fa fa_h_s_arrmul16_fa9_2_out(.a(h_s_arrmul16_and9_2[0]), .b(h_s_arrmul16_fa10_1_xor1[0]), .cin(h_s_arrmul16_fa8_2_or0[0]), .fa_xor1(h_s_arrmul16_fa9_2_xor1), .fa_or0(h_s_arrmul16_fa9_2_or0));
  and_gate and_gate_h_s_arrmul16_and10_2(.a(a[10]), .b(b[2]), .out(h_s_arrmul16_and10_2));
  fa fa_h_s_arrmul16_fa10_2_out(.a(h_s_arrmul16_and10_2[0]), .b(h_s_arrmul16_fa11_1_xor1[0]), .cin(h_s_arrmul16_fa9_2_or0[0]), .fa_xor1(h_s_arrmul16_fa10_2_xor1), .fa_or0(h_s_arrmul16_fa10_2_or0));
  and_gate and_gate_h_s_arrmul16_and11_2(.a(a[11]), .b(b[2]), .out(h_s_arrmul16_and11_2));
  fa fa_h_s_arrmul16_fa11_2_out(.a(h_s_arrmul16_and11_2[0]), .b(h_s_arrmul16_fa12_1_xor1[0]), .cin(h_s_arrmul16_fa10_2_or0[0]), .fa_xor1(h_s_arrmul16_fa11_2_xor1), .fa_or0(h_s_arrmul16_fa11_2_or0));
  and_gate and_gate_h_s_arrmul16_and12_2(.a(a[12]), .b(b[2]), .out(h_s_arrmul16_and12_2));
  fa fa_h_s_arrmul16_fa12_2_out(.a(h_s_arrmul16_and12_2[0]), .b(h_s_arrmul16_fa13_1_xor1[0]), .cin(h_s_arrmul16_fa11_2_or0[0]), .fa_xor1(h_s_arrmul16_fa12_2_xor1), .fa_or0(h_s_arrmul16_fa12_2_or0));
  and_gate and_gate_h_s_arrmul16_and13_2(.a(a[13]), .b(b[2]), .out(h_s_arrmul16_and13_2));
  fa fa_h_s_arrmul16_fa13_2_out(.a(h_s_arrmul16_and13_2[0]), .b(h_s_arrmul16_fa14_1_xor1[0]), .cin(h_s_arrmul16_fa12_2_or0[0]), .fa_xor1(h_s_arrmul16_fa13_2_xor1), .fa_or0(h_s_arrmul16_fa13_2_or0));
  and_gate and_gate_h_s_arrmul16_and14_2(.a(a[14]), .b(b[2]), .out(h_s_arrmul16_and14_2));
  fa fa_h_s_arrmul16_fa14_2_out(.a(h_s_arrmul16_and14_2[0]), .b(h_s_arrmul16_fa15_1_xor1[0]), .cin(h_s_arrmul16_fa13_2_or0[0]), .fa_xor1(h_s_arrmul16_fa14_2_xor1), .fa_or0(h_s_arrmul16_fa14_2_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_2(.a(a[15]), .b(b[2]), .out(h_s_arrmul16_nand15_2));
  fa fa_h_s_arrmul16_fa15_2_out(.a(h_s_arrmul16_nand15_2[0]), .b(h_s_arrmul16_fa15_1_or0[0]), .cin(h_s_arrmul16_fa14_2_or0[0]), .fa_xor1(h_s_arrmul16_fa15_2_xor1), .fa_or0(h_s_arrmul16_fa15_2_or0));
  and_gate and_gate_h_s_arrmul16_and0_3(.a(a[0]), .b(b[3]), .out(h_s_arrmul16_and0_3));
  ha ha_h_s_arrmul16_ha0_3_out(.a(h_s_arrmul16_and0_3[0]), .b(h_s_arrmul16_fa1_2_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_3_xor0), .ha_and0(h_s_arrmul16_ha0_3_and0));
  and_gate and_gate_h_s_arrmul16_and1_3(.a(a[1]), .b(b[3]), .out(h_s_arrmul16_and1_3));
  fa fa_h_s_arrmul16_fa1_3_out(.a(h_s_arrmul16_and1_3[0]), .b(h_s_arrmul16_fa2_2_xor1[0]), .cin(h_s_arrmul16_ha0_3_and0[0]), .fa_xor1(h_s_arrmul16_fa1_3_xor1), .fa_or0(h_s_arrmul16_fa1_3_or0));
  and_gate and_gate_h_s_arrmul16_and2_3(.a(a[2]), .b(b[3]), .out(h_s_arrmul16_and2_3));
  fa fa_h_s_arrmul16_fa2_3_out(.a(h_s_arrmul16_and2_3[0]), .b(h_s_arrmul16_fa3_2_xor1[0]), .cin(h_s_arrmul16_fa1_3_or0[0]), .fa_xor1(h_s_arrmul16_fa2_3_xor1), .fa_or0(h_s_arrmul16_fa2_3_or0));
  and_gate and_gate_h_s_arrmul16_and3_3(.a(a[3]), .b(b[3]), .out(h_s_arrmul16_and3_3));
  fa fa_h_s_arrmul16_fa3_3_out(.a(h_s_arrmul16_and3_3[0]), .b(h_s_arrmul16_fa4_2_xor1[0]), .cin(h_s_arrmul16_fa2_3_or0[0]), .fa_xor1(h_s_arrmul16_fa3_3_xor1), .fa_or0(h_s_arrmul16_fa3_3_or0));
  and_gate and_gate_h_s_arrmul16_and4_3(.a(a[4]), .b(b[3]), .out(h_s_arrmul16_and4_3));
  fa fa_h_s_arrmul16_fa4_3_out(.a(h_s_arrmul16_and4_3[0]), .b(h_s_arrmul16_fa5_2_xor1[0]), .cin(h_s_arrmul16_fa3_3_or0[0]), .fa_xor1(h_s_arrmul16_fa4_3_xor1), .fa_or0(h_s_arrmul16_fa4_3_or0));
  and_gate and_gate_h_s_arrmul16_and5_3(.a(a[5]), .b(b[3]), .out(h_s_arrmul16_and5_3));
  fa fa_h_s_arrmul16_fa5_3_out(.a(h_s_arrmul16_and5_3[0]), .b(h_s_arrmul16_fa6_2_xor1[0]), .cin(h_s_arrmul16_fa4_3_or0[0]), .fa_xor1(h_s_arrmul16_fa5_3_xor1), .fa_or0(h_s_arrmul16_fa5_3_or0));
  and_gate and_gate_h_s_arrmul16_and6_3(.a(a[6]), .b(b[3]), .out(h_s_arrmul16_and6_3));
  fa fa_h_s_arrmul16_fa6_3_out(.a(h_s_arrmul16_and6_3[0]), .b(h_s_arrmul16_fa7_2_xor1[0]), .cin(h_s_arrmul16_fa5_3_or0[0]), .fa_xor1(h_s_arrmul16_fa6_3_xor1), .fa_or0(h_s_arrmul16_fa6_3_or0));
  and_gate and_gate_h_s_arrmul16_and7_3(.a(a[7]), .b(b[3]), .out(h_s_arrmul16_and7_3));
  fa fa_h_s_arrmul16_fa7_3_out(.a(h_s_arrmul16_and7_3[0]), .b(h_s_arrmul16_fa8_2_xor1[0]), .cin(h_s_arrmul16_fa6_3_or0[0]), .fa_xor1(h_s_arrmul16_fa7_3_xor1), .fa_or0(h_s_arrmul16_fa7_3_or0));
  and_gate and_gate_h_s_arrmul16_and8_3(.a(a[8]), .b(b[3]), .out(h_s_arrmul16_and8_3));
  fa fa_h_s_arrmul16_fa8_3_out(.a(h_s_arrmul16_and8_3[0]), .b(h_s_arrmul16_fa9_2_xor1[0]), .cin(h_s_arrmul16_fa7_3_or0[0]), .fa_xor1(h_s_arrmul16_fa8_3_xor1), .fa_or0(h_s_arrmul16_fa8_3_or0));
  and_gate and_gate_h_s_arrmul16_and9_3(.a(a[9]), .b(b[3]), .out(h_s_arrmul16_and9_3));
  fa fa_h_s_arrmul16_fa9_3_out(.a(h_s_arrmul16_and9_3[0]), .b(h_s_arrmul16_fa10_2_xor1[0]), .cin(h_s_arrmul16_fa8_3_or0[0]), .fa_xor1(h_s_arrmul16_fa9_3_xor1), .fa_or0(h_s_arrmul16_fa9_3_or0));
  and_gate and_gate_h_s_arrmul16_and10_3(.a(a[10]), .b(b[3]), .out(h_s_arrmul16_and10_3));
  fa fa_h_s_arrmul16_fa10_3_out(.a(h_s_arrmul16_and10_3[0]), .b(h_s_arrmul16_fa11_2_xor1[0]), .cin(h_s_arrmul16_fa9_3_or0[0]), .fa_xor1(h_s_arrmul16_fa10_3_xor1), .fa_or0(h_s_arrmul16_fa10_3_or0));
  and_gate and_gate_h_s_arrmul16_and11_3(.a(a[11]), .b(b[3]), .out(h_s_arrmul16_and11_3));
  fa fa_h_s_arrmul16_fa11_3_out(.a(h_s_arrmul16_and11_3[0]), .b(h_s_arrmul16_fa12_2_xor1[0]), .cin(h_s_arrmul16_fa10_3_or0[0]), .fa_xor1(h_s_arrmul16_fa11_3_xor1), .fa_or0(h_s_arrmul16_fa11_3_or0));
  and_gate and_gate_h_s_arrmul16_and12_3(.a(a[12]), .b(b[3]), .out(h_s_arrmul16_and12_3));
  fa fa_h_s_arrmul16_fa12_3_out(.a(h_s_arrmul16_and12_3[0]), .b(h_s_arrmul16_fa13_2_xor1[0]), .cin(h_s_arrmul16_fa11_3_or0[0]), .fa_xor1(h_s_arrmul16_fa12_3_xor1), .fa_or0(h_s_arrmul16_fa12_3_or0));
  and_gate and_gate_h_s_arrmul16_and13_3(.a(a[13]), .b(b[3]), .out(h_s_arrmul16_and13_3));
  fa fa_h_s_arrmul16_fa13_3_out(.a(h_s_arrmul16_and13_3[0]), .b(h_s_arrmul16_fa14_2_xor1[0]), .cin(h_s_arrmul16_fa12_3_or0[0]), .fa_xor1(h_s_arrmul16_fa13_3_xor1), .fa_or0(h_s_arrmul16_fa13_3_or0));
  and_gate and_gate_h_s_arrmul16_and14_3(.a(a[14]), .b(b[3]), .out(h_s_arrmul16_and14_3));
  fa fa_h_s_arrmul16_fa14_3_out(.a(h_s_arrmul16_and14_3[0]), .b(h_s_arrmul16_fa15_2_xor1[0]), .cin(h_s_arrmul16_fa13_3_or0[0]), .fa_xor1(h_s_arrmul16_fa14_3_xor1), .fa_or0(h_s_arrmul16_fa14_3_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_3(.a(a[15]), .b(b[3]), .out(h_s_arrmul16_nand15_3));
  fa fa_h_s_arrmul16_fa15_3_out(.a(h_s_arrmul16_nand15_3[0]), .b(h_s_arrmul16_fa15_2_or0[0]), .cin(h_s_arrmul16_fa14_3_or0[0]), .fa_xor1(h_s_arrmul16_fa15_3_xor1), .fa_or0(h_s_arrmul16_fa15_3_or0));
  and_gate and_gate_h_s_arrmul16_and0_4(.a(a[0]), .b(b[4]), .out(h_s_arrmul16_and0_4));
  ha ha_h_s_arrmul16_ha0_4_out(.a(h_s_arrmul16_and0_4[0]), .b(h_s_arrmul16_fa1_3_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_4_xor0), .ha_and0(h_s_arrmul16_ha0_4_and0));
  and_gate and_gate_h_s_arrmul16_and1_4(.a(a[1]), .b(b[4]), .out(h_s_arrmul16_and1_4));
  fa fa_h_s_arrmul16_fa1_4_out(.a(h_s_arrmul16_and1_4[0]), .b(h_s_arrmul16_fa2_3_xor1[0]), .cin(h_s_arrmul16_ha0_4_and0[0]), .fa_xor1(h_s_arrmul16_fa1_4_xor1), .fa_or0(h_s_arrmul16_fa1_4_or0));
  and_gate and_gate_h_s_arrmul16_and2_4(.a(a[2]), .b(b[4]), .out(h_s_arrmul16_and2_4));
  fa fa_h_s_arrmul16_fa2_4_out(.a(h_s_arrmul16_and2_4[0]), .b(h_s_arrmul16_fa3_3_xor1[0]), .cin(h_s_arrmul16_fa1_4_or0[0]), .fa_xor1(h_s_arrmul16_fa2_4_xor1), .fa_or0(h_s_arrmul16_fa2_4_or0));
  and_gate and_gate_h_s_arrmul16_and3_4(.a(a[3]), .b(b[4]), .out(h_s_arrmul16_and3_4));
  fa fa_h_s_arrmul16_fa3_4_out(.a(h_s_arrmul16_and3_4[0]), .b(h_s_arrmul16_fa4_3_xor1[0]), .cin(h_s_arrmul16_fa2_4_or0[0]), .fa_xor1(h_s_arrmul16_fa3_4_xor1), .fa_or0(h_s_arrmul16_fa3_4_or0));
  and_gate and_gate_h_s_arrmul16_and4_4(.a(a[4]), .b(b[4]), .out(h_s_arrmul16_and4_4));
  fa fa_h_s_arrmul16_fa4_4_out(.a(h_s_arrmul16_and4_4[0]), .b(h_s_arrmul16_fa5_3_xor1[0]), .cin(h_s_arrmul16_fa3_4_or0[0]), .fa_xor1(h_s_arrmul16_fa4_4_xor1), .fa_or0(h_s_arrmul16_fa4_4_or0));
  and_gate and_gate_h_s_arrmul16_and5_4(.a(a[5]), .b(b[4]), .out(h_s_arrmul16_and5_4));
  fa fa_h_s_arrmul16_fa5_4_out(.a(h_s_arrmul16_and5_4[0]), .b(h_s_arrmul16_fa6_3_xor1[0]), .cin(h_s_arrmul16_fa4_4_or0[0]), .fa_xor1(h_s_arrmul16_fa5_4_xor1), .fa_or0(h_s_arrmul16_fa5_4_or0));
  and_gate and_gate_h_s_arrmul16_and6_4(.a(a[6]), .b(b[4]), .out(h_s_arrmul16_and6_4));
  fa fa_h_s_arrmul16_fa6_4_out(.a(h_s_arrmul16_and6_4[0]), .b(h_s_arrmul16_fa7_3_xor1[0]), .cin(h_s_arrmul16_fa5_4_or0[0]), .fa_xor1(h_s_arrmul16_fa6_4_xor1), .fa_or0(h_s_arrmul16_fa6_4_or0));
  and_gate and_gate_h_s_arrmul16_and7_4(.a(a[7]), .b(b[4]), .out(h_s_arrmul16_and7_4));
  fa fa_h_s_arrmul16_fa7_4_out(.a(h_s_arrmul16_and7_4[0]), .b(h_s_arrmul16_fa8_3_xor1[0]), .cin(h_s_arrmul16_fa6_4_or0[0]), .fa_xor1(h_s_arrmul16_fa7_4_xor1), .fa_or0(h_s_arrmul16_fa7_4_or0));
  and_gate and_gate_h_s_arrmul16_and8_4(.a(a[8]), .b(b[4]), .out(h_s_arrmul16_and8_4));
  fa fa_h_s_arrmul16_fa8_4_out(.a(h_s_arrmul16_and8_4[0]), .b(h_s_arrmul16_fa9_3_xor1[0]), .cin(h_s_arrmul16_fa7_4_or0[0]), .fa_xor1(h_s_arrmul16_fa8_4_xor1), .fa_or0(h_s_arrmul16_fa8_4_or0));
  and_gate and_gate_h_s_arrmul16_and9_4(.a(a[9]), .b(b[4]), .out(h_s_arrmul16_and9_4));
  fa fa_h_s_arrmul16_fa9_4_out(.a(h_s_arrmul16_and9_4[0]), .b(h_s_arrmul16_fa10_3_xor1[0]), .cin(h_s_arrmul16_fa8_4_or0[0]), .fa_xor1(h_s_arrmul16_fa9_4_xor1), .fa_or0(h_s_arrmul16_fa9_4_or0));
  and_gate and_gate_h_s_arrmul16_and10_4(.a(a[10]), .b(b[4]), .out(h_s_arrmul16_and10_4));
  fa fa_h_s_arrmul16_fa10_4_out(.a(h_s_arrmul16_and10_4[0]), .b(h_s_arrmul16_fa11_3_xor1[0]), .cin(h_s_arrmul16_fa9_4_or0[0]), .fa_xor1(h_s_arrmul16_fa10_4_xor1), .fa_or0(h_s_arrmul16_fa10_4_or0));
  and_gate and_gate_h_s_arrmul16_and11_4(.a(a[11]), .b(b[4]), .out(h_s_arrmul16_and11_4));
  fa fa_h_s_arrmul16_fa11_4_out(.a(h_s_arrmul16_and11_4[0]), .b(h_s_arrmul16_fa12_3_xor1[0]), .cin(h_s_arrmul16_fa10_4_or0[0]), .fa_xor1(h_s_arrmul16_fa11_4_xor1), .fa_or0(h_s_arrmul16_fa11_4_or0));
  and_gate and_gate_h_s_arrmul16_and12_4(.a(a[12]), .b(b[4]), .out(h_s_arrmul16_and12_4));
  fa fa_h_s_arrmul16_fa12_4_out(.a(h_s_arrmul16_and12_4[0]), .b(h_s_arrmul16_fa13_3_xor1[0]), .cin(h_s_arrmul16_fa11_4_or0[0]), .fa_xor1(h_s_arrmul16_fa12_4_xor1), .fa_or0(h_s_arrmul16_fa12_4_or0));
  and_gate and_gate_h_s_arrmul16_and13_4(.a(a[13]), .b(b[4]), .out(h_s_arrmul16_and13_4));
  fa fa_h_s_arrmul16_fa13_4_out(.a(h_s_arrmul16_and13_4[0]), .b(h_s_arrmul16_fa14_3_xor1[0]), .cin(h_s_arrmul16_fa12_4_or0[0]), .fa_xor1(h_s_arrmul16_fa13_4_xor1), .fa_or0(h_s_arrmul16_fa13_4_or0));
  and_gate and_gate_h_s_arrmul16_and14_4(.a(a[14]), .b(b[4]), .out(h_s_arrmul16_and14_4));
  fa fa_h_s_arrmul16_fa14_4_out(.a(h_s_arrmul16_and14_4[0]), .b(h_s_arrmul16_fa15_3_xor1[0]), .cin(h_s_arrmul16_fa13_4_or0[0]), .fa_xor1(h_s_arrmul16_fa14_4_xor1), .fa_or0(h_s_arrmul16_fa14_4_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_4(.a(a[15]), .b(b[4]), .out(h_s_arrmul16_nand15_4));
  fa fa_h_s_arrmul16_fa15_4_out(.a(h_s_arrmul16_nand15_4[0]), .b(h_s_arrmul16_fa15_3_or0[0]), .cin(h_s_arrmul16_fa14_4_or0[0]), .fa_xor1(h_s_arrmul16_fa15_4_xor1), .fa_or0(h_s_arrmul16_fa15_4_or0));
  and_gate and_gate_h_s_arrmul16_and0_5(.a(a[0]), .b(b[5]), .out(h_s_arrmul16_and0_5));
  ha ha_h_s_arrmul16_ha0_5_out(.a(h_s_arrmul16_and0_5[0]), .b(h_s_arrmul16_fa1_4_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_5_xor0), .ha_and0(h_s_arrmul16_ha0_5_and0));
  and_gate and_gate_h_s_arrmul16_and1_5(.a(a[1]), .b(b[5]), .out(h_s_arrmul16_and1_5));
  fa fa_h_s_arrmul16_fa1_5_out(.a(h_s_arrmul16_and1_5[0]), .b(h_s_arrmul16_fa2_4_xor1[0]), .cin(h_s_arrmul16_ha0_5_and0[0]), .fa_xor1(h_s_arrmul16_fa1_5_xor1), .fa_or0(h_s_arrmul16_fa1_5_or0));
  and_gate and_gate_h_s_arrmul16_and2_5(.a(a[2]), .b(b[5]), .out(h_s_arrmul16_and2_5));
  fa fa_h_s_arrmul16_fa2_5_out(.a(h_s_arrmul16_and2_5[0]), .b(h_s_arrmul16_fa3_4_xor1[0]), .cin(h_s_arrmul16_fa1_5_or0[0]), .fa_xor1(h_s_arrmul16_fa2_5_xor1), .fa_or0(h_s_arrmul16_fa2_5_or0));
  and_gate and_gate_h_s_arrmul16_and3_5(.a(a[3]), .b(b[5]), .out(h_s_arrmul16_and3_5));
  fa fa_h_s_arrmul16_fa3_5_out(.a(h_s_arrmul16_and3_5[0]), .b(h_s_arrmul16_fa4_4_xor1[0]), .cin(h_s_arrmul16_fa2_5_or0[0]), .fa_xor1(h_s_arrmul16_fa3_5_xor1), .fa_or0(h_s_arrmul16_fa3_5_or0));
  and_gate and_gate_h_s_arrmul16_and4_5(.a(a[4]), .b(b[5]), .out(h_s_arrmul16_and4_5));
  fa fa_h_s_arrmul16_fa4_5_out(.a(h_s_arrmul16_and4_5[0]), .b(h_s_arrmul16_fa5_4_xor1[0]), .cin(h_s_arrmul16_fa3_5_or0[0]), .fa_xor1(h_s_arrmul16_fa4_5_xor1), .fa_or0(h_s_arrmul16_fa4_5_or0));
  and_gate and_gate_h_s_arrmul16_and5_5(.a(a[5]), .b(b[5]), .out(h_s_arrmul16_and5_5));
  fa fa_h_s_arrmul16_fa5_5_out(.a(h_s_arrmul16_and5_5[0]), .b(h_s_arrmul16_fa6_4_xor1[0]), .cin(h_s_arrmul16_fa4_5_or0[0]), .fa_xor1(h_s_arrmul16_fa5_5_xor1), .fa_or0(h_s_arrmul16_fa5_5_or0));
  and_gate and_gate_h_s_arrmul16_and6_5(.a(a[6]), .b(b[5]), .out(h_s_arrmul16_and6_5));
  fa fa_h_s_arrmul16_fa6_5_out(.a(h_s_arrmul16_and6_5[0]), .b(h_s_arrmul16_fa7_4_xor1[0]), .cin(h_s_arrmul16_fa5_5_or0[0]), .fa_xor1(h_s_arrmul16_fa6_5_xor1), .fa_or0(h_s_arrmul16_fa6_5_or0));
  and_gate and_gate_h_s_arrmul16_and7_5(.a(a[7]), .b(b[5]), .out(h_s_arrmul16_and7_5));
  fa fa_h_s_arrmul16_fa7_5_out(.a(h_s_arrmul16_and7_5[0]), .b(h_s_arrmul16_fa8_4_xor1[0]), .cin(h_s_arrmul16_fa6_5_or0[0]), .fa_xor1(h_s_arrmul16_fa7_5_xor1), .fa_or0(h_s_arrmul16_fa7_5_or0));
  and_gate and_gate_h_s_arrmul16_and8_5(.a(a[8]), .b(b[5]), .out(h_s_arrmul16_and8_5));
  fa fa_h_s_arrmul16_fa8_5_out(.a(h_s_arrmul16_and8_5[0]), .b(h_s_arrmul16_fa9_4_xor1[0]), .cin(h_s_arrmul16_fa7_5_or0[0]), .fa_xor1(h_s_arrmul16_fa8_5_xor1), .fa_or0(h_s_arrmul16_fa8_5_or0));
  and_gate and_gate_h_s_arrmul16_and9_5(.a(a[9]), .b(b[5]), .out(h_s_arrmul16_and9_5));
  fa fa_h_s_arrmul16_fa9_5_out(.a(h_s_arrmul16_and9_5[0]), .b(h_s_arrmul16_fa10_4_xor1[0]), .cin(h_s_arrmul16_fa8_5_or0[0]), .fa_xor1(h_s_arrmul16_fa9_5_xor1), .fa_or0(h_s_arrmul16_fa9_5_or0));
  and_gate and_gate_h_s_arrmul16_and10_5(.a(a[10]), .b(b[5]), .out(h_s_arrmul16_and10_5));
  fa fa_h_s_arrmul16_fa10_5_out(.a(h_s_arrmul16_and10_5[0]), .b(h_s_arrmul16_fa11_4_xor1[0]), .cin(h_s_arrmul16_fa9_5_or0[0]), .fa_xor1(h_s_arrmul16_fa10_5_xor1), .fa_or0(h_s_arrmul16_fa10_5_or0));
  and_gate and_gate_h_s_arrmul16_and11_5(.a(a[11]), .b(b[5]), .out(h_s_arrmul16_and11_5));
  fa fa_h_s_arrmul16_fa11_5_out(.a(h_s_arrmul16_and11_5[0]), .b(h_s_arrmul16_fa12_4_xor1[0]), .cin(h_s_arrmul16_fa10_5_or0[0]), .fa_xor1(h_s_arrmul16_fa11_5_xor1), .fa_or0(h_s_arrmul16_fa11_5_or0));
  and_gate and_gate_h_s_arrmul16_and12_5(.a(a[12]), .b(b[5]), .out(h_s_arrmul16_and12_5));
  fa fa_h_s_arrmul16_fa12_5_out(.a(h_s_arrmul16_and12_5[0]), .b(h_s_arrmul16_fa13_4_xor1[0]), .cin(h_s_arrmul16_fa11_5_or0[0]), .fa_xor1(h_s_arrmul16_fa12_5_xor1), .fa_or0(h_s_arrmul16_fa12_5_or0));
  and_gate and_gate_h_s_arrmul16_and13_5(.a(a[13]), .b(b[5]), .out(h_s_arrmul16_and13_5));
  fa fa_h_s_arrmul16_fa13_5_out(.a(h_s_arrmul16_and13_5[0]), .b(h_s_arrmul16_fa14_4_xor1[0]), .cin(h_s_arrmul16_fa12_5_or0[0]), .fa_xor1(h_s_arrmul16_fa13_5_xor1), .fa_or0(h_s_arrmul16_fa13_5_or0));
  and_gate and_gate_h_s_arrmul16_and14_5(.a(a[14]), .b(b[5]), .out(h_s_arrmul16_and14_5));
  fa fa_h_s_arrmul16_fa14_5_out(.a(h_s_arrmul16_and14_5[0]), .b(h_s_arrmul16_fa15_4_xor1[0]), .cin(h_s_arrmul16_fa13_5_or0[0]), .fa_xor1(h_s_arrmul16_fa14_5_xor1), .fa_or0(h_s_arrmul16_fa14_5_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_5(.a(a[15]), .b(b[5]), .out(h_s_arrmul16_nand15_5));
  fa fa_h_s_arrmul16_fa15_5_out(.a(h_s_arrmul16_nand15_5[0]), .b(h_s_arrmul16_fa15_4_or0[0]), .cin(h_s_arrmul16_fa14_5_or0[0]), .fa_xor1(h_s_arrmul16_fa15_5_xor1), .fa_or0(h_s_arrmul16_fa15_5_or0));
  and_gate and_gate_h_s_arrmul16_and0_6(.a(a[0]), .b(b[6]), .out(h_s_arrmul16_and0_6));
  ha ha_h_s_arrmul16_ha0_6_out(.a(h_s_arrmul16_and0_6[0]), .b(h_s_arrmul16_fa1_5_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_6_xor0), .ha_and0(h_s_arrmul16_ha0_6_and0));
  and_gate and_gate_h_s_arrmul16_and1_6(.a(a[1]), .b(b[6]), .out(h_s_arrmul16_and1_6));
  fa fa_h_s_arrmul16_fa1_6_out(.a(h_s_arrmul16_and1_6[0]), .b(h_s_arrmul16_fa2_5_xor1[0]), .cin(h_s_arrmul16_ha0_6_and0[0]), .fa_xor1(h_s_arrmul16_fa1_6_xor1), .fa_or0(h_s_arrmul16_fa1_6_or0));
  and_gate and_gate_h_s_arrmul16_and2_6(.a(a[2]), .b(b[6]), .out(h_s_arrmul16_and2_6));
  fa fa_h_s_arrmul16_fa2_6_out(.a(h_s_arrmul16_and2_6[0]), .b(h_s_arrmul16_fa3_5_xor1[0]), .cin(h_s_arrmul16_fa1_6_or0[0]), .fa_xor1(h_s_arrmul16_fa2_6_xor1), .fa_or0(h_s_arrmul16_fa2_6_or0));
  and_gate and_gate_h_s_arrmul16_and3_6(.a(a[3]), .b(b[6]), .out(h_s_arrmul16_and3_6));
  fa fa_h_s_arrmul16_fa3_6_out(.a(h_s_arrmul16_and3_6[0]), .b(h_s_arrmul16_fa4_5_xor1[0]), .cin(h_s_arrmul16_fa2_6_or0[0]), .fa_xor1(h_s_arrmul16_fa3_6_xor1), .fa_or0(h_s_arrmul16_fa3_6_or0));
  and_gate and_gate_h_s_arrmul16_and4_6(.a(a[4]), .b(b[6]), .out(h_s_arrmul16_and4_6));
  fa fa_h_s_arrmul16_fa4_6_out(.a(h_s_arrmul16_and4_6[0]), .b(h_s_arrmul16_fa5_5_xor1[0]), .cin(h_s_arrmul16_fa3_6_or0[0]), .fa_xor1(h_s_arrmul16_fa4_6_xor1), .fa_or0(h_s_arrmul16_fa4_6_or0));
  and_gate and_gate_h_s_arrmul16_and5_6(.a(a[5]), .b(b[6]), .out(h_s_arrmul16_and5_6));
  fa fa_h_s_arrmul16_fa5_6_out(.a(h_s_arrmul16_and5_6[0]), .b(h_s_arrmul16_fa6_5_xor1[0]), .cin(h_s_arrmul16_fa4_6_or0[0]), .fa_xor1(h_s_arrmul16_fa5_6_xor1), .fa_or0(h_s_arrmul16_fa5_6_or0));
  and_gate and_gate_h_s_arrmul16_and6_6(.a(a[6]), .b(b[6]), .out(h_s_arrmul16_and6_6));
  fa fa_h_s_arrmul16_fa6_6_out(.a(h_s_arrmul16_and6_6[0]), .b(h_s_arrmul16_fa7_5_xor1[0]), .cin(h_s_arrmul16_fa5_6_or0[0]), .fa_xor1(h_s_arrmul16_fa6_6_xor1), .fa_or0(h_s_arrmul16_fa6_6_or0));
  and_gate and_gate_h_s_arrmul16_and7_6(.a(a[7]), .b(b[6]), .out(h_s_arrmul16_and7_6));
  fa fa_h_s_arrmul16_fa7_6_out(.a(h_s_arrmul16_and7_6[0]), .b(h_s_arrmul16_fa8_5_xor1[0]), .cin(h_s_arrmul16_fa6_6_or0[0]), .fa_xor1(h_s_arrmul16_fa7_6_xor1), .fa_or0(h_s_arrmul16_fa7_6_or0));
  and_gate and_gate_h_s_arrmul16_and8_6(.a(a[8]), .b(b[6]), .out(h_s_arrmul16_and8_6));
  fa fa_h_s_arrmul16_fa8_6_out(.a(h_s_arrmul16_and8_6[0]), .b(h_s_arrmul16_fa9_5_xor1[0]), .cin(h_s_arrmul16_fa7_6_or0[0]), .fa_xor1(h_s_arrmul16_fa8_6_xor1), .fa_or0(h_s_arrmul16_fa8_6_or0));
  and_gate and_gate_h_s_arrmul16_and9_6(.a(a[9]), .b(b[6]), .out(h_s_arrmul16_and9_6));
  fa fa_h_s_arrmul16_fa9_6_out(.a(h_s_arrmul16_and9_6[0]), .b(h_s_arrmul16_fa10_5_xor1[0]), .cin(h_s_arrmul16_fa8_6_or0[0]), .fa_xor1(h_s_arrmul16_fa9_6_xor1), .fa_or0(h_s_arrmul16_fa9_6_or0));
  and_gate and_gate_h_s_arrmul16_and10_6(.a(a[10]), .b(b[6]), .out(h_s_arrmul16_and10_6));
  fa fa_h_s_arrmul16_fa10_6_out(.a(h_s_arrmul16_and10_6[0]), .b(h_s_arrmul16_fa11_5_xor1[0]), .cin(h_s_arrmul16_fa9_6_or0[0]), .fa_xor1(h_s_arrmul16_fa10_6_xor1), .fa_or0(h_s_arrmul16_fa10_6_or0));
  and_gate and_gate_h_s_arrmul16_and11_6(.a(a[11]), .b(b[6]), .out(h_s_arrmul16_and11_6));
  fa fa_h_s_arrmul16_fa11_6_out(.a(h_s_arrmul16_and11_6[0]), .b(h_s_arrmul16_fa12_5_xor1[0]), .cin(h_s_arrmul16_fa10_6_or0[0]), .fa_xor1(h_s_arrmul16_fa11_6_xor1), .fa_or0(h_s_arrmul16_fa11_6_or0));
  and_gate and_gate_h_s_arrmul16_and12_6(.a(a[12]), .b(b[6]), .out(h_s_arrmul16_and12_6));
  fa fa_h_s_arrmul16_fa12_6_out(.a(h_s_arrmul16_and12_6[0]), .b(h_s_arrmul16_fa13_5_xor1[0]), .cin(h_s_arrmul16_fa11_6_or0[0]), .fa_xor1(h_s_arrmul16_fa12_6_xor1), .fa_or0(h_s_arrmul16_fa12_6_or0));
  and_gate and_gate_h_s_arrmul16_and13_6(.a(a[13]), .b(b[6]), .out(h_s_arrmul16_and13_6));
  fa fa_h_s_arrmul16_fa13_6_out(.a(h_s_arrmul16_and13_6[0]), .b(h_s_arrmul16_fa14_5_xor1[0]), .cin(h_s_arrmul16_fa12_6_or0[0]), .fa_xor1(h_s_arrmul16_fa13_6_xor1), .fa_or0(h_s_arrmul16_fa13_6_or0));
  and_gate and_gate_h_s_arrmul16_and14_6(.a(a[14]), .b(b[6]), .out(h_s_arrmul16_and14_6));
  fa fa_h_s_arrmul16_fa14_6_out(.a(h_s_arrmul16_and14_6[0]), .b(h_s_arrmul16_fa15_5_xor1[0]), .cin(h_s_arrmul16_fa13_6_or0[0]), .fa_xor1(h_s_arrmul16_fa14_6_xor1), .fa_or0(h_s_arrmul16_fa14_6_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_6(.a(a[15]), .b(b[6]), .out(h_s_arrmul16_nand15_6));
  fa fa_h_s_arrmul16_fa15_6_out(.a(h_s_arrmul16_nand15_6[0]), .b(h_s_arrmul16_fa15_5_or0[0]), .cin(h_s_arrmul16_fa14_6_or0[0]), .fa_xor1(h_s_arrmul16_fa15_6_xor1), .fa_or0(h_s_arrmul16_fa15_6_or0));
  and_gate and_gate_h_s_arrmul16_and0_7(.a(a[0]), .b(b[7]), .out(h_s_arrmul16_and0_7));
  ha ha_h_s_arrmul16_ha0_7_out(.a(h_s_arrmul16_and0_7[0]), .b(h_s_arrmul16_fa1_6_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_7_xor0), .ha_and0(h_s_arrmul16_ha0_7_and0));
  and_gate and_gate_h_s_arrmul16_and1_7(.a(a[1]), .b(b[7]), .out(h_s_arrmul16_and1_7));
  fa fa_h_s_arrmul16_fa1_7_out(.a(h_s_arrmul16_and1_7[0]), .b(h_s_arrmul16_fa2_6_xor1[0]), .cin(h_s_arrmul16_ha0_7_and0[0]), .fa_xor1(h_s_arrmul16_fa1_7_xor1), .fa_or0(h_s_arrmul16_fa1_7_or0));
  and_gate and_gate_h_s_arrmul16_and2_7(.a(a[2]), .b(b[7]), .out(h_s_arrmul16_and2_7));
  fa fa_h_s_arrmul16_fa2_7_out(.a(h_s_arrmul16_and2_7[0]), .b(h_s_arrmul16_fa3_6_xor1[0]), .cin(h_s_arrmul16_fa1_7_or0[0]), .fa_xor1(h_s_arrmul16_fa2_7_xor1), .fa_or0(h_s_arrmul16_fa2_7_or0));
  and_gate and_gate_h_s_arrmul16_and3_7(.a(a[3]), .b(b[7]), .out(h_s_arrmul16_and3_7));
  fa fa_h_s_arrmul16_fa3_7_out(.a(h_s_arrmul16_and3_7[0]), .b(h_s_arrmul16_fa4_6_xor1[0]), .cin(h_s_arrmul16_fa2_7_or0[0]), .fa_xor1(h_s_arrmul16_fa3_7_xor1), .fa_or0(h_s_arrmul16_fa3_7_or0));
  and_gate and_gate_h_s_arrmul16_and4_7(.a(a[4]), .b(b[7]), .out(h_s_arrmul16_and4_7));
  fa fa_h_s_arrmul16_fa4_7_out(.a(h_s_arrmul16_and4_7[0]), .b(h_s_arrmul16_fa5_6_xor1[0]), .cin(h_s_arrmul16_fa3_7_or0[0]), .fa_xor1(h_s_arrmul16_fa4_7_xor1), .fa_or0(h_s_arrmul16_fa4_7_or0));
  and_gate and_gate_h_s_arrmul16_and5_7(.a(a[5]), .b(b[7]), .out(h_s_arrmul16_and5_7));
  fa fa_h_s_arrmul16_fa5_7_out(.a(h_s_arrmul16_and5_7[0]), .b(h_s_arrmul16_fa6_6_xor1[0]), .cin(h_s_arrmul16_fa4_7_or0[0]), .fa_xor1(h_s_arrmul16_fa5_7_xor1), .fa_or0(h_s_arrmul16_fa5_7_or0));
  and_gate and_gate_h_s_arrmul16_and6_7(.a(a[6]), .b(b[7]), .out(h_s_arrmul16_and6_7));
  fa fa_h_s_arrmul16_fa6_7_out(.a(h_s_arrmul16_and6_7[0]), .b(h_s_arrmul16_fa7_6_xor1[0]), .cin(h_s_arrmul16_fa5_7_or0[0]), .fa_xor1(h_s_arrmul16_fa6_7_xor1), .fa_or0(h_s_arrmul16_fa6_7_or0));
  and_gate and_gate_h_s_arrmul16_and7_7(.a(a[7]), .b(b[7]), .out(h_s_arrmul16_and7_7));
  fa fa_h_s_arrmul16_fa7_7_out(.a(h_s_arrmul16_and7_7[0]), .b(h_s_arrmul16_fa8_6_xor1[0]), .cin(h_s_arrmul16_fa6_7_or0[0]), .fa_xor1(h_s_arrmul16_fa7_7_xor1), .fa_or0(h_s_arrmul16_fa7_7_or0));
  and_gate and_gate_h_s_arrmul16_and8_7(.a(a[8]), .b(b[7]), .out(h_s_arrmul16_and8_7));
  fa fa_h_s_arrmul16_fa8_7_out(.a(h_s_arrmul16_and8_7[0]), .b(h_s_arrmul16_fa9_6_xor1[0]), .cin(h_s_arrmul16_fa7_7_or0[0]), .fa_xor1(h_s_arrmul16_fa8_7_xor1), .fa_or0(h_s_arrmul16_fa8_7_or0));
  and_gate and_gate_h_s_arrmul16_and9_7(.a(a[9]), .b(b[7]), .out(h_s_arrmul16_and9_7));
  fa fa_h_s_arrmul16_fa9_7_out(.a(h_s_arrmul16_and9_7[0]), .b(h_s_arrmul16_fa10_6_xor1[0]), .cin(h_s_arrmul16_fa8_7_or0[0]), .fa_xor1(h_s_arrmul16_fa9_7_xor1), .fa_or0(h_s_arrmul16_fa9_7_or0));
  and_gate and_gate_h_s_arrmul16_and10_7(.a(a[10]), .b(b[7]), .out(h_s_arrmul16_and10_7));
  fa fa_h_s_arrmul16_fa10_7_out(.a(h_s_arrmul16_and10_7[0]), .b(h_s_arrmul16_fa11_6_xor1[0]), .cin(h_s_arrmul16_fa9_7_or0[0]), .fa_xor1(h_s_arrmul16_fa10_7_xor1), .fa_or0(h_s_arrmul16_fa10_7_or0));
  and_gate and_gate_h_s_arrmul16_and11_7(.a(a[11]), .b(b[7]), .out(h_s_arrmul16_and11_7));
  fa fa_h_s_arrmul16_fa11_7_out(.a(h_s_arrmul16_and11_7[0]), .b(h_s_arrmul16_fa12_6_xor1[0]), .cin(h_s_arrmul16_fa10_7_or0[0]), .fa_xor1(h_s_arrmul16_fa11_7_xor1), .fa_or0(h_s_arrmul16_fa11_7_or0));
  and_gate and_gate_h_s_arrmul16_and12_7(.a(a[12]), .b(b[7]), .out(h_s_arrmul16_and12_7));
  fa fa_h_s_arrmul16_fa12_7_out(.a(h_s_arrmul16_and12_7[0]), .b(h_s_arrmul16_fa13_6_xor1[0]), .cin(h_s_arrmul16_fa11_7_or0[0]), .fa_xor1(h_s_arrmul16_fa12_7_xor1), .fa_or0(h_s_arrmul16_fa12_7_or0));
  and_gate and_gate_h_s_arrmul16_and13_7(.a(a[13]), .b(b[7]), .out(h_s_arrmul16_and13_7));
  fa fa_h_s_arrmul16_fa13_7_out(.a(h_s_arrmul16_and13_7[0]), .b(h_s_arrmul16_fa14_6_xor1[0]), .cin(h_s_arrmul16_fa12_7_or0[0]), .fa_xor1(h_s_arrmul16_fa13_7_xor1), .fa_or0(h_s_arrmul16_fa13_7_or0));
  and_gate and_gate_h_s_arrmul16_and14_7(.a(a[14]), .b(b[7]), .out(h_s_arrmul16_and14_7));
  fa fa_h_s_arrmul16_fa14_7_out(.a(h_s_arrmul16_and14_7[0]), .b(h_s_arrmul16_fa15_6_xor1[0]), .cin(h_s_arrmul16_fa13_7_or0[0]), .fa_xor1(h_s_arrmul16_fa14_7_xor1), .fa_or0(h_s_arrmul16_fa14_7_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_7(.a(a[15]), .b(b[7]), .out(h_s_arrmul16_nand15_7));
  fa fa_h_s_arrmul16_fa15_7_out(.a(h_s_arrmul16_nand15_7[0]), .b(h_s_arrmul16_fa15_6_or0[0]), .cin(h_s_arrmul16_fa14_7_or0[0]), .fa_xor1(h_s_arrmul16_fa15_7_xor1), .fa_or0(h_s_arrmul16_fa15_7_or0));
  and_gate and_gate_h_s_arrmul16_and0_8(.a(a[0]), .b(b[8]), .out(h_s_arrmul16_and0_8));
  ha ha_h_s_arrmul16_ha0_8_out(.a(h_s_arrmul16_and0_8[0]), .b(h_s_arrmul16_fa1_7_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_8_xor0), .ha_and0(h_s_arrmul16_ha0_8_and0));
  and_gate and_gate_h_s_arrmul16_and1_8(.a(a[1]), .b(b[8]), .out(h_s_arrmul16_and1_8));
  fa fa_h_s_arrmul16_fa1_8_out(.a(h_s_arrmul16_and1_8[0]), .b(h_s_arrmul16_fa2_7_xor1[0]), .cin(h_s_arrmul16_ha0_8_and0[0]), .fa_xor1(h_s_arrmul16_fa1_8_xor1), .fa_or0(h_s_arrmul16_fa1_8_or0));
  and_gate and_gate_h_s_arrmul16_and2_8(.a(a[2]), .b(b[8]), .out(h_s_arrmul16_and2_8));
  fa fa_h_s_arrmul16_fa2_8_out(.a(h_s_arrmul16_and2_8[0]), .b(h_s_arrmul16_fa3_7_xor1[0]), .cin(h_s_arrmul16_fa1_8_or0[0]), .fa_xor1(h_s_arrmul16_fa2_8_xor1), .fa_or0(h_s_arrmul16_fa2_8_or0));
  and_gate and_gate_h_s_arrmul16_and3_8(.a(a[3]), .b(b[8]), .out(h_s_arrmul16_and3_8));
  fa fa_h_s_arrmul16_fa3_8_out(.a(h_s_arrmul16_and3_8[0]), .b(h_s_arrmul16_fa4_7_xor1[0]), .cin(h_s_arrmul16_fa2_8_or0[0]), .fa_xor1(h_s_arrmul16_fa3_8_xor1), .fa_or0(h_s_arrmul16_fa3_8_or0));
  and_gate and_gate_h_s_arrmul16_and4_8(.a(a[4]), .b(b[8]), .out(h_s_arrmul16_and4_8));
  fa fa_h_s_arrmul16_fa4_8_out(.a(h_s_arrmul16_and4_8[0]), .b(h_s_arrmul16_fa5_7_xor1[0]), .cin(h_s_arrmul16_fa3_8_or0[0]), .fa_xor1(h_s_arrmul16_fa4_8_xor1), .fa_or0(h_s_arrmul16_fa4_8_or0));
  and_gate and_gate_h_s_arrmul16_and5_8(.a(a[5]), .b(b[8]), .out(h_s_arrmul16_and5_8));
  fa fa_h_s_arrmul16_fa5_8_out(.a(h_s_arrmul16_and5_8[0]), .b(h_s_arrmul16_fa6_7_xor1[0]), .cin(h_s_arrmul16_fa4_8_or0[0]), .fa_xor1(h_s_arrmul16_fa5_8_xor1), .fa_or0(h_s_arrmul16_fa5_8_or0));
  and_gate and_gate_h_s_arrmul16_and6_8(.a(a[6]), .b(b[8]), .out(h_s_arrmul16_and6_8));
  fa fa_h_s_arrmul16_fa6_8_out(.a(h_s_arrmul16_and6_8[0]), .b(h_s_arrmul16_fa7_7_xor1[0]), .cin(h_s_arrmul16_fa5_8_or0[0]), .fa_xor1(h_s_arrmul16_fa6_8_xor1), .fa_or0(h_s_arrmul16_fa6_8_or0));
  and_gate and_gate_h_s_arrmul16_and7_8(.a(a[7]), .b(b[8]), .out(h_s_arrmul16_and7_8));
  fa fa_h_s_arrmul16_fa7_8_out(.a(h_s_arrmul16_and7_8[0]), .b(h_s_arrmul16_fa8_7_xor1[0]), .cin(h_s_arrmul16_fa6_8_or0[0]), .fa_xor1(h_s_arrmul16_fa7_8_xor1), .fa_or0(h_s_arrmul16_fa7_8_or0));
  and_gate and_gate_h_s_arrmul16_and8_8(.a(a[8]), .b(b[8]), .out(h_s_arrmul16_and8_8));
  fa fa_h_s_arrmul16_fa8_8_out(.a(h_s_arrmul16_and8_8[0]), .b(h_s_arrmul16_fa9_7_xor1[0]), .cin(h_s_arrmul16_fa7_8_or0[0]), .fa_xor1(h_s_arrmul16_fa8_8_xor1), .fa_or0(h_s_arrmul16_fa8_8_or0));
  and_gate and_gate_h_s_arrmul16_and9_8(.a(a[9]), .b(b[8]), .out(h_s_arrmul16_and9_8));
  fa fa_h_s_arrmul16_fa9_8_out(.a(h_s_arrmul16_and9_8[0]), .b(h_s_arrmul16_fa10_7_xor1[0]), .cin(h_s_arrmul16_fa8_8_or0[0]), .fa_xor1(h_s_arrmul16_fa9_8_xor1), .fa_or0(h_s_arrmul16_fa9_8_or0));
  and_gate and_gate_h_s_arrmul16_and10_8(.a(a[10]), .b(b[8]), .out(h_s_arrmul16_and10_8));
  fa fa_h_s_arrmul16_fa10_8_out(.a(h_s_arrmul16_and10_8[0]), .b(h_s_arrmul16_fa11_7_xor1[0]), .cin(h_s_arrmul16_fa9_8_or0[0]), .fa_xor1(h_s_arrmul16_fa10_8_xor1), .fa_or0(h_s_arrmul16_fa10_8_or0));
  and_gate and_gate_h_s_arrmul16_and11_8(.a(a[11]), .b(b[8]), .out(h_s_arrmul16_and11_8));
  fa fa_h_s_arrmul16_fa11_8_out(.a(h_s_arrmul16_and11_8[0]), .b(h_s_arrmul16_fa12_7_xor1[0]), .cin(h_s_arrmul16_fa10_8_or0[0]), .fa_xor1(h_s_arrmul16_fa11_8_xor1), .fa_or0(h_s_arrmul16_fa11_8_or0));
  and_gate and_gate_h_s_arrmul16_and12_8(.a(a[12]), .b(b[8]), .out(h_s_arrmul16_and12_8));
  fa fa_h_s_arrmul16_fa12_8_out(.a(h_s_arrmul16_and12_8[0]), .b(h_s_arrmul16_fa13_7_xor1[0]), .cin(h_s_arrmul16_fa11_8_or0[0]), .fa_xor1(h_s_arrmul16_fa12_8_xor1), .fa_or0(h_s_arrmul16_fa12_8_or0));
  and_gate and_gate_h_s_arrmul16_and13_8(.a(a[13]), .b(b[8]), .out(h_s_arrmul16_and13_8));
  fa fa_h_s_arrmul16_fa13_8_out(.a(h_s_arrmul16_and13_8[0]), .b(h_s_arrmul16_fa14_7_xor1[0]), .cin(h_s_arrmul16_fa12_8_or0[0]), .fa_xor1(h_s_arrmul16_fa13_8_xor1), .fa_or0(h_s_arrmul16_fa13_8_or0));
  and_gate and_gate_h_s_arrmul16_and14_8(.a(a[14]), .b(b[8]), .out(h_s_arrmul16_and14_8));
  fa fa_h_s_arrmul16_fa14_8_out(.a(h_s_arrmul16_and14_8[0]), .b(h_s_arrmul16_fa15_7_xor1[0]), .cin(h_s_arrmul16_fa13_8_or0[0]), .fa_xor1(h_s_arrmul16_fa14_8_xor1), .fa_or0(h_s_arrmul16_fa14_8_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_8(.a(a[15]), .b(b[8]), .out(h_s_arrmul16_nand15_8));
  fa fa_h_s_arrmul16_fa15_8_out(.a(h_s_arrmul16_nand15_8[0]), .b(h_s_arrmul16_fa15_7_or0[0]), .cin(h_s_arrmul16_fa14_8_or0[0]), .fa_xor1(h_s_arrmul16_fa15_8_xor1), .fa_or0(h_s_arrmul16_fa15_8_or0));
  and_gate and_gate_h_s_arrmul16_and0_9(.a(a[0]), .b(b[9]), .out(h_s_arrmul16_and0_9));
  ha ha_h_s_arrmul16_ha0_9_out(.a(h_s_arrmul16_and0_9[0]), .b(h_s_arrmul16_fa1_8_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_9_xor0), .ha_and0(h_s_arrmul16_ha0_9_and0));
  and_gate and_gate_h_s_arrmul16_and1_9(.a(a[1]), .b(b[9]), .out(h_s_arrmul16_and1_9));
  fa fa_h_s_arrmul16_fa1_9_out(.a(h_s_arrmul16_and1_9[0]), .b(h_s_arrmul16_fa2_8_xor1[0]), .cin(h_s_arrmul16_ha0_9_and0[0]), .fa_xor1(h_s_arrmul16_fa1_9_xor1), .fa_or0(h_s_arrmul16_fa1_9_or0));
  and_gate and_gate_h_s_arrmul16_and2_9(.a(a[2]), .b(b[9]), .out(h_s_arrmul16_and2_9));
  fa fa_h_s_arrmul16_fa2_9_out(.a(h_s_arrmul16_and2_9[0]), .b(h_s_arrmul16_fa3_8_xor1[0]), .cin(h_s_arrmul16_fa1_9_or0[0]), .fa_xor1(h_s_arrmul16_fa2_9_xor1), .fa_or0(h_s_arrmul16_fa2_9_or0));
  and_gate and_gate_h_s_arrmul16_and3_9(.a(a[3]), .b(b[9]), .out(h_s_arrmul16_and3_9));
  fa fa_h_s_arrmul16_fa3_9_out(.a(h_s_arrmul16_and3_9[0]), .b(h_s_arrmul16_fa4_8_xor1[0]), .cin(h_s_arrmul16_fa2_9_or0[0]), .fa_xor1(h_s_arrmul16_fa3_9_xor1), .fa_or0(h_s_arrmul16_fa3_9_or0));
  and_gate and_gate_h_s_arrmul16_and4_9(.a(a[4]), .b(b[9]), .out(h_s_arrmul16_and4_9));
  fa fa_h_s_arrmul16_fa4_9_out(.a(h_s_arrmul16_and4_9[0]), .b(h_s_arrmul16_fa5_8_xor1[0]), .cin(h_s_arrmul16_fa3_9_or0[0]), .fa_xor1(h_s_arrmul16_fa4_9_xor1), .fa_or0(h_s_arrmul16_fa4_9_or0));
  and_gate and_gate_h_s_arrmul16_and5_9(.a(a[5]), .b(b[9]), .out(h_s_arrmul16_and5_9));
  fa fa_h_s_arrmul16_fa5_9_out(.a(h_s_arrmul16_and5_9[0]), .b(h_s_arrmul16_fa6_8_xor1[0]), .cin(h_s_arrmul16_fa4_9_or0[0]), .fa_xor1(h_s_arrmul16_fa5_9_xor1), .fa_or0(h_s_arrmul16_fa5_9_or0));
  and_gate and_gate_h_s_arrmul16_and6_9(.a(a[6]), .b(b[9]), .out(h_s_arrmul16_and6_9));
  fa fa_h_s_arrmul16_fa6_9_out(.a(h_s_arrmul16_and6_9[0]), .b(h_s_arrmul16_fa7_8_xor1[0]), .cin(h_s_arrmul16_fa5_9_or0[0]), .fa_xor1(h_s_arrmul16_fa6_9_xor1), .fa_or0(h_s_arrmul16_fa6_9_or0));
  and_gate and_gate_h_s_arrmul16_and7_9(.a(a[7]), .b(b[9]), .out(h_s_arrmul16_and7_9));
  fa fa_h_s_arrmul16_fa7_9_out(.a(h_s_arrmul16_and7_9[0]), .b(h_s_arrmul16_fa8_8_xor1[0]), .cin(h_s_arrmul16_fa6_9_or0[0]), .fa_xor1(h_s_arrmul16_fa7_9_xor1), .fa_or0(h_s_arrmul16_fa7_9_or0));
  and_gate and_gate_h_s_arrmul16_and8_9(.a(a[8]), .b(b[9]), .out(h_s_arrmul16_and8_9));
  fa fa_h_s_arrmul16_fa8_9_out(.a(h_s_arrmul16_and8_9[0]), .b(h_s_arrmul16_fa9_8_xor1[0]), .cin(h_s_arrmul16_fa7_9_or0[0]), .fa_xor1(h_s_arrmul16_fa8_9_xor1), .fa_or0(h_s_arrmul16_fa8_9_or0));
  and_gate and_gate_h_s_arrmul16_and9_9(.a(a[9]), .b(b[9]), .out(h_s_arrmul16_and9_9));
  fa fa_h_s_arrmul16_fa9_9_out(.a(h_s_arrmul16_and9_9[0]), .b(h_s_arrmul16_fa10_8_xor1[0]), .cin(h_s_arrmul16_fa8_9_or0[0]), .fa_xor1(h_s_arrmul16_fa9_9_xor1), .fa_or0(h_s_arrmul16_fa9_9_or0));
  and_gate and_gate_h_s_arrmul16_and10_9(.a(a[10]), .b(b[9]), .out(h_s_arrmul16_and10_9));
  fa fa_h_s_arrmul16_fa10_9_out(.a(h_s_arrmul16_and10_9[0]), .b(h_s_arrmul16_fa11_8_xor1[0]), .cin(h_s_arrmul16_fa9_9_or0[0]), .fa_xor1(h_s_arrmul16_fa10_9_xor1), .fa_or0(h_s_arrmul16_fa10_9_or0));
  and_gate and_gate_h_s_arrmul16_and11_9(.a(a[11]), .b(b[9]), .out(h_s_arrmul16_and11_9));
  fa fa_h_s_arrmul16_fa11_9_out(.a(h_s_arrmul16_and11_9[0]), .b(h_s_arrmul16_fa12_8_xor1[0]), .cin(h_s_arrmul16_fa10_9_or0[0]), .fa_xor1(h_s_arrmul16_fa11_9_xor1), .fa_or0(h_s_arrmul16_fa11_9_or0));
  and_gate and_gate_h_s_arrmul16_and12_9(.a(a[12]), .b(b[9]), .out(h_s_arrmul16_and12_9));
  fa fa_h_s_arrmul16_fa12_9_out(.a(h_s_arrmul16_and12_9[0]), .b(h_s_arrmul16_fa13_8_xor1[0]), .cin(h_s_arrmul16_fa11_9_or0[0]), .fa_xor1(h_s_arrmul16_fa12_9_xor1), .fa_or0(h_s_arrmul16_fa12_9_or0));
  and_gate and_gate_h_s_arrmul16_and13_9(.a(a[13]), .b(b[9]), .out(h_s_arrmul16_and13_9));
  fa fa_h_s_arrmul16_fa13_9_out(.a(h_s_arrmul16_and13_9[0]), .b(h_s_arrmul16_fa14_8_xor1[0]), .cin(h_s_arrmul16_fa12_9_or0[0]), .fa_xor1(h_s_arrmul16_fa13_9_xor1), .fa_or0(h_s_arrmul16_fa13_9_or0));
  and_gate and_gate_h_s_arrmul16_and14_9(.a(a[14]), .b(b[9]), .out(h_s_arrmul16_and14_9));
  fa fa_h_s_arrmul16_fa14_9_out(.a(h_s_arrmul16_and14_9[0]), .b(h_s_arrmul16_fa15_8_xor1[0]), .cin(h_s_arrmul16_fa13_9_or0[0]), .fa_xor1(h_s_arrmul16_fa14_9_xor1), .fa_or0(h_s_arrmul16_fa14_9_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_9(.a(a[15]), .b(b[9]), .out(h_s_arrmul16_nand15_9));
  fa fa_h_s_arrmul16_fa15_9_out(.a(h_s_arrmul16_nand15_9[0]), .b(h_s_arrmul16_fa15_8_or0[0]), .cin(h_s_arrmul16_fa14_9_or0[0]), .fa_xor1(h_s_arrmul16_fa15_9_xor1), .fa_or0(h_s_arrmul16_fa15_9_or0));
  and_gate and_gate_h_s_arrmul16_and0_10(.a(a[0]), .b(b[10]), .out(h_s_arrmul16_and0_10));
  ha ha_h_s_arrmul16_ha0_10_out(.a(h_s_arrmul16_and0_10[0]), .b(h_s_arrmul16_fa1_9_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_10_xor0), .ha_and0(h_s_arrmul16_ha0_10_and0));
  and_gate and_gate_h_s_arrmul16_and1_10(.a(a[1]), .b(b[10]), .out(h_s_arrmul16_and1_10));
  fa fa_h_s_arrmul16_fa1_10_out(.a(h_s_arrmul16_and1_10[0]), .b(h_s_arrmul16_fa2_9_xor1[0]), .cin(h_s_arrmul16_ha0_10_and0[0]), .fa_xor1(h_s_arrmul16_fa1_10_xor1), .fa_or0(h_s_arrmul16_fa1_10_or0));
  and_gate and_gate_h_s_arrmul16_and2_10(.a(a[2]), .b(b[10]), .out(h_s_arrmul16_and2_10));
  fa fa_h_s_arrmul16_fa2_10_out(.a(h_s_arrmul16_and2_10[0]), .b(h_s_arrmul16_fa3_9_xor1[0]), .cin(h_s_arrmul16_fa1_10_or0[0]), .fa_xor1(h_s_arrmul16_fa2_10_xor1), .fa_or0(h_s_arrmul16_fa2_10_or0));
  and_gate and_gate_h_s_arrmul16_and3_10(.a(a[3]), .b(b[10]), .out(h_s_arrmul16_and3_10));
  fa fa_h_s_arrmul16_fa3_10_out(.a(h_s_arrmul16_and3_10[0]), .b(h_s_arrmul16_fa4_9_xor1[0]), .cin(h_s_arrmul16_fa2_10_or0[0]), .fa_xor1(h_s_arrmul16_fa3_10_xor1), .fa_or0(h_s_arrmul16_fa3_10_or0));
  and_gate and_gate_h_s_arrmul16_and4_10(.a(a[4]), .b(b[10]), .out(h_s_arrmul16_and4_10));
  fa fa_h_s_arrmul16_fa4_10_out(.a(h_s_arrmul16_and4_10[0]), .b(h_s_arrmul16_fa5_9_xor1[0]), .cin(h_s_arrmul16_fa3_10_or0[0]), .fa_xor1(h_s_arrmul16_fa4_10_xor1), .fa_or0(h_s_arrmul16_fa4_10_or0));
  and_gate and_gate_h_s_arrmul16_and5_10(.a(a[5]), .b(b[10]), .out(h_s_arrmul16_and5_10));
  fa fa_h_s_arrmul16_fa5_10_out(.a(h_s_arrmul16_and5_10[0]), .b(h_s_arrmul16_fa6_9_xor1[0]), .cin(h_s_arrmul16_fa4_10_or0[0]), .fa_xor1(h_s_arrmul16_fa5_10_xor1), .fa_or0(h_s_arrmul16_fa5_10_or0));
  and_gate and_gate_h_s_arrmul16_and6_10(.a(a[6]), .b(b[10]), .out(h_s_arrmul16_and6_10));
  fa fa_h_s_arrmul16_fa6_10_out(.a(h_s_arrmul16_and6_10[0]), .b(h_s_arrmul16_fa7_9_xor1[0]), .cin(h_s_arrmul16_fa5_10_or0[0]), .fa_xor1(h_s_arrmul16_fa6_10_xor1), .fa_or0(h_s_arrmul16_fa6_10_or0));
  and_gate and_gate_h_s_arrmul16_and7_10(.a(a[7]), .b(b[10]), .out(h_s_arrmul16_and7_10));
  fa fa_h_s_arrmul16_fa7_10_out(.a(h_s_arrmul16_and7_10[0]), .b(h_s_arrmul16_fa8_9_xor1[0]), .cin(h_s_arrmul16_fa6_10_or0[0]), .fa_xor1(h_s_arrmul16_fa7_10_xor1), .fa_or0(h_s_arrmul16_fa7_10_or0));
  and_gate and_gate_h_s_arrmul16_and8_10(.a(a[8]), .b(b[10]), .out(h_s_arrmul16_and8_10));
  fa fa_h_s_arrmul16_fa8_10_out(.a(h_s_arrmul16_and8_10[0]), .b(h_s_arrmul16_fa9_9_xor1[0]), .cin(h_s_arrmul16_fa7_10_or0[0]), .fa_xor1(h_s_arrmul16_fa8_10_xor1), .fa_or0(h_s_arrmul16_fa8_10_or0));
  and_gate and_gate_h_s_arrmul16_and9_10(.a(a[9]), .b(b[10]), .out(h_s_arrmul16_and9_10));
  fa fa_h_s_arrmul16_fa9_10_out(.a(h_s_arrmul16_and9_10[0]), .b(h_s_arrmul16_fa10_9_xor1[0]), .cin(h_s_arrmul16_fa8_10_or0[0]), .fa_xor1(h_s_arrmul16_fa9_10_xor1), .fa_or0(h_s_arrmul16_fa9_10_or0));
  and_gate and_gate_h_s_arrmul16_and10_10(.a(a[10]), .b(b[10]), .out(h_s_arrmul16_and10_10));
  fa fa_h_s_arrmul16_fa10_10_out(.a(h_s_arrmul16_and10_10[0]), .b(h_s_arrmul16_fa11_9_xor1[0]), .cin(h_s_arrmul16_fa9_10_or0[0]), .fa_xor1(h_s_arrmul16_fa10_10_xor1), .fa_or0(h_s_arrmul16_fa10_10_or0));
  and_gate and_gate_h_s_arrmul16_and11_10(.a(a[11]), .b(b[10]), .out(h_s_arrmul16_and11_10));
  fa fa_h_s_arrmul16_fa11_10_out(.a(h_s_arrmul16_and11_10[0]), .b(h_s_arrmul16_fa12_9_xor1[0]), .cin(h_s_arrmul16_fa10_10_or0[0]), .fa_xor1(h_s_arrmul16_fa11_10_xor1), .fa_or0(h_s_arrmul16_fa11_10_or0));
  and_gate and_gate_h_s_arrmul16_and12_10(.a(a[12]), .b(b[10]), .out(h_s_arrmul16_and12_10));
  fa fa_h_s_arrmul16_fa12_10_out(.a(h_s_arrmul16_and12_10[0]), .b(h_s_arrmul16_fa13_9_xor1[0]), .cin(h_s_arrmul16_fa11_10_or0[0]), .fa_xor1(h_s_arrmul16_fa12_10_xor1), .fa_or0(h_s_arrmul16_fa12_10_or0));
  and_gate and_gate_h_s_arrmul16_and13_10(.a(a[13]), .b(b[10]), .out(h_s_arrmul16_and13_10));
  fa fa_h_s_arrmul16_fa13_10_out(.a(h_s_arrmul16_and13_10[0]), .b(h_s_arrmul16_fa14_9_xor1[0]), .cin(h_s_arrmul16_fa12_10_or0[0]), .fa_xor1(h_s_arrmul16_fa13_10_xor1), .fa_or0(h_s_arrmul16_fa13_10_or0));
  and_gate and_gate_h_s_arrmul16_and14_10(.a(a[14]), .b(b[10]), .out(h_s_arrmul16_and14_10));
  fa fa_h_s_arrmul16_fa14_10_out(.a(h_s_arrmul16_and14_10[0]), .b(h_s_arrmul16_fa15_9_xor1[0]), .cin(h_s_arrmul16_fa13_10_or0[0]), .fa_xor1(h_s_arrmul16_fa14_10_xor1), .fa_or0(h_s_arrmul16_fa14_10_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_10(.a(a[15]), .b(b[10]), .out(h_s_arrmul16_nand15_10));
  fa fa_h_s_arrmul16_fa15_10_out(.a(h_s_arrmul16_nand15_10[0]), .b(h_s_arrmul16_fa15_9_or0[0]), .cin(h_s_arrmul16_fa14_10_or0[0]), .fa_xor1(h_s_arrmul16_fa15_10_xor1), .fa_or0(h_s_arrmul16_fa15_10_or0));
  and_gate and_gate_h_s_arrmul16_and0_11(.a(a[0]), .b(b[11]), .out(h_s_arrmul16_and0_11));
  ha ha_h_s_arrmul16_ha0_11_out(.a(h_s_arrmul16_and0_11[0]), .b(h_s_arrmul16_fa1_10_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_11_xor0), .ha_and0(h_s_arrmul16_ha0_11_and0));
  and_gate and_gate_h_s_arrmul16_and1_11(.a(a[1]), .b(b[11]), .out(h_s_arrmul16_and1_11));
  fa fa_h_s_arrmul16_fa1_11_out(.a(h_s_arrmul16_and1_11[0]), .b(h_s_arrmul16_fa2_10_xor1[0]), .cin(h_s_arrmul16_ha0_11_and0[0]), .fa_xor1(h_s_arrmul16_fa1_11_xor1), .fa_or0(h_s_arrmul16_fa1_11_or0));
  and_gate and_gate_h_s_arrmul16_and2_11(.a(a[2]), .b(b[11]), .out(h_s_arrmul16_and2_11));
  fa fa_h_s_arrmul16_fa2_11_out(.a(h_s_arrmul16_and2_11[0]), .b(h_s_arrmul16_fa3_10_xor1[0]), .cin(h_s_arrmul16_fa1_11_or0[0]), .fa_xor1(h_s_arrmul16_fa2_11_xor1), .fa_or0(h_s_arrmul16_fa2_11_or0));
  and_gate and_gate_h_s_arrmul16_and3_11(.a(a[3]), .b(b[11]), .out(h_s_arrmul16_and3_11));
  fa fa_h_s_arrmul16_fa3_11_out(.a(h_s_arrmul16_and3_11[0]), .b(h_s_arrmul16_fa4_10_xor1[0]), .cin(h_s_arrmul16_fa2_11_or0[0]), .fa_xor1(h_s_arrmul16_fa3_11_xor1), .fa_or0(h_s_arrmul16_fa3_11_or0));
  and_gate and_gate_h_s_arrmul16_and4_11(.a(a[4]), .b(b[11]), .out(h_s_arrmul16_and4_11));
  fa fa_h_s_arrmul16_fa4_11_out(.a(h_s_arrmul16_and4_11[0]), .b(h_s_arrmul16_fa5_10_xor1[0]), .cin(h_s_arrmul16_fa3_11_or0[0]), .fa_xor1(h_s_arrmul16_fa4_11_xor1), .fa_or0(h_s_arrmul16_fa4_11_or0));
  and_gate and_gate_h_s_arrmul16_and5_11(.a(a[5]), .b(b[11]), .out(h_s_arrmul16_and5_11));
  fa fa_h_s_arrmul16_fa5_11_out(.a(h_s_arrmul16_and5_11[0]), .b(h_s_arrmul16_fa6_10_xor1[0]), .cin(h_s_arrmul16_fa4_11_or0[0]), .fa_xor1(h_s_arrmul16_fa5_11_xor1), .fa_or0(h_s_arrmul16_fa5_11_or0));
  and_gate and_gate_h_s_arrmul16_and6_11(.a(a[6]), .b(b[11]), .out(h_s_arrmul16_and6_11));
  fa fa_h_s_arrmul16_fa6_11_out(.a(h_s_arrmul16_and6_11[0]), .b(h_s_arrmul16_fa7_10_xor1[0]), .cin(h_s_arrmul16_fa5_11_or0[0]), .fa_xor1(h_s_arrmul16_fa6_11_xor1), .fa_or0(h_s_arrmul16_fa6_11_or0));
  and_gate and_gate_h_s_arrmul16_and7_11(.a(a[7]), .b(b[11]), .out(h_s_arrmul16_and7_11));
  fa fa_h_s_arrmul16_fa7_11_out(.a(h_s_arrmul16_and7_11[0]), .b(h_s_arrmul16_fa8_10_xor1[0]), .cin(h_s_arrmul16_fa6_11_or0[0]), .fa_xor1(h_s_arrmul16_fa7_11_xor1), .fa_or0(h_s_arrmul16_fa7_11_or0));
  and_gate and_gate_h_s_arrmul16_and8_11(.a(a[8]), .b(b[11]), .out(h_s_arrmul16_and8_11));
  fa fa_h_s_arrmul16_fa8_11_out(.a(h_s_arrmul16_and8_11[0]), .b(h_s_arrmul16_fa9_10_xor1[0]), .cin(h_s_arrmul16_fa7_11_or0[0]), .fa_xor1(h_s_arrmul16_fa8_11_xor1), .fa_or0(h_s_arrmul16_fa8_11_or0));
  and_gate and_gate_h_s_arrmul16_and9_11(.a(a[9]), .b(b[11]), .out(h_s_arrmul16_and9_11));
  fa fa_h_s_arrmul16_fa9_11_out(.a(h_s_arrmul16_and9_11[0]), .b(h_s_arrmul16_fa10_10_xor1[0]), .cin(h_s_arrmul16_fa8_11_or0[0]), .fa_xor1(h_s_arrmul16_fa9_11_xor1), .fa_or0(h_s_arrmul16_fa9_11_or0));
  and_gate and_gate_h_s_arrmul16_and10_11(.a(a[10]), .b(b[11]), .out(h_s_arrmul16_and10_11));
  fa fa_h_s_arrmul16_fa10_11_out(.a(h_s_arrmul16_and10_11[0]), .b(h_s_arrmul16_fa11_10_xor1[0]), .cin(h_s_arrmul16_fa9_11_or0[0]), .fa_xor1(h_s_arrmul16_fa10_11_xor1), .fa_or0(h_s_arrmul16_fa10_11_or0));
  and_gate and_gate_h_s_arrmul16_and11_11(.a(a[11]), .b(b[11]), .out(h_s_arrmul16_and11_11));
  fa fa_h_s_arrmul16_fa11_11_out(.a(h_s_arrmul16_and11_11[0]), .b(h_s_arrmul16_fa12_10_xor1[0]), .cin(h_s_arrmul16_fa10_11_or0[0]), .fa_xor1(h_s_arrmul16_fa11_11_xor1), .fa_or0(h_s_arrmul16_fa11_11_or0));
  and_gate and_gate_h_s_arrmul16_and12_11(.a(a[12]), .b(b[11]), .out(h_s_arrmul16_and12_11));
  fa fa_h_s_arrmul16_fa12_11_out(.a(h_s_arrmul16_and12_11[0]), .b(h_s_arrmul16_fa13_10_xor1[0]), .cin(h_s_arrmul16_fa11_11_or0[0]), .fa_xor1(h_s_arrmul16_fa12_11_xor1), .fa_or0(h_s_arrmul16_fa12_11_or0));
  and_gate and_gate_h_s_arrmul16_and13_11(.a(a[13]), .b(b[11]), .out(h_s_arrmul16_and13_11));
  fa fa_h_s_arrmul16_fa13_11_out(.a(h_s_arrmul16_and13_11[0]), .b(h_s_arrmul16_fa14_10_xor1[0]), .cin(h_s_arrmul16_fa12_11_or0[0]), .fa_xor1(h_s_arrmul16_fa13_11_xor1), .fa_or0(h_s_arrmul16_fa13_11_or0));
  and_gate and_gate_h_s_arrmul16_and14_11(.a(a[14]), .b(b[11]), .out(h_s_arrmul16_and14_11));
  fa fa_h_s_arrmul16_fa14_11_out(.a(h_s_arrmul16_and14_11[0]), .b(h_s_arrmul16_fa15_10_xor1[0]), .cin(h_s_arrmul16_fa13_11_or0[0]), .fa_xor1(h_s_arrmul16_fa14_11_xor1), .fa_or0(h_s_arrmul16_fa14_11_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_11(.a(a[15]), .b(b[11]), .out(h_s_arrmul16_nand15_11));
  fa fa_h_s_arrmul16_fa15_11_out(.a(h_s_arrmul16_nand15_11[0]), .b(h_s_arrmul16_fa15_10_or0[0]), .cin(h_s_arrmul16_fa14_11_or0[0]), .fa_xor1(h_s_arrmul16_fa15_11_xor1), .fa_or0(h_s_arrmul16_fa15_11_or0));
  and_gate and_gate_h_s_arrmul16_and0_12(.a(a[0]), .b(b[12]), .out(h_s_arrmul16_and0_12));
  ha ha_h_s_arrmul16_ha0_12_out(.a(h_s_arrmul16_and0_12[0]), .b(h_s_arrmul16_fa1_11_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_12_xor0), .ha_and0(h_s_arrmul16_ha0_12_and0));
  and_gate and_gate_h_s_arrmul16_and1_12(.a(a[1]), .b(b[12]), .out(h_s_arrmul16_and1_12));
  fa fa_h_s_arrmul16_fa1_12_out(.a(h_s_arrmul16_and1_12[0]), .b(h_s_arrmul16_fa2_11_xor1[0]), .cin(h_s_arrmul16_ha0_12_and0[0]), .fa_xor1(h_s_arrmul16_fa1_12_xor1), .fa_or0(h_s_arrmul16_fa1_12_or0));
  and_gate and_gate_h_s_arrmul16_and2_12(.a(a[2]), .b(b[12]), .out(h_s_arrmul16_and2_12));
  fa fa_h_s_arrmul16_fa2_12_out(.a(h_s_arrmul16_and2_12[0]), .b(h_s_arrmul16_fa3_11_xor1[0]), .cin(h_s_arrmul16_fa1_12_or0[0]), .fa_xor1(h_s_arrmul16_fa2_12_xor1), .fa_or0(h_s_arrmul16_fa2_12_or0));
  and_gate and_gate_h_s_arrmul16_and3_12(.a(a[3]), .b(b[12]), .out(h_s_arrmul16_and3_12));
  fa fa_h_s_arrmul16_fa3_12_out(.a(h_s_arrmul16_and3_12[0]), .b(h_s_arrmul16_fa4_11_xor1[0]), .cin(h_s_arrmul16_fa2_12_or0[0]), .fa_xor1(h_s_arrmul16_fa3_12_xor1), .fa_or0(h_s_arrmul16_fa3_12_or0));
  and_gate and_gate_h_s_arrmul16_and4_12(.a(a[4]), .b(b[12]), .out(h_s_arrmul16_and4_12));
  fa fa_h_s_arrmul16_fa4_12_out(.a(h_s_arrmul16_and4_12[0]), .b(h_s_arrmul16_fa5_11_xor1[0]), .cin(h_s_arrmul16_fa3_12_or0[0]), .fa_xor1(h_s_arrmul16_fa4_12_xor1), .fa_or0(h_s_arrmul16_fa4_12_or0));
  and_gate and_gate_h_s_arrmul16_and5_12(.a(a[5]), .b(b[12]), .out(h_s_arrmul16_and5_12));
  fa fa_h_s_arrmul16_fa5_12_out(.a(h_s_arrmul16_and5_12[0]), .b(h_s_arrmul16_fa6_11_xor1[0]), .cin(h_s_arrmul16_fa4_12_or0[0]), .fa_xor1(h_s_arrmul16_fa5_12_xor1), .fa_or0(h_s_arrmul16_fa5_12_or0));
  and_gate and_gate_h_s_arrmul16_and6_12(.a(a[6]), .b(b[12]), .out(h_s_arrmul16_and6_12));
  fa fa_h_s_arrmul16_fa6_12_out(.a(h_s_arrmul16_and6_12[0]), .b(h_s_arrmul16_fa7_11_xor1[0]), .cin(h_s_arrmul16_fa5_12_or0[0]), .fa_xor1(h_s_arrmul16_fa6_12_xor1), .fa_or0(h_s_arrmul16_fa6_12_or0));
  and_gate and_gate_h_s_arrmul16_and7_12(.a(a[7]), .b(b[12]), .out(h_s_arrmul16_and7_12));
  fa fa_h_s_arrmul16_fa7_12_out(.a(h_s_arrmul16_and7_12[0]), .b(h_s_arrmul16_fa8_11_xor1[0]), .cin(h_s_arrmul16_fa6_12_or0[0]), .fa_xor1(h_s_arrmul16_fa7_12_xor1), .fa_or0(h_s_arrmul16_fa7_12_or0));
  and_gate and_gate_h_s_arrmul16_and8_12(.a(a[8]), .b(b[12]), .out(h_s_arrmul16_and8_12));
  fa fa_h_s_arrmul16_fa8_12_out(.a(h_s_arrmul16_and8_12[0]), .b(h_s_arrmul16_fa9_11_xor1[0]), .cin(h_s_arrmul16_fa7_12_or0[0]), .fa_xor1(h_s_arrmul16_fa8_12_xor1), .fa_or0(h_s_arrmul16_fa8_12_or0));
  and_gate and_gate_h_s_arrmul16_and9_12(.a(a[9]), .b(b[12]), .out(h_s_arrmul16_and9_12));
  fa fa_h_s_arrmul16_fa9_12_out(.a(h_s_arrmul16_and9_12[0]), .b(h_s_arrmul16_fa10_11_xor1[0]), .cin(h_s_arrmul16_fa8_12_or0[0]), .fa_xor1(h_s_arrmul16_fa9_12_xor1), .fa_or0(h_s_arrmul16_fa9_12_or0));
  and_gate and_gate_h_s_arrmul16_and10_12(.a(a[10]), .b(b[12]), .out(h_s_arrmul16_and10_12));
  fa fa_h_s_arrmul16_fa10_12_out(.a(h_s_arrmul16_and10_12[0]), .b(h_s_arrmul16_fa11_11_xor1[0]), .cin(h_s_arrmul16_fa9_12_or0[0]), .fa_xor1(h_s_arrmul16_fa10_12_xor1), .fa_or0(h_s_arrmul16_fa10_12_or0));
  and_gate and_gate_h_s_arrmul16_and11_12(.a(a[11]), .b(b[12]), .out(h_s_arrmul16_and11_12));
  fa fa_h_s_arrmul16_fa11_12_out(.a(h_s_arrmul16_and11_12[0]), .b(h_s_arrmul16_fa12_11_xor1[0]), .cin(h_s_arrmul16_fa10_12_or0[0]), .fa_xor1(h_s_arrmul16_fa11_12_xor1), .fa_or0(h_s_arrmul16_fa11_12_or0));
  and_gate and_gate_h_s_arrmul16_and12_12(.a(a[12]), .b(b[12]), .out(h_s_arrmul16_and12_12));
  fa fa_h_s_arrmul16_fa12_12_out(.a(h_s_arrmul16_and12_12[0]), .b(h_s_arrmul16_fa13_11_xor1[0]), .cin(h_s_arrmul16_fa11_12_or0[0]), .fa_xor1(h_s_arrmul16_fa12_12_xor1), .fa_or0(h_s_arrmul16_fa12_12_or0));
  and_gate and_gate_h_s_arrmul16_and13_12(.a(a[13]), .b(b[12]), .out(h_s_arrmul16_and13_12));
  fa fa_h_s_arrmul16_fa13_12_out(.a(h_s_arrmul16_and13_12[0]), .b(h_s_arrmul16_fa14_11_xor1[0]), .cin(h_s_arrmul16_fa12_12_or0[0]), .fa_xor1(h_s_arrmul16_fa13_12_xor1), .fa_or0(h_s_arrmul16_fa13_12_or0));
  and_gate and_gate_h_s_arrmul16_and14_12(.a(a[14]), .b(b[12]), .out(h_s_arrmul16_and14_12));
  fa fa_h_s_arrmul16_fa14_12_out(.a(h_s_arrmul16_and14_12[0]), .b(h_s_arrmul16_fa15_11_xor1[0]), .cin(h_s_arrmul16_fa13_12_or0[0]), .fa_xor1(h_s_arrmul16_fa14_12_xor1), .fa_or0(h_s_arrmul16_fa14_12_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_12(.a(a[15]), .b(b[12]), .out(h_s_arrmul16_nand15_12));
  fa fa_h_s_arrmul16_fa15_12_out(.a(h_s_arrmul16_nand15_12[0]), .b(h_s_arrmul16_fa15_11_or0[0]), .cin(h_s_arrmul16_fa14_12_or0[0]), .fa_xor1(h_s_arrmul16_fa15_12_xor1), .fa_or0(h_s_arrmul16_fa15_12_or0));
  and_gate and_gate_h_s_arrmul16_and0_13(.a(a[0]), .b(b[13]), .out(h_s_arrmul16_and0_13));
  ha ha_h_s_arrmul16_ha0_13_out(.a(h_s_arrmul16_and0_13[0]), .b(h_s_arrmul16_fa1_12_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_13_xor0), .ha_and0(h_s_arrmul16_ha0_13_and0));
  and_gate and_gate_h_s_arrmul16_and1_13(.a(a[1]), .b(b[13]), .out(h_s_arrmul16_and1_13));
  fa fa_h_s_arrmul16_fa1_13_out(.a(h_s_arrmul16_and1_13[0]), .b(h_s_arrmul16_fa2_12_xor1[0]), .cin(h_s_arrmul16_ha0_13_and0[0]), .fa_xor1(h_s_arrmul16_fa1_13_xor1), .fa_or0(h_s_arrmul16_fa1_13_or0));
  and_gate and_gate_h_s_arrmul16_and2_13(.a(a[2]), .b(b[13]), .out(h_s_arrmul16_and2_13));
  fa fa_h_s_arrmul16_fa2_13_out(.a(h_s_arrmul16_and2_13[0]), .b(h_s_arrmul16_fa3_12_xor1[0]), .cin(h_s_arrmul16_fa1_13_or0[0]), .fa_xor1(h_s_arrmul16_fa2_13_xor1), .fa_or0(h_s_arrmul16_fa2_13_or0));
  and_gate and_gate_h_s_arrmul16_and3_13(.a(a[3]), .b(b[13]), .out(h_s_arrmul16_and3_13));
  fa fa_h_s_arrmul16_fa3_13_out(.a(h_s_arrmul16_and3_13[0]), .b(h_s_arrmul16_fa4_12_xor1[0]), .cin(h_s_arrmul16_fa2_13_or0[0]), .fa_xor1(h_s_arrmul16_fa3_13_xor1), .fa_or0(h_s_arrmul16_fa3_13_or0));
  and_gate and_gate_h_s_arrmul16_and4_13(.a(a[4]), .b(b[13]), .out(h_s_arrmul16_and4_13));
  fa fa_h_s_arrmul16_fa4_13_out(.a(h_s_arrmul16_and4_13[0]), .b(h_s_arrmul16_fa5_12_xor1[0]), .cin(h_s_arrmul16_fa3_13_or0[0]), .fa_xor1(h_s_arrmul16_fa4_13_xor1), .fa_or0(h_s_arrmul16_fa4_13_or0));
  and_gate and_gate_h_s_arrmul16_and5_13(.a(a[5]), .b(b[13]), .out(h_s_arrmul16_and5_13));
  fa fa_h_s_arrmul16_fa5_13_out(.a(h_s_arrmul16_and5_13[0]), .b(h_s_arrmul16_fa6_12_xor1[0]), .cin(h_s_arrmul16_fa4_13_or0[0]), .fa_xor1(h_s_arrmul16_fa5_13_xor1), .fa_or0(h_s_arrmul16_fa5_13_or0));
  and_gate and_gate_h_s_arrmul16_and6_13(.a(a[6]), .b(b[13]), .out(h_s_arrmul16_and6_13));
  fa fa_h_s_arrmul16_fa6_13_out(.a(h_s_arrmul16_and6_13[0]), .b(h_s_arrmul16_fa7_12_xor1[0]), .cin(h_s_arrmul16_fa5_13_or0[0]), .fa_xor1(h_s_arrmul16_fa6_13_xor1), .fa_or0(h_s_arrmul16_fa6_13_or0));
  and_gate and_gate_h_s_arrmul16_and7_13(.a(a[7]), .b(b[13]), .out(h_s_arrmul16_and7_13));
  fa fa_h_s_arrmul16_fa7_13_out(.a(h_s_arrmul16_and7_13[0]), .b(h_s_arrmul16_fa8_12_xor1[0]), .cin(h_s_arrmul16_fa6_13_or0[0]), .fa_xor1(h_s_arrmul16_fa7_13_xor1), .fa_or0(h_s_arrmul16_fa7_13_or0));
  and_gate and_gate_h_s_arrmul16_and8_13(.a(a[8]), .b(b[13]), .out(h_s_arrmul16_and8_13));
  fa fa_h_s_arrmul16_fa8_13_out(.a(h_s_arrmul16_and8_13[0]), .b(h_s_arrmul16_fa9_12_xor1[0]), .cin(h_s_arrmul16_fa7_13_or0[0]), .fa_xor1(h_s_arrmul16_fa8_13_xor1), .fa_or0(h_s_arrmul16_fa8_13_or0));
  and_gate and_gate_h_s_arrmul16_and9_13(.a(a[9]), .b(b[13]), .out(h_s_arrmul16_and9_13));
  fa fa_h_s_arrmul16_fa9_13_out(.a(h_s_arrmul16_and9_13[0]), .b(h_s_arrmul16_fa10_12_xor1[0]), .cin(h_s_arrmul16_fa8_13_or0[0]), .fa_xor1(h_s_arrmul16_fa9_13_xor1), .fa_or0(h_s_arrmul16_fa9_13_or0));
  and_gate and_gate_h_s_arrmul16_and10_13(.a(a[10]), .b(b[13]), .out(h_s_arrmul16_and10_13));
  fa fa_h_s_arrmul16_fa10_13_out(.a(h_s_arrmul16_and10_13[0]), .b(h_s_arrmul16_fa11_12_xor1[0]), .cin(h_s_arrmul16_fa9_13_or0[0]), .fa_xor1(h_s_arrmul16_fa10_13_xor1), .fa_or0(h_s_arrmul16_fa10_13_or0));
  and_gate and_gate_h_s_arrmul16_and11_13(.a(a[11]), .b(b[13]), .out(h_s_arrmul16_and11_13));
  fa fa_h_s_arrmul16_fa11_13_out(.a(h_s_arrmul16_and11_13[0]), .b(h_s_arrmul16_fa12_12_xor1[0]), .cin(h_s_arrmul16_fa10_13_or0[0]), .fa_xor1(h_s_arrmul16_fa11_13_xor1), .fa_or0(h_s_arrmul16_fa11_13_or0));
  and_gate and_gate_h_s_arrmul16_and12_13(.a(a[12]), .b(b[13]), .out(h_s_arrmul16_and12_13));
  fa fa_h_s_arrmul16_fa12_13_out(.a(h_s_arrmul16_and12_13[0]), .b(h_s_arrmul16_fa13_12_xor1[0]), .cin(h_s_arrmul16_fa11_13_or0[0]), .fa_xor1(h_s_arrmul16_fa12_13_xor1), .fa_or0(h_s_arrmul16_fa12_13_or0));
  and_gate and_gate_h_s_arrmul16_and13_13(.a(a[13]), .b(b[13]), .out(h_s_arrmul16_and13_13));
  fa fa_h_s_arrmul16_fa13_13_out(.a(h_s_arrmul16_and13_13[0]), .b(h_s_arrmul16_fa14_12_xor1[0]), .cin(h_s_arrmul16_fa12_13_or0[0]), .fa_xor1(h_s_arrmul16_fa13_13_xor1), .fa_or0(h_s_arrmul16_fa13_13_or0));
  and_gate and_gate_h_s_arrmul16_and14_13(.a(a[14]), .b(b[13]), .out(h_s_arrmul16_and14_13));
  fa fa_h_s_arrmul16_fa14_13_out(.a(h_s_arrmul16_and14_13[0]), .b(h_s_arrmul16_fa15_12_xor1[0]), .cin(h_s_arrmul16_fa13_13_or0[0]), .fa_xor1(h_s_arrmul16_fa14_13_xor1), .fa_or0(h_s_arrmul16_fa14_13_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_13(.a(a[15]), .b(b[13]), .out(h_s_arrmul16_nand15_13));
  fa fa_h_s_arrmul16_fa15_13_out(.a(h_s_arrmul16_nand15_13[0]), .b(h_s_arrmul16_fa15_12_or0[0]), .cin(h_s_arrmul16_fa14_13_or0[0]), .fa_xor1(h_s_arrmul16_fa15_13_xor1), .fa_or0(h_s_arrmul16_fa15_13_or0));
  and_gate and_gate_h_s_arrmul16_and0_14(.a(a[0]), .b(b[14]), .out(h_s_arrmul16_and0_14));
  ha ha_h_s_arrmul16_ha0_14_out(.a(h_s_arrmul16_and0_14[0]), .b(h_s_arrmul16_fa1_13_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_14_xor0), .ha_and0(h_s_arrmul16_ha0_14_and0));
  and_gate and_gate_h_s_arrmul16_and1_14(.a(a[1]), .b(b[14]), .out(h_s_arrmul16_and1_14));
  fa fa_h_s_arrmul16_fa1_14_out(.a(h_s_arrmul16_and1_14[0]), .b(h_s_arrmul16_fa2_13_xor1[0]), .cin(h_s_arrmul16_ha0_14_and0[0]), .fa_xor1(h_s_arrmul16_fa1_14_xor1), .fa_or0(h_s_arrmul16_fa1_14_or0));
  and_gate and_gate_h_s_arrmul16_and2_14(.a(a[2]), .b(b[14]), .out(h_s_arrmul16_and2_14));
  fa fa_h_s_arrmul16_fa2_14_out(.a(h_s_arrmul16_and2_14[0]), .b(h_s_arrmul16_fa3_13_xor1[0]), .cin(h_s_arrmul16_fa1_14_or0[0]), .fa_xor1(h_s_arrmul16_fa2_14_xor1), .fa_or0(h_s_arrmul16_fa2_14_or0));
  and_gate and_gate_h_s_arrmul16_and3_14(.a(a[3]), .b(b[14]), .out(h_s_arrmul16_and3_14));
  fa fa_h_s_arrmul16_fa3_14_out(.a(h_s_arrmul16_and3_14[0]), .b(h_s_arrmul16_fa4_13_xor1[0]), .cin(h_s_arrmul16_fa2_14_or0[0]), .fa_xor1(h_s_arrmul16_fa3_14_xor1), .fa_or0(h_s_arrmul16_fa3_14_or0));
  and_gate and_gate_h_s_arrmul16_and4_14(.a(a[4]), .b(b[14]), .out(h_s_arrmul16_and4_14));
  fa fa_h_s_arrmul16_fa4_14_out(.a(h_s_arrmul16_and4_14[0]), .b(h_s_arrmul16_fa5_13_xor1[0]), .cin(h_s_arrmul16_fa3_14_or0[0]), .fa_xor1(h_s_arrmul16_fa4_14_xor1), .fa_or0(h_s_arrmul16_fa4_14_or0));
  and_gate and_gate_h_s_arrmul16_and5_14(.a(a[5]), .b(b[14]), .out(h_s_arrmul16_and5_14));
  fa fa_h_s_arrmul16_fa5_14_out(.a(h_s_arrmul16_and5_14[0]), .b(h_s_arrmul16_fa6_13_xor1[0]), .cin(h_s_arrmul16_fa4_14_or0[0]), .fa_xor1(h_s_arrmul16_fa5_14_xor1), .fa_or0(h_s_arrmul16_fa5_14_or0));
  and_gate and_gate_h_s_arrmul16_and6_14(.a(a[6]), .b(b[14]), .out(h_s_arrmul16_and6_14));
  fa fa_h_s_arrmul16_fa6_14_out(.a(h_s_arrmul16_and6_14[0]), .b(h_s_arrmul16_fa7_13_xor1[0]), .cin(h_s_arrmul16_fa5_14_or0[0]), .fa_xor1(h_s_arrmul16_fa6_14_xor1), .fa_or0(h_s_arrmul16_fa6_14_or0));
  and_gate and_gate_h_s_arrmul16_and7_14(.a(a[7]), .b(b[14]), .out(h_s_arrmul16_and7_14));
  fa fa_h_s_arrmul16_fa7_14_out(.a(h_s_arrmul16_and7_14[0]), .b(h_s_arrmul16_fa8_13_xor1[0]), .cin(h_s_arrmul16_fa6_14_or0[0]), .fa_xor1(h_s_arrmul16_fa7_14_xor1), .fa_or0(h_s_arrmul16_fa7_14_or0));
  and_gate and_gate_h_s_arrmul16_and8_14(.a(a[8]), .b(b[14]), .out(h_s_arrmul16_and8_14));
  fa fa_h_s_arrmul16_fa8_14_out(.a(h_s_arrmul16_and8_14[0]), .b(h_s_arrmul16_fa9_13_xor1[0]), .cin(h_s_arrmul16_fa7_14_or0[0]), .fa_xor1(h_s_arrmul16_fa8_14_xor1), .fa_or0(h_s_arrmul16_fa8_14_or0));
  and_gate and_gate_h_s_arrmul16_and9_14(.a(a[9]), .b(b[14]), .out(h_s_arrmul16_and9_14));
  fa fa_h_s_arrmul16_fa9_14_out(.a(h_s_arrmul16_and9_14[0]), .b(h_s_arrmul16_fa10_13_xor1[0]), .cin(h_s_arrmul16_fa8_14_or0[0]), .fa_xor1(h_s_arrmul16_fa9_14_xor1), .fa_or0(h_s_arrmul16_fa9_14_or0));
  and_gate and_gate_h_s_arrmul16_and10_14(.a(a[10]), .b(b[14]), .out(h_s_arrmul16_and10_14));
  fa fa_h_s_arrmul16_fa10_14_out(.a(h_s_arrmul16_and10_14[0]), .b(h_s_arrmul16_fa11_13_xor1[0]), .cin(h_s_arrmul16_fa9_14_or0[0]), .fa_xor1(h_s_arrmul16_fa10_14_xor1), .fa_or0(h_s_arrmul16_fa10_14_or0));
  and_gate and_gate_h_s_arrmul16_and11_14(.a(a[11]), .b(b[14]), .out(h_s_arrmul16_and11_14));
  fa fa_h_s_arrmul16_fa11_14_out(.a(h_s_arrmul16_and11_14[0]), .b(h_s_arrmul16_fa12_13_xor1[0]), .cin(h_s_arrmul16_fa10_14_or0[0]), .fa_xor1(h_s_arrmul16_fa11_14_xor1), .fa_or0(h_s_arrmul16_fa11_14_or0));
  and_gate and_gate_h_s_arrmul16_and12_14(.a(a[12]), .b(b[14]), .out(h_s_arrmul16_and12_14));
  fa fa_h_s_arrmul16_fa12_14_out(.a(h_s_arrmul16_and12_14[0]), .b(h_s_arrmul16_fa13_13_xor1[0]), .cin(h_s_arrmul16_fa11_14_or0[0]), .fa_xor1(h_s_arrmul16_fa12_14_xor1), .fa_or0(h_s_arrmul16_fa12_14_or0));
  and_gate and_gate_h_s_arrmul16_and13_14(.a(a[13]), .b(b[14]), .out(h_s_arrmul16_and13_14));
  fa fa_h_s_arrmul16_fa13_14_out(.a(h_s_arrmul16_and13_14[0]), .b(h_s_arrmul16_fa14_13_xor1[0]), .cin(h_s_arrmul16_fa12_14_or0[0]), .fa_xor1(h_s_arrmul16_fa13_14_xor1), .fa_or0(h_s_arrmul16_fa13_14_or0));
  and_gate and_gate_h_s_arrmul16_and14_14(.a(a[14]), .b(b[14]), .out(h_s_arrmul16_and14_14));
  fa fa_h_s_arrmul16_fa14_14_out(.a(h_s_arrmul16_and14_14[0]), .b(h_s_arrmul16_fa15_13_xor1[0]), .cin(h_s_arrmul16_fa13_14_or0[0]), .fa_xor1(h_s_arrmul16_fa14_14_xor1), .fa_or0(h_s_arrmul16_fa14_14_or0));
  nand_gate nand_gate_h_s_arrmul16_nand15_14(.a(a[15]), .b(b[14]), .out(h_s_arrmul16_nand15_14));
  fa fa_h_s_arrmul16_fa15_14_out(.a(h_s_arrmul16_nand15_14[0]), .b(h_s_arrmul16_fa15_13_or0[0]), .cin(h_s_arrmul16_fa14_14_or0[0]), .fa_xor1(h_s_arrmul16_fa15_14_xor1), .fa_or0(h_s_arrmul16_fa15_14_or0));
  nand_gate nand_gate_h_s_arrmul16_nand0_15(.a(a[0]), .b(b[15]), .out(h_s_arrmul16_nand0_15));
  ha ha_h_s_arrmul16_ha0_15_out(.a(h_s_arrmul16_nand0_15[0]), .b(h_s_arrmul16_fa1_14_xor1[0]), .ha_xor0(h_s_arrmul16_ha0_15_xor0), .ha_and0(h_s_arrmul16_ha0_15_and0));
  nand_gate nand_gate_h_s_arrmul16_nand1_15(.a(a[1]), .b(b[15]), .out(h_s_arrmul16_nand1_15));
  fa fa_h_s_arrmul16_fa1_15_out(.a(h_s_arrmul16_nand1_15[0]), .b(h_s_arrmul16_fa2_14_xor1[0]), .cin(h_s_arrmul16_ha0_15_and0[0]), .fa_xor1(h_s_arrmul16_fa1_15_xor1), .fa_or0(h_s_arrmul16_fa1_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand2_15(.a(a[2]), .b(b[15]), .out(h_s_arrmul16_nand2_15));
  fa fa_h_s_arrmul16_fa2_15_out(.a(h_s_arrmul16_nand2_15[0]), .b(h_s_arrmul16_fa3_14_xor1[0]), .cin(h_s_arrmul16_fa1_15_or0[0]), .fa_xor1(h_s_arrmul16_fa2_15_xor1), .fa_or0(h_s_arrmul16_fa2_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand3_15(.a(a[3]), .b(b[15]), .out(h_s_arrmul16_nand3_15));
  fa fa_h_s_arrmul16_fa3_15_out(.a(h_s_arrmul16_nand3_15[0]), .b(h_s_arrmul16_fa4_14_xor1[0]), .cin(h_s_arrmul16_fa2_15_or0[0]), .fa_xor1(h_s_arrmul16_fa3_15_xor1), .fa_or0(h_s_arrmul16_fa3_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand4_15(.a(a[4]), .b(b[15]), .out(h_s_arrmul16_nand4_15));
  fa fa_h_s_arrmul16_fa4_15_out(.a(h_s_arrmul16_nand4_15[0]), .b(h_s_arrmul16_fa5_14_xor1[0]), .cin(h_s_arrmul16_fa3_15_or0[0]), .fa_xor1(h_s_arrmul16_fa4_15_xor1), .fa_or0(h_s_arrmul16_fa4_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand5_15(.a(a[5]), .b(b[15]), .out(h_s_arrmul16_nand5_15));
  fa fa_h_s_arrmul16_fa5_15_out(.a(h_s_arrmul16_nand5_15[0]), .b(h_s_arrmul16_fa6_14_xor1[0]), .cin(h_s_arrmul16_fa4_15_or0[0]), .fa_xor1(h_s_arrmul16_fa5_15_xor1), .fa_or0(h_s_arrmul16_fa5_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand6_15(.a(a[6]), .b(b[15]), .out(h_s_arrmul16_nand6_15));
  fa fa_h_s_arrmul16_fa6_15_out(.a(h_s_arrmul16_nand6_15[0]), .b(h_s_arrmul16_fa7_14_xor1[0]), .cin(h_s_arrmul16_fa5_15_or0[0]), .fa_xor1(h_s_arrmul16_fa6_15_xor1), .fa_or0(h_s_arrmul16_fa6_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand7_15(.a(a[7]), .b(b[15]), .out(h_s_arrmul16_nand7_15));
  fa fa_h_s_arrmul16_fa7_15_out(.a(h_s_arrmul16_nand7_15[0]), .b(h_s_arrmul16_fa8_14_xor1[0]), .cin(h_s_arrmul16_fa6_15_or0[0]), .fa_xor1(h_s_arrmul16_fa7_15_xor1), .fa_or0(h_s_arrmul16_fa7_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand8_15(.a(a[8]), .b(b[15]), .out(h_s_arrmul16_nand8_15));
  fa fa_h_s_arrmul16_fa8_15_out(.a(h_s_arrmul16_nand8_15[0]), .b(h_s_arrmul16_fa9_14_xor1[0]), .cin(h_s_arrmul16_fa7_15_or0[0]), .fa_xor1(h_s_arrmul16_fa8_15_xor1), .fa_or0(h_s_arrmul16_fa8_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand9_15(.a(a[9]), .b(b[15]), .out(h_s_arrmul16_nand9_15));
  fa fa_h_s_arrmul16_fa9_15_out(.a(h_s_arrmul16_nand9_15[0]), .b(h_s_arrmul16_fa10_14_xor1[0]), .cin(h_s_arrmul16_fa8_15_or0[0]), .fa_xor1(h_s_arrmul16_fa9_15_xor1), .fa_or0(h_s_arrmul16_fa9_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand10_15(.a(a[10]), .b(b[15]), .out(h_s_arrmul16_nand10_15));
  fa fa_h_s_arrmul16_fa10_15_out(.a(h_s_arrmul16_nand10_15[0]), .b(h_s_arrmul16_fa11_14_xor1[0]), .cin(h_s_arrmul16_fa9_15_or0[0]), .fa_xor1(h_s_arrmul16_fa10_15_xor1), .fa_or0(h_s_arrmul16_fa10_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand11_15(.a(a[11]), .b(b[15]), .out(h_s_arrmul16_nand11_15));
  fa fa_h_s_arrmul16_fa11_15_out(.a(h_s_arrmul16_nand11_15[0]), .b(h_s_arrmul16_fa12_14_xor1[0]), .cin(h_s_arrmul16_fa10_15_or0[0]), .fa_xor1(h_s_arrmul16_fa11_15_xor1), .fa_or0(h_s_arrmul16_fa11_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand12_15(.a(a[12]), .b(b[15]), .out(h_s_arrmul16_nand12_15));
  fa fa_h_s_arrmul16_fa12_15_out(.a(h_s_arrmul16_nand12_15[0]), .b(h_s_arrmul16_fa13_14_xor1[0]), .cin(h_s_arrmul16_fa11_15_or0[0]), .fa_xor1(h_s_arrmul16_fa12_15_xor1), .fa_or0(h_s_arrmul16_fa12_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand13_15(.a(a[13]), .b(b[15]), .out(h_s_arrmul16_nand13_15));
  fa fa_h_s_arrmul16_fa13_15_out(.a(h_s_arrmul16_nand13_15[0]), .b(h_s_arrmul16_fa14_14_xor1[0]), .cin(h_s_arrmul16_fa12_15_or0[0]), .fa_xor1(h_s_arrmul16_fa13_15_xor1), .fa_or0(h_s_arrmul16_fa13_15_or0));
  nand_gate nand_gate_h_s_arrmul16_nand14_15(.a(a[14]), .b(b[15]), .out(h_s_arrmul16_nand14_15));
  fa fa_h_s_arrmul16_fa14_15_out(.a(h_s_arrmul16_nand14_15[0]), .b(h_s_arrmul16_fa15_14_xor1[0]), .cin(h_s_arrmul16_fa13_15_or0[0]), .fa_xor1(h_s_arrmul16_fa14_15_xor1), .fa_or0(h_s_arrmul16_fa14_15_or0));
  and_gate and_gate_h_s_arrmul16_and15_15(.a(a[15]), .b(b[15]), .out(h_s_arrmul16_and15_15));
  fa fa_h_s_arrmul16_fa15_15_out(.a(h_s_arrmul16_and15_15[0]), .b(h_s_arrmul16_fa15_14_or0[0]), .cin(h_s_arrmul16_fa14_15_or0[0]), .fa_xor1(h_s_arrmul16_fa15_15_xor1), .fa_or0(h_s_arrmul16_fa15_15_or0));
  not_gate not_gate_h_s_arrmul16_xor16_15(.a(h_s_arrmul16_fa15_15_or0[0]), .out(h_s_arrmul16_xor16_15));

  assign h_s_arrmul16_out[0] = h_s_arrmul16_and0_0[0];
  assign h_s_arrmul16_out[1] = h_s_arrmul16_ha0_1_xor0[0];
  assign h_s_arrmul16_out[2] = h_s_arrmul16_ha0_2_xor0[0];
  assign h_s_arrmul16_out[3] = h_s_arrmul16_ha0_3_xor0[0];
  assign h_s_arrmul16_out[4] = h_s_arrmul16_ha0_4_xor0[0];
  assign h_s_arrmul16_out[5] = h_s_arrmul16_ha0_5_xor0[0];
  assign h_s_arrmul16_out[6] = h_s_arrmul16_ha0_6_xor0[0];
  assign h_s_arrmul16_out[7] = h_s_arrmul16_ha0_7_xor0[0];
  assign h_s_arrmul16_out[8] = h_s_arrmul16_ha0_8_xor0[0];
  assign h_s_arrmul16_out[9] = h_s_arrmul16_ha0_9_xor0[0];
  assign h_s_arrmul16_out[10] = h_s_arrmul16_ha0_10_xor0[0];
  assign h_s_arrmul16_out[11] = h_s_arrmul16_ha0_11_xor0[0];
  assign h_s_arrmul16_out[12] = h_s_arrmul16_ha0_12_xor0[0];
  assign h_s_arrmul16_out[13] = h_s_arrmul16_ha0_13_xor0[0];
  assign h_s_arrmul16_out[14] = h_s_arrmul16_ha0_14_xor0[0];
  assign h_s_arrmul16_out[15] = h_s_arrmul16_ha0_15_xor0[0];
  assign h_s_arrmul16_out[16] = h_s_arrmul16_fa1_15_xor1[0];
  assign h_s_arrmul16_out[17] = h_s_arrmul16_fa2_15_xor1[0];
  assign h_s_arrmul16_out[18] = h_s_arrmul16_fa3_15_xor1[0];
  assign h_s_arrmul16_out[19] = h_s_arrmul16_fa4_15_xor1[0];
  assign h_s_arrmul16_out[20] = h_s_arrmul16_fa5_15_xor1[0];
  assign h_s_arrmul16_out[21] = h_s_arrmul16_fa6_15_xor1[0];
  assign h_s_arrmul16_out[22] = h_s_arrmul16_fa7_15_xor1[0];
  assign h_s_arrmul16_out[23] = h_s_arrmul16_fa8_15_xor1[0];
  assign h_s_arrmul16_out[24] = h_s_arrmul16_fa9_15_xor1[0];
  assign h_s_arrmul16_out[25] = h_s_arrmul16_fa10_15_xor1[0];
  assign h_s_arrmul16_out[26] = h_s_arrmul16_fa11_15_xor1[0];
  assign h_s_arrmul16_out[27] = h_s_arrmul16_fa12_15_xor1[0];
  assign h_s_arrmul16_out[28] = h_s_arrmul16_fa13_15_xor1[0];
  assign h_s_arrmul16_out[29] = h_s_arrmul16_fa14_15_xor1[0];
  assign h_s_arrmul16_out[30] = h_s_arrmul16_fa15_15_xor1[0];
  assign h_s_arrmul16_out[31] = h_s_arrmul16_xor16_15[0];
endmodule