module u_cla32(input [31:0] a, input [31:0] b, output [32:0] u_cla32_out);
  wire u_cla32_pg_logic0_or0;
  wire u_cla32_pg_logic0_and0;
  wire u_cla32_pg_logic0_xor0;
  wire u_cla32_pg_logic1_or0;
  wire u_cla32_pg_logic1_and0;
  wire u_cla32_pg_logic1_xor0;
  wire u_cla32_xor1;
  wire u_cla32_and0;
  wire u_cla32_or0;
  wire u_cla32_pg_logic2_or0;
  wire u_cla32_pg_logic2_and0;
  wire u_cla32_pg_logic2_xor0;
  wire u_cla32_xor2;
  wire u_cla32_and1;
  wire u_cla32_and2;
  wire u_cla32_and3;
  wire u_cla32_and4;
  wire u_cla32_or1;
  wire u_cla32_or2;
  wire u_cla32_pg_logic3_or0;
  wire u_cla32_pg_logic3_and0;
  wire u_cla32_pg_logic3_xor0;
  wire u_cla32_xor3;
  wire u_cla32_and5;
  wire u_cla32_and6;
  wire u_cla32_and7;
  wire u_cla32_and8;
  wire u_cla32_and9;
  wire u_cla32_and10;
  wire u_cla32_and11;
  wire u_cla32_or3;
  wire u_cla32_or4;
  wire u_cla32_or5;
  wire u_cla32_pg_logic4_or0;
  wire u_cla32_pg_logic4_and0;
  wire u_cla32_pg_logic4_xor0;
  wire u_cla32_xor4;
  wire u_cla32_and12;
  wire u_cla32_or6;
  wire u_cla32_pg_logic5_or0;
  wire u_cla32_pg_logic5_and0;
  wire u_cla32_pg_logic5_xor0;
  wire u_cla32_xor5;
  wire u_cla32_and13;
  wire u_cla32_and14;
  wire u_cla32_and15;
  wire u_cla32_or7;
  wire u_cla32_or8;
  wire u_cla32_pg_logic6_or0;
  wire u_cla32_pg_logic6_and0;
  wire u_cla32_pg_logic6_xor0;
  wire u_cla32_xor6;
  wire u_cla32_and16;
  wire u_cla32_and17;
  wire u_cla32_and18;
  wire u_cla32_and19;
  wire u_cla32_and20;
  wire u_cla32_and21;
  wire u_cla32_or9;
  wire u_cla32_or10;
  wire u_cla32_or11;
  wire u_cla32_pg_logic7_or0;
  wire u_cla32_pg_logic7_and0;
  wire u_cla32_pg_logic7_xor0;
  wire u_cla32_xor7;
  wire u_cla32_and22;
  wire u_cla32_and23;
  wire u_cla32_and24;
  wire u_cla32_and25;
  wire u_cla32_and26;
  wire u_cla32_and27;
  wire u_cla32_and28;
  wire u_cla32_and29;
  wire u_cla32_and30;
  wire u_cla32_and31;
  wire u_cla32_or12;
  wire u_cla32_or13;
  wire u_cla32_or14;
  wire u_cla32_or15;
  wire u_cla32_pg_logic8_or0;
  wire u_cla32_pg_logic8_and0;
  wire u_cla32_pg_logic8_xor0;
  wire u_cla32_xor8;
  wire u_cla32_and32;
  wire u_cla32_or16;
  wire u_cla32_pg_logic9_or0;
  wire u_cla32_pg_logic9_and0;
  wire u_cla32_pg_logic9_xor0;
  wire u_cla32_xor9;
  wire u_cla32_and33;
  wire u_cla32_and34;
  wire u_cla32_and35;
  wire u_cla32_or17;
  wire u_cla32_or18;
  wire u_cla32_pg_logic10_or0;
  wire u_cla32_pg_logic10_and0;
  wire u_cla32_pg_logic10_xor0;
  wire u_cla32_xor10;
  wire u_cla32_and36;
  wire u_cla32_and37;
  wire u_cla32_and38;
  wire u_cla32_and39;
  wire u_cla32_and40;
  wire u_cla32_and41;
  wire u_cla32_or19;
  wire u_cla32_or20;
  wire u_cla32_or21;
  wire u_cla32_pg_logic11_or0;
  wire u_cla32_pg_logic11_and0;
  wire u_cla32_pg_logic11_xor0;
  wire u_cla32_xor11;
  wire u_cla32_and42;
  wire u_cla32_and43;
  wire u_cla32_and44;
  wire u_cla32_and45;
  wire u_cla32_and46;
  wire u_cla32_and47;
  wire u_cla32_and48;
  wire u_cla32_and49;
  wire u_cla32_and50;
  wire u_cla32_and51;
  wire u_cla32_or22;
  wire u_cla32_or23;
  wire u_cla32_or24;
  wire u_cla32_or25;
  wire u_cla32_pg_logic12_or0;
  wire u_cla32_pg_logic12_and0;
  wire u_cla32_pg_logic12_xor0;
  wire u_cla32_xor12;
  wire u_cla32_and52;
  wire u_cla32_or26;
  wire u_cla32_pg_logic13_or0;
  wire u_cla32_pg_logic13_and0;
  wire u_cla32_pg_logic13_xor0;
  wire u_cla32_xor13;
  wire u_cla32_and53;
  wire u_cla32_and54;
  wire u_cla32_and55;
  wire u_cla32_or27;
  wire u_cla32_or28;
  wire u_cla32_pg_logic14_or0;
  wire u_cla32_pg_logic14_and0;
  wire u_cla32_pg_logic14_xor0;
  wire u_cla32_xor14;
  wire u_cla32_and56;
  wire u_cla32_and57;
  wire u_cla32_and58;
  wire u_cla32_and59;
  wire u_cla32_and60;
  wire u_cla32_and61;
  wire u_cla32_or29;
  wire u_cla32_or30;
  wire u_cla32_or31;
  wire u_cla32_pg_logic15_or0;
  wire u_cla32_pg_logic15_and0;
  wire u_cla32_pg_logic15_xor0;
  wire u_cla32_xor15;
  wire u_cla32_and62;
  wire u_cla32_and63;
  wire u_cla32_and64;
  wire u_cla32_and65;
  wire u_cla32_and66;
  wire u_cla32_and67;
  wire u_cla32_and68;
  wire u_cla32_and69;
  wire u_cla32_and70;
  wire u_cla32_and71;
  wire u_cla32_or32;
  wire u_cla32_or33;
  wire u_cla32_or34;
  wire u_cla32_or35;
  wire u_cla32_pg_logic16_or0;
  wire u_cla32_pg_logic16_and0;
  wire u_cla32_pg_logic16_xor0;
  wire u_cla32_xor16;
  wire u_cla32_and72;
  wire u_cla32_or36;
  wire u_cla32_pg_logic17_or0;
  wire u_cla32_pg_logic17_and0;
  wire u_cla32_pg_logic17_xor0;
  wire u_cla32_xor17;
  wire u_cla32_and73;
  wire u_cla32_and74;
  wire u_cla32_and75;
  wire u_cla32_or37;
  wire u_cla32_or38;
  wire u_cla32_pg_logic18_or0;
  wire u_cla32_pg_logic18_and0;
  wire u_cla32_pg_logic18_xor0;
  wire u_cla32_xor18;
  wire u_cla32_and76;
  wire u_cla32_and77;
  wire u_cla32_and78;
  wire u_cla32_and79;
  wire u_cla32_and80;
  wire u_cla32_and81;
  wire u_cla32_or39;
  wire u_cla32_or40;
  wire u_cla32_or41;
  wire u_cla32_pg_logic19_or0;
  wire u_cla32_pg_logic19_and0;
  wire u_cla32_pg_logic19_xor0;
  wire u_cla32_xor19;
  wire u_cla32_and82;
  wire u_cla32_and83;
  wire u_cla32_and84;
  wire u_cla32_and85;
  wire u_cla32_and86;
  wire u_cla32_and87;
  wire u_cla32_and88;
  wire u_cla32_and89;
  wire u_cla32_and90;
  wire u_cla32_and91;
  wire u_cla32_or42;
  wire u_cla32_or43;
  wire u_cla32_or44;
  wire u_cla32_or45;
  wire u_cla32_pg_logic20_or0;
  wire u_cla32_pg_logic20_and0;
  wire u_cla32_pg_logic20_xor0;
  wire u_cla32_xor20;
  wire u_cla32_and92;
  wire u_cla32_or46;
  wire u_cla32_pg_logic21_or0;
  wire u_cla32_pg_logic21_and0;
  wire u_cla32_pg_logic21_xor0;
  wire u_cla32_xor21;
  wire u_cla32_and93;
  wire u_cla32_and94;
  wire u_cla32_and95;
  wire u_cla32_or47;
  wire u_cla32_or48;
  wire u_cla32_pg_logic22_or0;
  wire u_cla32_pg_logic22_and0;
  wire u_cla32_pg_logic22_xor0;
  wire u_cla32_xor22;
  wire u_cla32_and96;
  wire u_cla32_and97;
  wire u_cla32_and98;
  wire u_cla32_and99;
  wire u_cla32_and100;
  wire u_cla32_and101;
  wire u_cla32_or49;
  wire u_cla32_or50;
  wire u_cla32_or51;
  wire u_cla32_pg_logic23_or0;
  wire u_cla32_pg_logic23_and0;
  wire u_cla32_pg_logic23_xor0;
  wire u_cla32_xor23;
  wire u_cla32_and102;
  wire u_cla32_and103;
  wire u_cla32_and104;
  wire u_cla32_and105;
  wire u_cla32_and106;
  wire u_cla32_and107;
  wire u_cla32_and108;
  wire u_cla32_and109;
  wire u_cla32_and110;
  wire u_cla32_and111;
  wire u_cla32_or52;
  wire u_cla32_or53;
  wire u_cla32_or54;
  wire u_cla32_or55;
  wire u_cla32_pg_logic24_or0;
  wire u_cla32_pg_logic24_and0;
  wire u_cla32_pg_logic24_xor0;
  wire u_cla32_xor24;
  wire u_cla32_and112;
  wire u_cla32_or56;
  wire u_cla32_pg_logic25_or0;
  wire u_cla32_pg_logic25_and0;
  wire u_cla32_pg_logic25_xor0;
  wire u_cla32_xor25;
  wire u_cla32_and113;
  wire u_cla32_and114;
  wire u_cla32_and115;
  wire u_cla32_or57;
  wire u_cla32_or58;
  wire u_cla32_pg_logic26_or0;
  wire u_cla32_pg_logic26_and0;
  wire u_cla32_pg_logic26_xor0;
  wire u_cla32_xor26;
  wire u_cla32_and116;
  wire u_cla32_and117;
  wire u_cla32_and118;
  wire u_cla32_and119;
  wire u_cla32_and120;
  wire u_cla32_and121;
  wire u_cla32_or59;
  wire u_cla32_or60;
  wire u_cla32_or61;
  wire u_cla32_pg_logic27_or0;
  wire u_cla32_pg_logic27_and0;
  wire u_cla32_pg_logic27_xor0;
  wire u_cla32_xor27;
  wire u_cla32_and122;
  wire u_cla32_and123;
  wire u_cla32_and124;
  wire u_cla32_and125;
  wire u_cla32_and126;
  wire u_cla32_and127;
  wire u_cla32_and128;
  wire u_cla32_and129;
  wire u_cla32_and130;
  wire u_cla32_and131;
  wire u_cla32_or62;
  wire u_cla32_or63;
  wire u_cla32_or64;
  wire u_cla32_or65;
  wire u_cla32_pg_logic28_or0;
  wire u_cla32_pg_logic28_and0;
  wire u_cla32_pg_logic28_xor0;
  wire u_cla32_xor28;
  wire u_cla32_and132;
  wire u_cla32_or66;
  wire u_cla32_pg_logic29_or0;
  wire u_cla32_pg_logic29_and0;
  wire u_cla32_pg_logic29_xor0;
  wire u_cla32_xor29;
  wire u_cla32_and133;
  wire u_cla32_and134;
  wire u_cla32_and135;
  wire u_cla32_or67;
  wire u_cla32_or68;
  wire u_cla32_pg_logic30_or0;
  wire u_cla32_pg_logic30_and0;
  wire u_cla32_pg_logic30_xor0;
  wire u_cla32_xor30;
  wire u_cla32_and136;
  wire u_cla32_and137;
  wire u_cla32_and138;
  wire u_cla32_and139;
  wire u_cla32_and140;
  wire u_cla32_and141;
  wire u_cla32_or69;
  wire u_cla32_or70;
  wire u_cla32_or71;
  wire u_cla32_pg_logic31_or0;
  wire u_cla32_pg_logic31_and0;
  wire u_cla32_pg_logic31_xor0;
  wire u_cla32_xor31;
  wire u_cla32_and142;
  wire u_cla32_and143;
  wire u_cla32_and144;
  wire u_cla32_and145;
  wire u_cla32_and146;
  wire u_cla32_and147;
  wire u_cla32_and148;
  wire u_cla32_and149;
  wire u_cla32_and150;
  wire u_cla32_and151;
  wire u_cla32_or72;
  wire u_cla32_or73;
  wire u_cla32_or74;
  wire u_cla32_or75;

  assign u_cla32_pg_logic0_or0 = a[0] | b[0];
  assign u_cla32_pg_logic0_and0 = a[0] & b[0];
  assign u_cla32_pg_logic0_xor0 = a[0] ^ b[0];
  assign u_cla32_pg_logic1_or0 = a[1] | b[1];
  assign u_cla32_pg_logic1_and0 = a[1] & b[1];
  assign u_cla32_pg_logic1_xor0 = a[1] ^ b[1];
  assign u_cla32_xor1 = u_cla32_pg_logic1_xor0 ^ u_cla32_pg_logic0_and0;
  assign u_cla32_and0 = u_cla32_pg_logic0_and0 & u_cla32_pg_logic1_or0;
  assign u_cla32_or0 = u_cla32_pg_logic1_and0 | u_cla32_and0;
  assign u_cla32_pg_logic2_or0 = a[2] | b[2];
  assign u_cla32_pg_logic2_and0 = a[2] & b[2];
  assign u_cla32_pg_logic2_xor0 = a[2] ^ b[2];
  assign u_cla32_xor2 = u_cla32_pg_logic2_xor0 ^ u_cla32_or0;
  assign u_cla32_and1 = u_cla32_pg_logic2_or0 & u_cla32_pg_logic0_or0;
  assign u_cla32_and2 = u_cla32_pg_logic0_and0 & u_cla32_pg_logic2_or0;
  assign u_cla32_and3 = u_cla32_and2 & u_cla32_pg_logic1_or0;
  assign u_cla32_and4 = u_cla32_pg_logic1_and0 & u_cla32_pg_logic2_or0;
  assign u_cla32_or1 = u_cla32_and3 | u_cla32_and4;
  assign u_cla32_or2 = u_cla32_pg_logic2_and0 | u_cla32_or1;
  assign u_cla32_pg_logic3_or0 = a[3] | b[3];
  assign u_cla32_pg_logic3_and0 = a[3] & b[3];
  assign u_cla32_pg_logic3_xor0 = a[3] ^ b[3];
  assign u_cla32_xor3 = u_cla32_pg_logic3_xor0 ^ u_cla32_or2;
  assign u_cla32_and5 = u_cla32_pg_logic3_or0 & u_cla32_pg_logic1_or0;
  assign u_cla32_and6 = u_cla32_pg_logic0_and0 & u_cla32_pg_logic2_or0;
  assign u_cla32_and7 = u_cla32_pg_logic3_or0 & u_cla32_pg_logic1_or0;
  assign u_cla32_and8 = u_cla32_and6 & u_cla32_and7;
  assign u_cla32_and9 = u_cla32_pg_logic1_and0 & u_cla32_pg_logic3_or0;
  assign u_cla32_and10 = u_cla32_and9 & u_cla32_pg_logic2_or0;
  assign u_cla32_and11 = u_cla32_pg_logic2_and0 & u_cla32_pg_logic3_or0;
  assign u_cla32_or3 = u_cla32_and8 | u_cla32_and11;
  assign u_cla32_or4 = u_cla32_and10 | u_cla32_or3;
  assign u_cla32_or5 = u_cla32_pg_logic3_and0 | u_cla32_or4;
  assign u_cla32_pg_logic4_or0 = a[4] | b[4];
  assign u_cla32_pg_logic4_and0 = a[4] & b[4];
  assign u_cla32_pg_logic4_xor0 = a[4] ^ b[4];
  assign u_cla32_xor4 = u_cla32_pg_logic4_xor0 ^ u_cla32_or5;
  assign u_cla32_and12 = u_cla32_or5 & u_cla32_pg_logic4_or0;
  assign u_cla32_or6 = u_cla32_pg_logic4_and0 | u_cla32_and12;
  assign u_cla32_pg_logic5_or0 = a[5] | b[5];
  assign u_cla32_pg_logic5_and0 = a[5] & b[5];
  assign u_cla32_pg_logic5_xor0 = a[5] ^ b[5];
  assign u_cla32_xor5 = u_cla32_pg_logic5_xor0 ^ u_cla32_or6;
  assign u_cla32_and13 = u_cla32_or5 & u_cla32_pg_logic5_or0;
  assign u_cla32_and14 = u_cla32_and13 & u_cla32_pg_logic4_or0;
  assign u_cla32_and15 = u_cla32_pg_logic4_and0 & u_cla32_pg_logic5_or0;
  assign u_cla32_or7 = u_cla32_and14 | u_cla32_and15;
  assign u_cla32_or8 = u_cla32_pg_logic5_and0 | u_cla32_or7;
  assign u_cla32_pg_logic6_or0 = a[6] | b[6];
  assign u_cla32_pg_logic6_and0 = a[6] & b[6];
  assign u_cla32_pg_logic6_xor0 = a[6] ^ b[6];
  assign u_cla32_xor6 = u_cla32_pg_logic6_xor0 ^ u_cla32_or8;
  assign u_cla32_and16 = u_cla32_or5 & u_cla32_pg_logic5_or0;
  assign u_cla32_and17 = u_cla32_pg_logic6_or0 & u_cla32_pg_logic4_or0;
  assign u_cla32_and18 = u_cla32_and16 & u_cla32_and17;
  assign u_cla32_and19 = u_cla32_pg_logic4_and0 & u_cla32_pg_logic6_or0;
  assign u_cla32_and20 = u_cla32_and19 & u_cla32_pg_logic5_or0;
  assign u_cla32_and21 = u_cla32_pg_logic5_and0 & u_cla32_pg_logic6_or0;
  assign u_cla32_or9 = u_cla32_and18 | u_cla32_and20;
  assign u_cla32_or10 = u_cla32_or9 | u_cla32_and21;
  assign u_cla32_or11 = u_cla32_pg_logic6_and0 | u_cla32_or10;
  assign u_cla32_pg_logic7_or0 = a[7] | b[7];
  assign u_cla32_pg_logic7_and0 = a[7] & b[7];
  assign u_cla32_pg_logic7_xor0 = a[7] ^ b[7];
  assign u_cla32_xor7 = u_cla32_pg_logic7_xor0 ^ u_cla32_or11;
  assign u_cla32_and22 = u_cla32_or5 & u_cla32_pg_logic6_or0;
  assign u_cla32_and23 = u_cla32_pg_logic7_or0 & u_cla32_pg_logic5_or0;
  assign u_cla32_and24 = u_cla32_and22 & u_cla32_and23;
  assign u_cla32_and25 = u_cla32_and24 & u_cla32_pg_logic4_or0;
  assign u_cla32_and26 = u_cla32_pg_logic4_and0 & u_cla32_pg_logic6_or0;
  assign u_cla32_and27 = u_cla32_pg_logic7_or0 & u_cla32_pg_logic5_or0;
  assign u_cla32_and28 = u_cla32_and26 & u_cla32_and27;
  assign u_cla32_and29 = u_cla32_pg_logic5_and0 & u_cla32_pg_logic7_or0;
  assign u_cla32_and30 = u_cla32_and29 & u_cla32_pg_logic6_or0;
  assign u_cla32_and31 = u_cla32_pg_logic6_and0 & u_cla32_pg_logic7_or0;
  assign u_cla32_or12 = u_cla32_and25 | u_cla32_and30;
  assign u_cla32_or13 = u_cla32_and28 | u_cla32_and31;
  assign u_cla32_or14 = u_cla32_or12 | u_cla32_or13;
  assign u_cla32_or15 = u_cla32_pg_logic7_and0 | u_cla32_or14;
  assign u_cla32_pg_logic8_or0 = a[8] | b[8];
  assign u_cla32_pg_logic8_and0 = a[8] & b[8];
  assign u_cla32_pg_logic8_xor0 = a[8] ^ b[8];
  assign u_cla32_xor8 = u_cla32_pg_logic8_xor0 ^ u_cla32_or15;
  assign u_cla32_and32 = u_cla32_or15 & u_cla32_pg_logic8_or0;
  assign u_cla32_or16 = u_cla32_pg_logic8_and0 | u_cla32_and32;
  assign u_cla32_pg_logic9_or0 = a[9] | b[9];
  assign u_cla32_pg_logic9_and0 = a[9] & b[9];
  assign u_cla32_pg_logic9_xor0 = a[9] ^ b[9];
  assign u_cla32_xor9 = u_cla32_pg_logic9_xor0 ^ u_cla32_or16;
  assign u_cla32_and33 = u_cla32_or15 & u_cla32_pg_logic9_or0;
  assign u_cla32_and34 = u_cla32_and33 & u_cla32_pg_logic8_or0;
  assign u_cla32_and35 = u_cla32_pg_logic8_and0 & u_cla32_pg_logic9_or0;
  assign u_cla32_or17 = u_cla32_and34 | u_cla32_and35;
  assign u_cla32_or18 = u_cla32_pg_logic9_and0 | u_cla32_or17;
  assign u_cla32_pg_logic10_or0 = a[10] | b[10];
  assign u_cla32_pg_logic10_and0 = a[10] & b[10];
  assign u_cla32_pg_logic10_xor0 = a[10] ^ b[10];
  assign u_cla32_xor10 = u_cla32_pg_logic10_xor0 ^ u_cla32_or18;
  assign u_cla32_and36 = u_cla32_or15 & u_cla32_pg_logic9_or0;
  assign u_cla32_and37 = u_cla32_pg_logic10_or0 & u_cla32_pg_logic8_or0;
  assign u_cla32_and38 = u_cla32_and36 & u_cla32_and37;
  assign u_cla32_and39 = u_cla32_pg_logic8_and0 & u_cla32_pg_logic10_or0;
  assign u_cla32_and40 = u_cla32_and39 & u_cla32_pg_logic9_or0;
  assign u_cla32_and41 = u_cla32_pg_logic9_and0 & u_cla32_pg_logic10_or0;
  assign u_cla32_or19 = u_cla32_and38 | u_cla32_and40;
  assign u_cla32_or20 = u_cla32_or19 | u_cla32_and41;
  assign u_cla32_or21 = u_cla32_pg_logic10_and0 | u_cla32_or20;
  assign u_cla32_pg_logic11_or0 = a[11] | b[11];
  assign u_cla32_pg_logic11_and0 = a[11] & b[11];
  assign u_cla32_pg_logic11_xor0 = a[11] ^ b[11];
  assign u_cla32_xor11 = u_cla32_pg_logic11_xor0 ^ u_cla32_or21;
  assign u_cla32_and42 = u_cla32_or15 & u_cla32_pg_logic10_or0;
  assign u_cla32_and43 = u_cla32_pg_logic11_or0 & u_cla32_pg_logic9_or0;
  assign u_cla32_and44 = u_cla32_and42 & u_cla32_and43;
  assign u_cla32_and45 = u_cla32_and44 & u_cla32_pg_logic8_or0;
  assign u_cla32_and46 = u_cla32_pg_logic8_and0 & u_cla32_pg_logic10_or0;
  assign u_cla32_and47 = u_cla32_pg_logic11_or0 & u_cla32_pg_logic9_or0;
  assign u_cla32_and48 = u_cla32_and46 & u_cla32_and47;
  assign u_cla32_and49 = u_cla32_pg_logic9_and0 & u_cla32_pg_logic11_or0;
  assign u_cla32_and50 = u_cla32_and49 & u_cla32_pg_logic10_or0;
  assign u_cla32_and51 = u_cla32_pg_logic10_and0 & u_cla32_pg_logic11_or0;
  assign u_cla32_or22 = u_cla32_and45 | u_cla32_and50;
  assign u_cla32_or23 = u_cla32_and48 | u_cla32_and51;
  assign u_cla32_or24 = u_cla32_or22 | u_cla32_or23;
  assign u_cla32_or25 = u_cla32_pg_logic11_and0 | u_cla32_or24;
  assign u_cla32_pg_logic12_or0 = a[12] | b[12];
  assign u_cla32_pg_logic12_and0 = a[12] & b[12];
  assign u_cla32_pg_logic12_xor0 = a[12] ^ b[12];
  assign u_cla32_xor12 = u_cla32_pg_logic12_xor0 ^ u_cla32_or25;
  assign u_cla32_and52 = u_cla32_or25 & u_cla32_pg_logic12_or0;
  assign u_cla32_or26 = u_cla32_pg_logic12_and0 | u_cla32_and52;
  assign u_cla32_pg_logic13_or0 = a[13] | b[13];
  assign u_cla32_pg_logic13_and0 = a[13] & b[13];
  assign u_cla32_pg_logic13_xor0 = a[13] ^ b[13];
  assign u_cla32_xor13 = u_cla32_pg_logic13_xor0 ^ u_cla32_or26;
  assign u_cla32_and53 = u_cla32_or25 & u_cla32_pg_logic13_or0;
  assign u_cla32_and54 = u_cla32_and53 & u_cla32_pg_logic12_or0;
  assign u_cla32_and55 = u_cla32_pg_logic12_and0 & u_cla32_pg_logic13_or0;
  assign u_cla32_or27 = u_cla32_and54 | u_cla32_and55;
  assign u_cla32_or28 = u_cla32_pg_logic13_and0 | u_cla32_or27;
  assign u_cla32_pg_logic14_or0 = a[14] | b[14];
  assign u_cla32_pg_logic14_and0 = a[14] & b[14];
  assign u_cla32_pg_logic14_xor0 = a[14] ^ b[14];
  assign u_cla32_xor14 = u_cla32_pg_logic14_xor0 ^ u_cla32_or28;
  assign u_cla32_and56 = u_cla32_or25 & u_cla32_pg_logic13_or0;
  assign u_cla32_and57 = u_cla32_pg_logic14_or0 & u_cla32_pg_logic12_or0;
  assign u_cla32_and58 = u_cla32_and56 & u_cla32_and57;
  assign u_cla32_and59 = u_cla32_pg_logic12_and0 & u_cla32_pg_logic14_or0;
  assign u_cla32_and60 = u_cla32_and59 & u_cla32_pg_logic13_or0;
  assign u_cla32_and61 = u_cla32_pg_logic13_and0 & u_cla32_pg_logic14_or0;
  assign u_cla32_or29 = u_cla32_and58 | u_cla32_and60;
  assign u_cla32_or30 = u_cla32_or29 | u_cla32_and61;
  assign u_cla32_or31 = u_cla32_pg_logic14_and0 | u_cla32_or30;
  assign u_cla32_pg_logic15_or0 = a[15] | b[15];
  assign u_cla32_pg_logic15_and0 = a[15] & b[15];
  assign u_cla32_pg_logic15_xor0 = a[15] ^ b[15];
  assign u_cla32_xor15 = u_cla32_pg_logic15_xor0 ^ u_cla32_or31;
  assign u_cla32_and62 = u_cla32_or25 & u_cla32_pg_logic14_or0;
  assign u_cla32_and63 = u_cla32_pg_logic15_or0 & u_cla32_pg_logic13_or0;
  assign u_cla32_and64 = u_cla32_and62 & u_cla32_and63;
  assign u_cla32_and65 = u_cla32_and64 & u_cla32_pg_logic12_or0;
  assign u_cla32_and66 = u_cla32_pg_logic12_and0 & u_cla32_pg_logic14_or0;
  assign u_cla32_and67 = u_cla32_pg_logic15_or0 & u_cla32_pg_logic13_or0;
  assign u_cla32_and68 = u_cla32_and66 & u_cla32_and67;
  assign u_cla32_and69 = u_cla32_pg_logic13_and0 & u_cla32_pg_logic15_or0;
  assign u_cla32_and70 = u_cla32_and69 & u_cla32_pg_logic14_or0;
  assign u_cla32_and71 = u_cla32_pg_logic14_and0 & u_cla32_pg_logic15_or0;
  assign u_cla32_or32 = u_cla32_and65 | u_cla32_and70;
  assign u_cla32_or33 = u_cla32_and68 | u_cla32_and71;
  assign u_cla32_or34 = u_cla32_or32 | u_cla32_or33;
  assign u_cla32_or35 = u_cla32_pg_logic15_and0 | u_cla32_or34;
  assign u_cla32_pg_logic16_or0 = a[16] | b[16];
  assign u_cla32_pg_logic16_and0 = a[16] & b[16];
  assign u_cla32_pg_logic16_xor0 = a[16] ^ b[16];
  assign u_cla32_xor16 = u_cla32_pg_logic16_xor0 ^ u_cla32_or35;
  assign u_cla32_and72 = u_cla32_or35 & u_cla32_pg_logic16_or0;
  assign u_cla32_or36 = u_cla32_pg_logic16_and0 | u_cla32_and72;
  assign u_cla32_pg_logic17_or0 = a[17] | b[17];
  assign u_cla32_pg_logic17_and0 = a[17] & b[17];
  assign u_cla32_pg_logic17_xor0 = a[17] ^ b[17];
  assign u_cla32_xor17 = u_cla32_pg_logic17_xor0 ^ u_cla32_or36;
  assign u_cla32_and73 = u_cla32_or35 & u_cla32_pg_logic17_or0;
  assign u_cla32_and74 = u_cla32_and73 & u_cla32_pg_logic16_or0;
  assign u_cla32_and75 = u_cla32_pg_logic16_and0 & u_cla32_pg_logic17_or0;
  assign u_cla32_or37 = u_cla32_and74 | u_cla32_and75;
  assign u_cla32_or38 = u_cla32_pg_logic17_and0 | u_cla32_or37;
  assign u_cla32_pg_logic18_or0 = a[18] | b[18];
  assign u_cla32_pg_logic18_and0 = a[18] & b[18];
  assign u_cla32_pg_logic18_xor0 = a[18] ^ b[18];
  assign u_cla32_xor18 = u_cla32_pg_logic18_xor0 ^ u_cla32_or38;
  assign u_cla32_and76 = u_cla32_or35 & u_cla32_pg_logic17_or0;
  assign u_cla32_and77 = u_cla32_pg_logic18_or0 & u_cla32_pg_logic16_or0;
  assign u_cla32_and78 = u_cla32_and76 & u_cla32_and77;
  assign u_cla32_and79 = u_cla32_pg_logic16_and0 & u_cla32_pg_logic18_or0;
  assign u_cla32_and80 = u_cla32_and79 & u_cla32_pg_logic17_or0;
  assign u_cla32_and81 = u_cla32_pg_logic17_and0 & u_cla32_pg_logic18_or0;
  assign u_cla32_or39 = u_cla32_and78 | u_cla32_and80;
  assign u_cla32_or40 = u_cla32_or39 | u_cla32_and81;
  assign u_cla32_or41 = u_cla32_pg_logic18_and0 | u_cla32_or40;
  assign u_cla32_pg_logic19_or0 = a[19] | b[19];
  assign u_cla32_pg_logic19_and0 = a[19] & b[19];
  assign u_cla32_pg_logic19_xor0 = a[19] ^ b[19];
  assign u_cla32_xor19 = u_cla32_pg_logic19_xor0 ^ u_cla32_or41;
  assign u_cla32_and82 = u_cla32_or35 & u_cla32_pg_logic18_or0;
  assign u_cla32_and83 = u_cla32_pg_logic19_or0 & u_cla32_pg_logic17_or0;
  assign u_cla32_and84 = u_cla32_and82 & u_cla32_and83;
  assign u_cla32_and85 = u_cla32_and84 & u_cla32_pg_logic16_or0;
  assign u_cla32_and86 = u_cla32_pg_logic16_and0 & u_cla32_pg_logic18_or0;
  assign u_cla32_and87 = u_cla32_pg_logic19_or0 & u_cla32_pg_logic17_or0;
  assign u_cla32_and88 = u_cla32_and86 & u_cla32_and87;
  assign u_cla32_and89 = u_cla32_pg_logic17_and0 & u_cla32_pg_logic19_or0;
  assign u_cla32_and90 = u_cla32_and89 & u_cla32_pg_logic18_or0;
  assign u_cla32_and91 = u_cla32_pg_logic18_and0 & u_cla32_pg_logic19_or0;
  assign u_cla32_or42 = u_cla32_and85 | u_cla32_and90;
  assign u_cla32_or43 = u_cla32_and88 | u_cla32_and91;
  assign u_cla32_or44 = u_cla32_or42 | u_cla32_or43;
  assign u_cla32_or45 = u_cla32_pg_logic19_and0 | u_cla32_or44;
  assign u_cla32_pg_logic20_or0 = a[20] | b[20];
  assign u_cla32_pg_logic20_and0 = a[20] & b[20];
  assign u_cla32_pg_logic20_xor0 = a[20] ^ b[20];
  assign u_cla32_xor20 = u_cla32_pg_logic20_xor0 ^ u_cla32_or45;
  assign u_cla32_and92 = u_cla32_or45 & u_cla32_pg_logic20_or0;
  assign u_cla32_or46 = u_cla32_pg_logic20_and0 | u_cla32_and92;
  assign u_cla32_pg_logic21_or0 = a[21] | b[21];
  assign u_cla32_pg_logic21_and0 = a[21] & b[21];
  assign u_cla32_pg_logic21_xor0 = a[21] ^ b[21];
  assign u_cla32_xor21 = u_cla32_pg_logic21_xor0 ^ u_cla32_or46;
  assign u_cla32_and93 = u_cla32_or45 & u_cla32_pg_logic21_or0;
  assign u_cla32_and94 = u_cla32_and93 & u_cla32_pg_logic20_or0;
  assign u_cla32_and95 = u_cla32_pg_logic20_and0 & u_cla32_pg_logic21_or0;
  assign u_cla32_or47 = u_cla32_and94 | u_cla32_and95;
  assign u_cla32_or48 = u_cla32_pg_logic21_and0 | u_cla32_or47;
  assign u_cla32_pg_logic22_or0 = a[22] | b[22];
  assign u_cla32_pg_logic22_and0 = a[22] & b[22];
  assign u_cla32_pg_logic22_xor0 = a[22] ^ b[22];
  assign u_cla32_xor22 = u_cla32_pg_logic22_xor0 ^ u_cla32_or48;
  assign u_cla32_and96 = u_cla32_or45 & u_cla32_pg_logic21_or0;
  assign u_cla32_and97 = u_cla32_pg_logic22_or0 & u_cla32_pg_logic20_or0;
  assign u_cla32_and98 = u_cla32_and96 & u_cla32_and97;
  assign u_cla32_and99 = u_cla32_pg_logic20_and0 & u_cla32_pg_logic22_or0;
  assign u_cla32_and100 = u_cla32_and99 & u_cla32_pg_logic21_or0;
  assign u_cla32_and101 = u_cla32_pg_logic21_and0 & u_cla32_pg_logic22_or0;
  assign u_cla32_or49 = u_cla32_and98 | u_cla32_and100;
  assign u_cla32_or50 = u_cla32_or49 | u_cla32_and101;
  assign u_cla32_or51 = u_cla32_pg_logic22_and0 | u_cla32_or50;
  assign u_cla32_pg_logic23_or0 = a[23] | b[23];
  assign u_cla32_pg_logic23_and0 = a[23] & b[23];
  assign u_cla32_pg_logic23_xor0 = a[23] ^ b[23];
  assign u_cla32_xor23 = u_cla32_pg_logic23_xor0 ^ u_cla32_or51;
  assign u_cla32_and102 = u_cla32_or45 & u_cla32_pg_logic22_or0;
  assign u_cla32_and103 = u_cla32_pg_logic23_or0 & u_cla32_pg_logic21_or0;
  assign u_cla32_and104 = u_cla32_and102 & u_cla32_and103;
  assign u_cla32_and105 = u_cla32_and104 & u_cla32_pg_logic20_or0;
  assign u_cla32_and106 = u_cla32_pg_logic20_and0 & u_cla32_pg_logic22_or0;
  assign u_cla32_and107 = u_cla32_pg_logic23_or0 & u_cla32_pg_logic21_or0;
  assign u_cla32_and108 = u_cla32_and106 & u_cla32_and107;
  assign u_cla32_and109 = u_cla32_pg_logic21_and0 & u_cla32_pg_logic23_or0;
  assign u_cla32_and110 = u_cla32_and109 & u_cla32_pg_logic22_or0;
  assign u_cla32_and111 = u_cla32_pg_logic22_and0 & u_cla32_pg_logic23_or0;
  assign u_cla32_or52 = u_cla32_and105 | u_cla32_and110;
  assign u_cla32_or53 = u_cla32_and108 | u_cla32_and111;
  assign u_cla32_or54 = u_cla32_or52 | u_cla32_or53;
  assign u_cla32_or55 = u_cla32_pg_logic23_and0 | u_cla32_or54;
  assign u_cla32_pg_logic24_or0 = a[24] | b[24];
  assign u_cla32_pg_logic24_and0 = a[24] & b[24];
  assign u_cla32_pg_logic24_xor0 = a[24] ^ b[24];
  assign u_cla32_xor24 = u_cla32_pg_logic24_xor0 ^ u_cla32_or55;
  assign u_cla32_and112 = u_cla32_or55 & u_cla32_pg_logic24_or0;
  assign u_cla32_or56 = u_cla32_pg_logic24_and0 | u_cla32_and112;
  assign u_cla32_pg_logic25_or0 = a[25] | b[25];
  assign u_cla32_pg_logic25_and0 = a[25] & b[25];
  assign u_cla32_pg_logic25_xor0 = a[25] ^ b[25];
  assign u_cla32_xor25 = u_cla32_pg_logic25_xor0 ^ u_cla32_or56;
  assign u_cla32_and113 = u_cla32_or55 & u_cla32_pg_logic25_or0;
  assign u_cla32_and114 = u_cla32_and113 & u_cla32_pg_logic24_or0;
  assign u_cla32_and115 = u_cla32_pg_logic24_and0 & u_cla32_pg_logic25_or0;
  assign u_cla32_or57 = u_cla32_and114 | u_cla32_and115;
  assign u_cla32_or58 = u_cla32_pg_logic25_and0 | u_cla32_or57;
  assign u_cla32_pg_logic26_or0 = a[26] | b[26];
  assign u_cla32_pg_logic26_and0 = a[26] & b[26];
  assign u_cla32_pg_logic26_xor0 = a[26] ^ b[26];
  assign u_cla32_xor26 = u_cla32_pg_logic26_xor0 ^ u_cla32_or58;
  assign u_cla32_and116 = u_cla32_or55 & u_cla32_pg_logic25_or0;
  assign u_cla32_and117 = u_cla32_pg_logic26_or0 & u_cla32_pg_logic24_or0;
  assign u_cla32_and118 = u_cla32_and116 & u_cla32_and117;
  assign u_cla32_and119 = u_cla32_pg_logic24_and0 & u_cla32_pg_logic26_or0;
  assign u_cla32_and120 = u_cla32_and119 & u_cla32_pg_logic25_or0;
  assign u_cla32_and121 = u_cla32_pg_logic25_and0 & u_cla32_pg_logic26_or0;
  assign u_cla32_or59 = u_cla32_and118 | u_cla32_and120;
  assign u_cla32_or60 = u_cla32_or59 | u_cla32_and121;
  assign u_cla32_or61 = u_cla32_pg_logic26_and0 | u_cla32_or60;
  assign u_cla32_pg_logic27_or0 = a[27] | b[27];
  assign u_cla32_pg_logic27_and0 = a[27] & b[27];
  assign u_cla32_pg_logic27_xor0 = a[27] ^ b[27];
  assign u_cla32_xor27 = u_cla32_pg_logic27_xor0 ^ u_cla32_or61;
  assign u_cla32_and122 = u_cla32_or55 & u_cla32_pg_logic26_or0;
  assign u_cla32_and123 = u_cla32_pg_logic27_or0 & u_cla32_pg_logic25_or0;
  assign u_cla32_and124 = u_cla32_and122 & u_cla32_and123;
  assign u_cla32_and125 = u_cla32_and124 & u_cla32_pg_logic24_or0;
  assign u_cla32_and126 = u_cla32_pg_logic24_and0 & u_cla32_pg_logic26_or0;
  assign u_cla32_and127 = u_cla32_pg_logic27_or0 & u_cla32_pg_logic25_or0;
  assign u_cla32_and128 = u_cla32_and126 & u_cla32_and127;
  assign u_cla32_and129 = u_cla32_pg_logic25_and0 & u_cla32_pg_logic27_or0;
  assign u_cla32_and130 = u_cla32_and129 & u_cla32_pg_logic26_or0;
  assign u_cla32_and131 = u_cla32_pg_logic26_and0 & u_cla32_pg_logic27_or0;
  assign u_cla32_or62 = u_cla32_and125 | u_cla32_and130;
  assign u_cla32_or63 = u_cla32_and128 | u_cla32_and131;
  assign u_cla32_or64 = u_cla32_or62 | u_cla32_or63;
  assign u_cla32_or65 = u_cla32_pg_logic27_and0 | u_cla32_or64;
  assign u_cla32_pg_logic28_or0 = a[28] | b[28];
  assign u_cla32_pg_logic28_and0 = a[28] & b[28];
  assign u_cla32_pg_logic28_xor0 = a[28] ^ b[28];
  assign u_cla32_xor28 = u_cla32_pg_logic28_xor0 ^ u_cla32_or65;
  assign u_cla32_and132 = u_cla32_or65 & u_cla32_pg_logic28_or0;
  assign u_cla32_or66 = u_cla32_pg_logic28_and0 | u_cla32_and132;
  assign u_cla32_pg_logic29_or0 = a[29] | b[29];
  assign u_cla32_pg_logic29_and0 = a[29] & b[29];
  assign u_cla32_pg_logic29_xor0 = a[29] ^ b[29];
  assign u_cla32_xor29 = u_cla32_pg_logic29_xor0 ^ u_cla32_or66;
  assign u_cla32_and133 = u_cla32_or65 & u_cla32_pg_logic29_or0;
  assign u_cla32_and134 = u_cla32_and133 & u_cla32_pg_logic28_or0;
  assign u_cla32_and135 = u_cla32_pg_logic28_and0 & u_cla32_pg_logic29_or0;
  assign u_cla32_or67 = u_cla32_and134 | u_cla32_and135;
  assign u_cla32_or68 = u_cla32_pg_logic29_and0 | u_cla32_or67;
  assign u_cla32_pg_logic30_or0 = a[30] | b[30];
  assign u_cla32_pg_logic30_and0 = a[30] & b[30];
  assign u_cla32_pg_logic30_xor0 = a[30] ^ b[30];
  assign u_cla32_xor30 = u_cla32_pg_logic30_xor0 ^ u_cla32_or68;
  assign u_cla32_and136 = u_cla32_or65 & u_cla32_pg_logic29_or0;
  assign u_cla32_and137 = u_cla32_pg_logic30_or0 & u_cla32_pg_logic28_or0;
  assign u_cla32_and138 = u_cla32_and136 & u_cla32_and137;
  assign u_cla32_and139 = u_cla32_pg_logic28_and0 & u_cla32_pg_logic30_or0;
  assign u_cla32_and140 = u_cla32_and139 & u_cla32_pg_logic29_or0;
  assign u_cla32_and141 = u_cla32_pg_logic29_and0 & u_cla32_pg_logic30_or0;
  assign u_cla32_or69 = u_cla32_and138 | u_cla32_and140;
  assign u_cla32_or70 = u_cla32_or69 | u_cla32_and141;
  assign u_cla32_or71 = u_cla32_pg_logic30_and0 | u_cla32_or70;
  assign u_cla32_pg_logic31_or0 = a[31] | b[31];
  assign u_cla32_pg_logic31_and0 = a[31] & b[31];
  assign u_cla32_pg_logic31_xor0 = a[31] ^ b[31];
  assign u_cla32_xor31 = u_cla32_pg_logic31_xor0 ^ u_cla32_or71;
  assign u_cla32_and142 = u_cla32_or65 & u_cla32_pg_logic30_or0;
  assign u_cla32_and143 = u_cla32_pg_logic31_or0 & u_cla32_pg_logic29_or0;
  assign u_cla32_and144 = u_cla32_and142 & u_cla32_and143;
  assign u_cla32_and145 = u_cla32_and144 & u_cla32_pg_logic28_or0;
  assign u_cla32_and146 = u_cla32_pg_logic28_and0 & u_cla32_pg_logic30_or0;
  assign u_cla32_and147 = u_cla32_pg_logic31_or0 & u_cla32_pg_logic29_or0;
  assign u_cla32_and148 = u_cla32_and146 & u_cla32_and147;
  assign u_cla32_and149 = u_cla32_pg_logic29_and0 & u_cla32_pg_logic31_or0;
  assign u_cla32_and150 = u_cla32_and149 & u_cla32_pg_logic30_or0;
  assign u_cla32_and151 = u_cla32_pg_logic30_and0 & u_cla32_pg_logic31_or0;
  assign u_cla32_or72 = u_cla32_and145 | u_cla32_and150;
  assign u_cla32_or73 = u_cla32_and148 | u_cla32_and151;
  assign u_cla32_or74 = u_cla32_or72 | u_cla32_or73;
  assign u_cla32_or75 = u_cla32_pg_logic31_and0 | u_cla32_or74;

  assign u_cla32_out[0] = u_cla32_pg_logic0_xor0;
  assign u_cla32_out[1] = u_cla32_xor1;
  assign u_cla32_out[2] = u_cla32_xor2;
  assign u_cla32_out[3] = u_cla32_xor3;
  assign u_cla32_out[4] = u_cla32_xor4;
  assign u_cla32_out[5] = u_cla32_xor5;
  assign u_cla32_out[6] = u_cla32_xor6;
  assign u_cla32_out[7] = u_cla32_xor7;
  assign u_cla32_out[8] = u_cla32_xor8;
  assign u_cla32_out[9] = u_cla32_xor9;
  assign u_cla32_out[10] = u_cla32_xor10;
  assign u_cla32_out[11] = u_cla32_xor11;
  assign u_cla32_out[12] = u_cla32_xor12;
  assign u_cla32_out[13] = u_cla32_xor13;
  assign u_cla32_out[14] = u_cla32_xor14;
  assign u_cla32_out[15] = u_cla32_xor15;
  assign u_cla32_out[16] = u_cla32_xor16;
  assign u_cla32_out[17] = u_cla32_xor17;
  assign u_cla32_out[18] = u_cla32_xor18;
  assign u_cla32_out[19] = u_cla32_xor19;
  assign u_cla32_out[20] = u_cla32_xor20;
  assign u_cla32_out[21] = u_cla32_xor21;
  assign u_cla32_out[22] = u_cla32_xor22;
  assign u_cla32_out[23] = u_cla32_xor23;
  assign u_cla32_out[24] = u_cla32_xor24;
  assign u_cla32_out[25] = u_cla32_xor25;
  assign u_cla32_out[26] = u_cla32_xor26;
  assign u_cla32_out[27] = u_cla32_xor27;
  assign u_cla32_out[28] = u_cla32_xor28;
  assign u_cla32_out[29] = u_cla32_xor29;
  assign u_cla32_out[30] = u_cla32_xor30;
  assign u_cla32_out[31] = u_cla32_xor31;
  assign u_cla32_out[32] = u_cla32_or75;
endmodule