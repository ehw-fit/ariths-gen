module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module nand_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a & _b);
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  xor_gate xor_gate_ha_y0(a, b, ha_y0);
  and_gate and_gate_ha_y1(a, b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_y0;
  wire fa_y1;
  wire fa_y3;

  xor_gate xor_gate_fa_y0(a, b, fa_y0);
  and_gate and_gate_fa_y1(a, b, fa_y1);
  and_gate and_gate_fa_y3(fa_y0, cin, fa_y3);

  xor_gate xor_gate_fa_y2(fa_y0, cin, fa_y2);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module h_s_arr_mul8(input [7:0] a, input [7:0] b, output [15:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire h_s_arr_mul8_xor_constant_wire_y0;
  wire h_s_arr_mul8_xnor_constant_wire_y0;
  wire constant_wire;
  wire h_s_arr_mul8_and_0_0_y0;
  wire h_s_arr_mul8_and_1_0_y0;
  wire h_s_arr_mul8_and_2_0_y0;
  wire h_s_arr_mul8_and_3_0_y0;
  wire h_s_arr_mul8_and_4_0_y0;
  wire h_s_arr_mul8_and_5_0_y0;
  wire h_s_arr_mul8_and_6_0_y0;
  wire h_s_arr_mul8_nand_7_0_y0;
  wire h_s_arr_mul8_and_0_1_y0;
  wire h_s_arr_mul8_ha_0_1_y0;
  wire h_s_arr_mul8_ha_0_1_y1;
  wire h_s_arr_mul8_and_1_1_y0;
  wire h_s_arr_mul8_fa_1_1_y2;
  wire h_s_arr_mul8_fa_1_1_y4;
  wire h_s_arr_mul8_and_2_1_y0;
  wire h_s_arr_mul8_fa_2_1_y2;
  wire h_s_arr_mul8_fa_2_1_y4;
  wire h_s_arr_mul8_and_3_1_y0;
  wire h_s_arr_mul8_fa_3_1_y2;
  wire h_s_arr_mul8_fa_3_1_y4;
  wire h_s_arr_mul8_and_4_1_y0;
  wire h_s_arr_mul8_fa_4_1_y2;
  wire h_s_arr_mul8_fa_4_1_y4;
  wire h_s_arr_mul8_and_5_1_y0;
  wire h_s_arr_mul8_fa_5_1_y2;
  wire h_s_arr_mul8_fa_5_1_y4;
  wire h_s_arr_mul8_and_6_1_y0;
  wire h_s_arr_mul8_fa_6_1_y2;
  wire h_s_arr_mul8_fa_6_1_y4;
  wire h_s_arr_mul8_nand_7_1_y0;
  wire h_s_arr_mul8_fa_7_1_y2;
  wire h_s_arr_mul8_fa_7_1_y4;
  wire h_s_arr_mul8_and_0_2_y0;
  wire h_s_arr_mul8_ha_0_2_y0;
  wire h_s_arr_mul8_ha_0_2_y1;
  wire h_s_arr_mul8_and_1_2_y0;
  wire h_s_arr_mul8_fa_1_2_y2;
  wire h_s_arr_mul8_fa_1_2_y4;
  wire h_s_arr_mul8_and_2_2_y0;
  wire h_s_arr_mul8_fa_2_2_y2;
  wire h_s_arr_mul8_fa_2_2_y4;
  wire h_s_arr_mul8_and_3_2_y0;
  wire h_s_arr_mul8_fa_3_2_y2;
  wire h_s_arr_mul8_fa_3_2_y4;
  wire h_s_arr_mul8_and_4_2_y0;
  wire h_s_arr_mul8_fa_4_2_y2;
  wire h_s_arr_mul8_fa_4_2_y4;
  wire h_s_arr_mul8_and_5_2_y0;
  wire h_s_arr_mul8_fa_5_2_y2;
  wire h_s_arr_mul8_fa_5_2_y4;
  wire h_s_arr_mul8_and_6_2_y0;
  wire h_s_arr_mul8_fa_6_2_y2;
  wire h_s_arr_mul8_fa_6_2_y4;
  wire h_s_arr_mul8_nand_7_2_y0;
  wire h_s_arr_mul8_fa_7_2_y2;
  wire h_s_arr_mul8_fa_7_2_y4;
  wire h_s_arr_mul8_and_0_3_y0;
  wire h_s_arr_mul8_ha_0_3_y0;
  wire h_s_arr_mul8_ha_0_3_y1;
  wire h_s_arr_mul8_and_1_3_y0;
  wire h_s_arr_mul8_fa_1_3_y2;
  wire h_s_arr_mul8_fa_1_3_y4;
  wire h_s_arr_mul8_and_2_3_y0;
  wire h_s_arr_mul8_fa_2_3_y2;
  wire h_s_arr_mul8_fa_2_3_y4;
  wire h_s_arr_mul8_and_3_3_y0;
  wire h_s_arr_mul8_fa_3_3_y2;
  wire h_s_arr_mul8_fa_3_3_y4;
  wire h_s_arr_mul8_and_4_3_y0;
  wire h_s_arr_mul8_fa_4_3_y2;
  wire h_s_arr_mul8_fa_4_3_y4;
  wire h_s_arr_mul8_and_5_3_y0;
  wire h_s_arr_mul8_fa_5_3_y2;
  wire h_s_arr_mul8_fa_5_3_y4;
  wire h_s_arr_mul8_and_6_3_y0;
  wire h_s_arr_mul8_fa_6_3_y2;
  wire h_s_arr_mul8_fa_6_3_y4;
  wire h_s_arr_mul8_nand_7_3_y0;
  wire h_s_arr_mul8_fa_7_3_y2;
  wire h_s_arr_mul8_fa_7_3_y4;
  wire h_s_arr_mul8_and_0_4_y0;
  wire h_s_arr_mul8_ha_0_4_y0;
  wire h_s_arr_mul8_ha_0_4_y1;
  wire h_s_arr_mul8_and_1_4_y0;
  wire h_s_arr_mul8_fa_1_4_y2;
  wire h_s_arr_mul8_fa_1_4_y4;
  wire h_s_arr_mul8_and_2_4_y0;
  wire h_s_arr_mul8_fa_2_4_y2;
  wire h_s_arr_mul8_fa_2_4_y4;
  wire h_s_arr_mul8_and_3_4_y0;
  wire h_s_arr_mul8_fa_3_4_y2;
  wire h_s_arr_mul8_fa_3_4_y4;
  wire h_s_arr_mul8_and_4_4_y0;
  wire h_s_arr_mul8_fa_4_4_y2;
  wire h_s_arr_mul8_fa_4_4_y4;
  wire h_s_arr_mul8_and_5_4_y0;
  wire h_s_arr_mul8_fa_5_4_y2;
  wire h_s_arr_mul8_fa_5_4_y4;
  wire h_s_arr_mul8_and_6_4_y0;
  wire h_s_arr_mul8_fa_6_4_y2;
  wire h_s_arr_mul8_fa_6_4_y4;
  wire h_s_arr_mul8_nand_7_4_y0;
  wire h_s_arr_mul8_fa_7_4_y2;
  wire h_s_arr_mul8_fa_7_4_y4;
  wire h_s_arr_mul8_and_0_5_y0;
  wire h_s_arr_mul8_ha_0_5_y0;
  wire h_s_arr_mul8_ha_0_5_y1;
  wire h_s_arr_mul8_and_1_5_y0;
  wire h_s_arr_mul8_fa_1_5_y2;
  wire h_s_arr_mul8_fa_1_5_y4;
  wire h_s_arr_mul8_and_2_5_y0;
  wire h_s_arr_mul8_fa_2_5_y2;
  wire h_s_arr_mul8_fa_2_5_y4;
  wire h_s_arr_mul8_and_3_5_y0;
  wire h_s_arr_mul8_fa_3_5_y2;
  wire h_s_arr_mul8_fa_3_5_y4;
  wire h_s_arr_mul8_and_4_5_y0;
  wire h_s_arr_mul8_fa_4_5_y2;
  wire h_s_arr_mul8_fa_4_5_y4;
  wire h_s_arr_mul8_and_5_5_y0;
  wire h_s_arr_mul8_fa_5_5_y2;
  wire h_s_arr_mul8_fa_5_5_y4;
  wire h_s_arr_mul8_and_6_5_y0;
  wire h_s_arr_mul8_fa_6_5_y2;
  wire h_s_arr_mul8_fa_6_5_y4;
  wire h_s_arr_mul8_nand_7_5_y0;
  wire h_s_arr_mul8_fa_7_5_y2;
  wire h_s_arr_mul8_fa_7_5_y4;
  wire h_s_arr_mul8_and_0_6_y0;
  wire h_s_arr_mul8_ha_0_6_y0;
  wire h_s_arr_mul8_ha_0_6_y1;
  wire h_s_arr_mul8_and_1_6_y0;
  wire h_s_arr_mul8_fa_1_6_y2;
  wire h_s_arr_mul8_fa_1_6_y4;
  wire h_s_arr_mul8_and_2_6_y0;
  wire h_s_arr_mul8_fa_2_6_y2;
  wire h_s_arr_mul8_fa_2_6_y4;
  wire h_s_arr_mul8_and_3_6_y0;
  wire h_s_arr_mul8_fa_3_6_y2;
  wire h_s_arr_mul8_fa_3_6_y4;
  wire h_s_arr_mul8_and_4_6_y0;
  wire h_s_arr_mul8_fa_4_6_y2;
  wire h_s_arr_mul8_fa_4_6_y4;
  wire h_s_arr_mul8_and_5_6_y0;
  wire h_s_arr_mul8_fa_5_6_y2;
  wire h_s_arr_mul8_fa_5_6_y4;
  wire h_s_arr_mul8_and_6_6_y0;
  wire h_s_arr_mul8_fa_6_6_y2;
  wire h_s_arr_mul8_fa_6_6_y4;
  wire h_s_arr_mul8_nand_7_6_y0;
  wire h_s_arr_mul8_fa_7_6_y2;
  wire h_s_arr_mul8_fa_7_6_y4;
  wire h_s_arr_mul8_nand_0_7_y0;
  wire h_s_arr_mul8_ha_0_7_y0;
  wire h_s_arr_mul8_ha_0_7_y1;
  wire h_s_arr_mul8_nand_1_7_y0;
  wire h_s_arr_mul8_fa_1_7_y2;
  wire h_s_arr_mul8_fa_1_7_y4;
  wire h_s_arr_mul8_nand_2_7_y0;
  wire h_s_arr_mul8_fa_2_7_y2;
  wire h_s_arr_mul8_fa_2_7_y4;
  wire h_s_arr_mul8_nand_3_7_y0;
  wire h_s_arr_mul8_fa_3_7_y2;
  wire h_s_arr_mul8_fa_3_7_y4;
  wire h_s_arr_mul8_nand_4_7_y0;
  wire h_s_arr_mul8_fa_4_7_y2;
  wire h_s_arr_mul8_fa_4_7_y4;
  wire h_s_arr_mul8_nand_5_7_y0;
  wire h_s_arr_mul8_fa_5_7_y2;
  wire h_s_arr_mul8_fa_5_7_y4;
  wire h_s_arr_mul8_nand_6_7_y0;
  wire h_s_arr_mul8_fa_6_7_y2;
  wire h_s_arr_mul8_fa_6_7_y4;
  wire h_s_arr_mul8_and_7_7_y0;
  wire h_s_arr_mul8_fa_7_7_y2;
  wire h_s_arr_mul8_fa_7_7_y4;
  wire h_s_arr_mul8_xor_8_7_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  xor_gate xor_gate_h_s_arr_mul8_xor_constant_wire_y0(a_0, b_0, h_s_arr_mul8_xor_constant_wire_y0);
  xnor_gate xnor_gate_h_s_arr_mul8_xnor_constant_wire_y0(a_0, b_0, h_s_arr_mul8_xnor_constant_wire_y0);
  or_gate or_gate_constant_wire(h_s_arr_mul8_xor_constant_wire_y0, h_s_arr_mul8_xnor_constant_wire_y0, constant_wire);
  and_gate and_gate_h_s_arr_mul8_and_0_0_y0(a_0, b_0, h_s_arr_mul8_and_0_0_y0);
  and_gate and_gate_h_s_arr_mul8_and_1_0_y0(a_1, b_0, h_s_arr_mul8_and_1_0_y0);
  and_gate and_gate_h_s_arr_mul8_and_2_0_y0(a_2, b_0, h_s_arr_mul8_and_2_0_y0);
  and_gate and_gate_h_s_arr_mul8_and_3_0_y0(a_3, b_0, h_s_arr_mul8_and_3_0_y0);
  and_gate and_gate_h_s_arr_mul8_and_4_0_y0(a_4, b_0, h_s_arr_mul8_and_4_0_y0);
  and_gate and_gate_h_s_arr_mul8_and_5_0_y0(a_5, b_0, h_s_arr_mul8_and_5_0_y0);
  and_gate and_gate_h_s_arr_mul8_and_6_0_y0(a_6, b_0, h_s_arr_mul8_and_6_0_y0);
  nand_gate nand_gate_h_s_arr_mul8_nand_7_0_y0(a_7, b_0, h_s_arr_mul8_nand_7_0_y0);
  and_gate and_gate_h_s_arr_mul8_and_0_1_y0(a_0, b_1, h_s_arr_mul8_and_0_1_y0);
  ha ha_h_s_arr_mul8_ha_0_1_y1(h_s_arr_mul8_and_0_1_y0, h_s_arr_mul8_and_1_0_y0, h_s_arr_mul8_ha_0_1_y0, h_s_arr_mul8_ha_0_1_y1);
  and_gate and_gate_h_s_arr_mul8_and_1_1_y0(a_1, b_1, h_s_arr_mul8_and_1_1_y0);
  fa fa_h_s_arr_mul8_fa_1_1_y4(h_s_arr_mul8_and_1_1_y0, h_s_arr_mul8_and_2_0_y0, h_s_arr_mul8_ha_0_1_y1, h_s_arr_mul8_fa_1_1_y2, h_s_arr_mul8_fa_1_1_y4);
  and_gate and_gate_h_s_arr_mul8_and_2_1_y0(a_2, b_1, h_s_arr_mul8_and_2_1_y0);
  fa fa_h_s_arr_mul8_fa_2_1_y4(h_s_arr_mul8_and_2_1_y0, h_s_arr_mul8_and_3_0_y0, h_s_arr_mul8_fa_1_1_y4, h_s_arr_mul8_fa_2_1_y2, h_s_arr_mul8_fa_2_1_y4);
  and_gate and_gate_h_s_arr_mul8_and_3_1_y0(a_3, b_1, h_s_arr_mul8_and_3_1_y0);
  fa fa_h_s_arr_mul8_fa_3_1_y4(h_s_arr_mul8_and_3_1_y0, h_s_arr_mul8_and_4_0_y0, h_s_arr_mul8_fa_2_1_y4, h_s_arr_mul8_fa_3_1_y2, h_s_arr_mul8_fa_3_1_y4);
  and_gate and_gate_h_s_arr_mul8_and_4_1_y0(a_4, b_1, h_s_arr_mul8_and_4_1_y0);
  fa fa_h_s_arr_mul8_fa_4_1_y4(h_s_arr_mul8_and_4_1_y0, h_s_arr_mul8_and_5_0_y0, h_s_arr_mul8_fa_3_1_y4, h_s_arr_mul8_fa_4_1_y2, h_s_arr_mul8_fa_4_1_y4);
  and_gate and_gate_h_s_arr_mul8_and_5_1_y0(a_5, b_1, h_s_arr_mul8_and_5_1_y0);
  fa fa_h_s_arr_mul8_fa_5_1_y4(h_s_arr_mul8_and_5_1_y0, h_s_arr_mul8_and_6_0_y0, h_s_arr_mul8_fa_4_1_y4, h_s_arr_mul8_fa_5_1_y2, h_s_arr_mul8_fa_5_1_y4);
  and_gate and_gate_h_s_arr_mul8_and_6_1_y0(a_6, b_1, h_s_arr_mul8_and_6_1_y0);
  fa fa_h_s_arr_mul8_fa_6_1_y4(h_s_arr_mul8_and_6_1_y0, h_s_arr_mul8_nand_7_0_y0, h_s_arr_mul8_fa_5_1_y4, h_s_arr_mul8_fa_6_1_y2, h_s_arr_mul8_fa_6_1_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_7_1_y0(a_7, b_1, h_s_arr_mul8_nand_7_1_y0);
  fa fa_h_s_arr_mul8_fa_7_1_y4(h_s_arr_mul8_nand_7_1_y0, constant_wire, h_s_arr_mul8_fa_6_1_y4, h_s_arr_mul8_fa_7_1_y2, h_s_arr_mul8_fa_7_1_y4);
  and_gate and_gate_h_s_arr_mul8_and_0_2_y0(a_0, b_2, h_s_arr_mul8_and_0_2_y0);
  ha ha_h_s_arr_mul8_ha_0_2_y1(h_s_arr_mul8_and_0_2_y0, h_s_arr_mul8_fa_1_1_y2, h_s_arr_mul8_ha_0_2_y0, h_s_arr_mul8_ha_0_2_y1);
  and_gate and_gate_h_s_arr_mul8_and_1_2_y0(a_1, b_2, h_s_arr_mul8_and_1_2_y0);
  fa fa_h_s_arr_mul8_fa_1_2_y4(h_s_arr_mul8_and_1_2_y0, h_s_arr_mul8_fa_2_1_y2, h_s_arr_mul8_ha_0_2_y1, h_s_arr_mul8_fa_1_2_y2, h_s_arr_mul8_fa_1_2_y4);
  and_gate and_gate_h_s_arr_mul8_and_2_2_y0(a_2, b_2, h_s_arr_mul8_and_2_2_y0);
  fa fa_h_s_arr_mul8_fa_2_2_y4(h_s_arr_mul8_and_2_2_y0, h_s_arr_mul8_fa_3_1_y2, h_s_arr_mul8_fa_1_2_y4, h_s_arr_mul8_fa_2_2_y2, h_s_arr_mul8_fa_2_2_y4);
  and_gate and_gate_h_s_arr_mul8_and_3_2_y0(a_3, b_2, h_s_arr_mul8_and_3_2_y0);
  fa fa_h_s_arr_mul8_fa_3_2_y4(h_s_arr_mul8_and_3_2_y0, h_s_arr_mul8_fa_4_1_y2, h_s_arr_mul8_fa_2_2_y4, h_s_arr_mul8_fa_3_2_y2, h_s_arr_mul8_fa_3_2_y4);
  and_gate and_gate_h_s_arr_mul8_and_4_2_y0(a_4, b_2, h_s_arr_mul8_and_4_2_y0);
  fa fa_h_s_arr_mul8_fa_4_2_y4(h_s_arr_mul8_and_4_2_y0, h_s_arr_mul8_fa_5_1_y2, h_s_arr_mul8_fa_3_2_y4, h_s_arr_mul8_fa_4_2_y2, h_s_arr_mul8_fa_4_2_y4);
  and_gate and_gate_h_s_arr_mul8_and_5_2_y0(a_5, b_2, h_s_arr_mul8_and_5_2_y0);
  fa fa_h_s_arr_mul8_fa_5_2_y4(h_s_arr_mul8_and_5_2_y0, h_s_arr_mul8_fa_6_1_y2, h_s_arr_mul8_fa_4_2_y4, h_s_arr_mul8_fa_5_2_y2, h_s_arr_mul8_fa_5_2_y4);
  and_gate and_gate_h_s_arr_mul8_and_6_2_y0(a_6, b_2, h_s_arr_mul8_and_6_2_y0);
  fa fa_h_s_arr_mul8_fa_6_2_y4(h_s_arr_mul8_and_6_2_y0, h_s_arr_mul8_fa_7_1_y2, h_s_arr_mul8_fa_5_2_y4, h_s_arr_mul8_fa_6_2_y2, h_s_arr_mul8_fa_6_2_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_7_2_y0(a_7, b_2, h_s_arr_mul8_nand_7_2_y0);
  fa fa_h_s_arr_mul8_fa_7_2_y4(h_s_arr_mul8_nand_7_2_y0, h_s_arr_mul8_fa_7_1_y4, h_s_arr_mul8_fa_6_2_y4, h_s_arr_mul8_fa_7_2_y2, h_s_arr_mul8_fa_7_2_y4);
  and_gate and_gate_h_s_arr_mul8_and_0_3_y0(a_0, b_3, h_s_arr_mul8_and_0_3_y0);
  ha ha_h_s_arr_mul8_ha_0_3_y1(h_s_arr_mul8_and_0_3_y0, h_s_arr_mul8_fa_1_2_y2, h_s_arr_mul8_ha_0_3_y0, h_s_arr_mul8_ha_0_3_y1);
  and_gate and_gate_h_s_arr_mul8_and_1_3_y0(a_1, b_3, h_s_arr_mul8_and_1_3_y0);
  fa fa_h_s_arr_mul8_fa_1_3_y4(h_s_arr_mul8_and_1_3_y0, h_s_arr_mul8_fa_2_2_y2, h_s_arr_mul8_ha_0_3_y1, h_s_arr_mul8_fa_1_3_y2, h_s_arr_mul8_fa_1_3_y4);
  and_gate and_gate_h_s_arr_mul8_and_2_3_y0(a_2, b_3, h_s_arr_mul8_and_2_3_y0);
  fa fa_h_s_arr_mul8_fa_2_3_y4(h_s_arr_mul8_and_2_3_y0, h_s_arr_mul8_fa_3_2_y2, h_s_arr_mul8_fa_1_3_y4, h_s_arr_mul8_fa_2_3_y2, h_s_arr_mul8_fa_2_3_y4);
  and_gate and_gate_h_s_arr_mul8_and_3_3_y0(a_3, b_3, h_s_arr_mul8_and_3_3_y0);
  fa fa_h_s_arr_mul8_fa_3_3_y4(h_s_arr_mul8_and_3_3_y0, h_s_arr_mul8_fa_4_2_y2, h_s_arr_mul8_fa_2_3_y4, h_s_arr_mul8_fa_3_3_y2, h_s_arr_mul8_fa_3_3_y4);
  and_gate and_gate_h_s_arr_mul8_and_4_3_y0(a_4, b_3, h_s_arr_mul8_and_4_3_y0);
  fa fa_h_s_arr_mul8_fa_4_3_y4(h_s_arr_mul8_and_4_3_y0, h_s_arr_mul8_fa_5_2_y2, h_s_arr_mul8_fa_3_3_y4, h_s_arr_mul8_fa_4_3_y2, h_s_arr_mul8_fa_4_3_y4);
  and_gate and_gate_h_s_arr_mul8_and_5_3_y0(a_5, b_3, h_s_arr_mul8_and_5_3_y0);
  fa fa_h_s_arr_mul8_fa_5_3_y4(h_s_arr_mul8_and_5_3_y0, h_s_arr_mul8_fa_6_2_y2, h_s_arr_mul8_fa_4_3_y4, h_s_arr_mul8_fa_5_3_y2, h_s_arr_mul8_fa_5_3_y4);
  and_gate and_gate_h_s_arr_mul8_and_6_3_y0(a_6, b_3, h_s_arr_mul8_and_6_3_y0);
  fa fa_h_s_arr_mul8_fa_6_3_y4(h_s_arr_mul8_and_6_3_y0, h_s_arr_mul8_fa_7_2_y2, h_s_arr_mul8_fa_5_3_y4, h_s_arr_mul8_fa_6_3_y2, h_s_arr_mul8_fa_6_3_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_7_3_y0(a_7, b_3, h_s_arr_mul8_nand_7_3_y0);
  fa fa_h_s_arr_mul8_fa_7_3_y4(h_s_arr_mul8_nand_7_3_y0, h_s_arr_mul8_fa_7_2_y4, h_s_arr_mul8_fa_6_3_y4, h_s_arr_mul8_fa_7_3_y2, h_s_arr_mul8_fa_7_3_y4);
  and_gate and_gate_h_s_arr_mul8_and_0_4_y0(a_0, b_4, h_s_arr_mul8_and_0_4_y0);
  ha ha_h_s_arr_mul8_ha_0_4_y1(h_s_arr_mul8_and_0_4_y0, h_s_arr_mul8_fa_1_3_y2, h_s_arr_mul8_ha_0_4_y0, h_s_arr_mul8_ha_0_4_y1);
  and_gate and_gate_h_s_arr_mul8_and_1_4_y0(a_1, b_4, h_s_arr_mul8_and_1_4_y0);
  fa fa_h_s_arr_mul8_fa_1_4_y4(h_s_arr_mul8_and_1_4_y0, h_s_arr_mul8_fa_2_3_y2, h_s_arr_mul8_ha_0_4_y1, h_s_arr_mul8_fa_1_4_y2, h_s_arr_mul8_fa_1_4_y4);
  and_gate and_gate_h_s_arr_mul8_and_2_4_y0(a_2, b_4, h_s_arr_mul8_and_2_4_y0);
  fa fa_h_s_arr_mul8_fa_2_4_y4(h_s_arr_mul8_and_2_4_y0, h_s_arr_mul8_fa_3_3_y2, h_s_arr_mul8_fa_1_4_y4, h_s_arr_mul8_fa_2_4_y2, h_s_arr_mul8_fa_2_4_y4);
  and_gate and_gate_h_s_arr_mul8_and_3_4_y0(a_3, b_4, h_s_arr_mul8_and_3_4_y0);
  fa fa_h_s_arr_mul8_fa_3_4_y4(h_s_arr_mul8_and_3_4_y0, h_s_arr_mul8_fa_4_3_y2, h_s_arr_mul8_fa_2_4_y4, h_s_arr_mul8_fa_3_4_y2, h_s_arr_mul8_fa_3_4_y4);
  and_gate and_gate_h_s_arr_mul8_and_4_4_y0(a_4, b_4, h_s_arr_mul8_and_4_4_y0);
  fa fa_h_s_arr_mul8_fa_4_4_y4(h_s_arr_mul8_and_4_4_y0, h_s_arr_mul8_fa_5_3_y2, h_s_arr_mul8_fa_3_4_y4, h_s_arr_mul8_fa_4_4_y2, h_s_arr_mul8_fa_4_4_y4);
  and_gate and_gate_h_s_arr_mul8_and_5_4_y0(a_5, b_4, h_s_arr_mul8_and_5_4_y0);
  fa fa_h_s_arr_mul8_fa_5_4_y4(h_s_arr_mul8_and_5_4_y0, h_s_arr_mul8_fa_6_3_y2, h_s_arr_mul8_fa_4_4_y4, h_s_arr_mul8_fa_5_4_y2, h_s_arr_mul8_fa_5_4_y4);
  and_gate and_gate_h_s_arr_mul8_and_6_4_y0(a_6, b_4, h_s_arr_mul8_and_6_4_y0);
  fa fa_h_s_arr_mul8_fa_6_4_y4(h_s_arr_mul8_and_6_4_y0, h_s_arr_mul8_fa_7_3_y2, h_s_arr_mul8_fa_5_4_y4, h_s_arr_mul8_fa_6_4_y2, h_s_arr_mul8_fa_6_4_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_7_4_y0(a_7, b_4, h_s_arr_mul8_nand_7_4_y0);
  fa fa_h_s_arr_mul8_fa_7_4_y4(h_s_arr_mul8_nand_7_4_y0, h_s_arr_mul8_fa_7_3_y4, h_s_arr_mul8_fa_6_4_y4, h_s_arr_mul8_fa_7_4_y2, h_s_arr_mul8_fa_7_4_y4);
  and_gate and_gate_h_s_arr_mul8_and_0_5_y0(a_0, b_5, h_s_arr_mul8_and_0_5_y0);
  ha ha_h_s_arr_mul8_ha_0_5_y1(h_s_arr_mul8_and_0_5_y0, h_s_arr_mul8_fa_1_4_y2, h_s_arr_mul8_ha_0_5_y0, h_s_arr_mul8_ha_0_5_y1);
  and_gate and_gate_h_s_arr_mul8_and_1_5_y0(a_1, b_5, h_s_arr_mul8_and_1_5_y0);
  fa fa_h_s_arr_mul8_fa_1_5_y4(h_s_arr_mul8_and_1_5_y0, h_s_arr_mul8_fa_2_4_y2, h_s_arr_mul8_ha_0_5_y1, h_s_arr_mul8_fa_1_5_y2, h_s_arr_mul8_fa_1_5_y4);
  and_gate and_gate_h_s_arr_mul8_and_2_5_y0(a_2, b_5, h_s_arr_mul8_and_2_5_y0);
  fa fa_h_s_arr_mul8_fa_2_5_y4(h_s_arr_mul8_and_2_5_y0, h_s_arr_mul8_fa_3_4_y2, h_s_arr_mul8_fa_1_5_y4, h_s_arr_mul8_fa_2_5_y2, h_s_arr_mul8_fa_2_5_y4);
  and_gate and_gate_h_s_arr_mul8_and_3_5_y0(a_3, b_5, h_s_arr_mul8_and_3_5_y0);
  fa fa_h_s_arr_mul8_fa_3_5_y4(h_s_arr_mul8_and_3_5_y0, h_s_arr_mul8_fa_4_4_y2, h_s_arr_mul8_fa_2_5_y4, h_s_arr_mul8_fa_3_5_y2, h_s_arr_mul8_fa_3_5_y4);
  and_gate and_gate_h_s_arr_mul8_and_4_5_y0(a_4, b_5, h_s_arr_mul8_and_4_5_y0);
  fa fa_h_s_arr_mul8_fa_4_5_y4(h_s_arr_mul8_and_4_5_y0, h_s_arr_mul8_fa_5_4_y2, h_s_arr_mul8_fa_3_5_y4, h_s_arr_mul8_fa_4_5_y2, h_s_arr_mul8_fa_4_5_y4);
  and_gate and_gate_h_s_arr_mul8_and_5_5_y0(a_5, b_5, h_s_arr_mul8_and_5_5_y0);
  fa fa_h_s_arr_mul8_fa_5_5_y4(h_s_arr_mul8_and_5_5_y0, h_s_arr_mul8_fa_6_4_y2, h_s_arr_mul8_fa_4_5_y4, h_s_arr_mul8_fa_5_5_y2, h_s_arr_mul8_fa_5_5_y4);
  and_gate and_gate_h_s_arr_mul8_and_6_5_y0(a_6, b_5, h_s_arr_mul8_and_6_5_y0);
  fa fa_h_s_arr_mul8_fa_6_5_y4(h_s_arr_mul8_and_6_5_y0, h_s_arr_mul8_fa_7_4_y2, h_s_arr_mul8_fa_5_5_y4, h_s_arr_mul8_fa_6_5_y2, h_s_arr_mul8_fa_6_5_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_7_5_y0(a_7, b_5, h_s_arr_mul8_nand_7_5_y0);
  fa fa_h_s_arr_mul8_fa_7_5_y4(h_s_arr_mul8_nand_7_5_y0, h_s_arr_mul8_fa_7_4_y4, h_s_arr_mul8_fa_6_5_y4, h_s_arr_mul8_fa_7_5_y2, h_s_arr_mul8_fa_7_5_y4);
  and_gate and_gate_h_s_arr_mul8_and_0_6_y0(a_0, b_6, h_s_arr_mul8_and_0_6_y0);
  ha ha_h_s_arr_mul8_ha_0_6_y1(h_s_arr_mul8_and_0_6_y0, h_s_arr_mul8_fa_1_5_y2, h_s_arr_mul8_ha_0_6_y0, h_s_arr_mul8_ha_0_6_y1);
  and_gate and_gate_h_s_arr_mul8_and_1_6_y0(a_1, b_6, h_s_arr_mul8_and_1_6_y0);
  fa fa_h_s_arr_mul8_fa_1_6_y4(h_s_arr_mul8_and_1_6_y0, h_s_arr_mul8_fa_2_5_y2, h_s_arr_mul8_ha_0_6_y1, h_s_arr_mul8_fa_1_6_y2, h_s_arr_mul8_fa_1_6_y4);
  and_gate and_gate_h_s_arr_mul8_and_2_6_y0(a_2, b_6, h_s_arr_mul8_and_2_6_y0);
  fa fa_h_s_arr_mul8_fa_2_6_y4(h_s_arr_mul8_and_2_6_y0, h_s_arr_mul8_fa_3_5_y2, h_s_arr_mul8_fa_1_6_y4, h_s_arr_mul8_fa_2_6_y2, h_s_arr_mul8_fa_2_6_y4);
  and_gate and_gate_h_s_arr_mul8_and_3_6_y0(a_3, b_6, h_s_arr_mul8_and_3_6_y0);
  fa fa_h_s_arr_mul8_fa_3_6_y4(h_s_arr_mul8_and_3_6_y0, h_s_arr_mul8_fa_4_5_y2, h_s_arr_mul8_fa_2_6_y4, h_s_arr_mul8_fa_3_6_y2, h_s_arr_mul8_fa_3_6_y4);
  and_gate and_gate_h_s_arr_mul8_and_4_6_y0(a_4, b_6, h_s_arr_mul8_and_4_6_y0);
  fa fa_h_s_arr_mul8_fa_4_6_y4(h_s_arr_mul8_and_4_6_y0, h_s_arr_mul8_fa_5_5_y2, h_s_arr_mul8_fa_3_6_y4, h_s_arr_mul8_fa_4_6_y2, h_s_arr_mul8_fa_4_6_y4);
  and_gate and_gate_h_s_arr_mul8_and_5_6_y0(a_5, b_6, h_s_arr_mul8_and_5_6_y0);
  fa fa_h_s_arr_mul8_fa_5_6_y4(h_s_arr_mul8_and_5_6_y0, h_s_arr_mul8_fa_6_5_y2, h_s_arr_mul8_fa_4_6_y4, h_s_arr_mul8_fa_5_6_y2, h_s_arr_mul8_fa_5_6_y4);
  and_gate and_gate_h_s_arr_mul8_and_6_6_y0(a_6, b_6, h_s_arr_mul8_and_6_6_y0);
  fa fa_h_s_arr_mul8_fa_6_6_y4(h_s_arr_mul8_and_6_6_y0, h_s_arr_mul8_fa_7_5_y2, h_s_arr_mul8_fa_5_6_y4, h_s_arr_mul8_fa_6_6_y2, h_s_arr_mul8_fa_6_6_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_7_6_y0(a_7, b_6, h_s_arr_mul8_nand_7_6_y0);
  fa fa_h_s_arr_mul8_fa_7_6_y4(h_s_arr_mul8_nand_7_6_y0, h_s_arr_mul8_fa_7_5_y4, h_s_arr_mul8_fa_6_6_y4, h_s_arr_mul8_fa_7_6_y2, h_s_arr_mul8_fa_7_6_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_0_7_y0(a_0, b_7, h_s_arr_mul8_nand_0_7_y0);
  ha ha_h_s_arr_mul8_ha_0_7_y1(h_s_arr_mul8_nand_0_7_y0, h_s_arr_mul8_fa_1_6_y2, h_s_arr_mul8_ha_0_7_y0, h_s_arr_mul8_ha_0_7_y1);
  nand_gate nand_gate_h_s_arr_mul8_nand_1_7_y0(a_1, b_7, h_s_arr_mul8_nand_1_7_y0);
  fa fa_h_s_arr_mul8_fa_1_7_y4(h_s_arr_mul8_nand_1_7_y0, h_s_arr_mul8_fa_2_6_y2, h_s_arr_mul8_ha_0_7_y1, h_s_arr_mul8_fa_1_7_y2, h_s_arr_mul8_fa_1_7_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_2_7_y0(a_2, b_7, h_s_arr_mul8_nand_2_7_y0);
  fa fa_h_s_arr_mul8_fa_2_7_y4(h_s_arr_mul8_nand_2_7_y0, h_s_arr_mul8_fa_3_6_y2, h_s_arr_mul8_fa_1_7_y4, h_s_arr_mul8_fa_2_7_y2, h_s_arr_mul8_fa_2_7_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_3_7_y0(a_3, b_7, h_s_arr_mul8_nand_3_7_y0);
  fa fa_h_s_arr_mul8_fa_3_7_y4(h_s_arr_mul8_nand_3_7_y0, h_s_arr_mul8_fa_4_6_y2, h_s_arr_mul8_fa_2_7_y4, h_s_arr_mul8_fa_3_7_y2, h_s_arr_mul8_fa_3_7_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_4_7_y0(a_4, b_7, h_s_arr_mul8_nand_4_7_y0);
  fa fa_h_s_arr_mul8_fa_4_7_y4(h_s_arr_mul8_nand_4_7_y0, h_s_arr_mul8_fa_5_6_y2, h_s_arr_mul8_fa_3_7_y4, h_s_arr_mul8_fa_4_7_y2, h_s_arr_mul8_fa_4_7_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_5_7_y0(a_5, b_7, h_s_arr_mul8_nand_5_7_y0);
  fa fa_h_s_arr_mul8_fa_5_7_y4(h_s_arr_mul8_nand_5_7_y0, h_s_arr_mul8_fa_6_6_y2, h_s_arr_mul8_fa_4_7_y4, h_s_arr_mul8_fa_5_7_y2, h_s_arr_mul8_fa_5_7_y4);
  nand_gate nand_gate_h_s_arr_mul8_nand_6_7_y0(a_6, b_7, h_s_arr_mul8_nand_6_7_y0);
  fa fa_h_s_arr_mul8_fa_6_7_y4(h_s_arr_mul8_nand_6_7_y0, h_s_arr_mul8_fa_7_6_y2, h_s_arr_mul8_fa_5_7_y4, h_s_arr_mul8_fa_6_7_y2, h_s_arr_mul8_fa_6_7_y4);
  and_gate and_gate_h_s_arr_mul8_and_7_7_y0(a_7, b_7, h_s_arr_mul8_and_7_7_y0);
  fa fa_h_s_arr_mul8_fa_7_7_y4(h_s_arr_mul8_and_7_7_y0, h_s_arr_mul8_fa_7_6_y4, h_s_arr_mul8_fa_6_7_y4, h_s_arr_mul8_fa_7_7_y2, h_s_arr_mul8_fa_7_7_y4);
  xor_gate xor_gate_h_s_arr_mul8_xor_8_7_y0(h_s_arr_mul8_fa_7_7_y4, constant_wire, h_s_arr_mul8_xor_8_7_y0);

  assign out[0] = h_s_arr_mul8_and_0_0_y0;
  assign out[1] = h_s_arr_mul8_ha_0_1_y0;
  assign out[2] = h_s_arr_mul8_ha_0_2_y0;
  assign out[3] = h_s_arr_mul8_ha_0_3_y0;
  assign out[4] = h_s_arr_mul8_ha_0_4_y0;
  assign out[5] = h_s_arr_mul8_ha_0_5_y0;
  assign out[6] = h_s_arr_mul8_ha_0_6_y0;
  assign out[7] = h_s_arr_mul8_ha_0_7_y0;
  assign out[8] = h_s_arr_mul8_fa_1_7_y2;
  assign out[9] = h_s_arr_mul8_fa_2_7_y2;
  assign out[10] = h_s_arr_mul8_fa_3_7_y2;
  assign out[11] = h_s_arr_mul8_fa_4_7_y2;
  assign out[12] = h_s_arr_mul8_fa_5_7_y2;
  assign out[13] = h_s_arr_mul8_fa_6_7_y2;
  assign out[14] = h_s_arr_mul8_fa_7_7_y2;
  assign out[15] = h_s_arr_mul8_xor_8_7_y0;
endmodule