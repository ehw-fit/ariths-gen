module f_s_cska32(input [31:0] a, input [31:0] b, output [32:0] f_s_cska32_out);
  wire f_s_cska32_xor0;
  wire f_s_cska32_ha0_xor0;
  wire f_s_cska32_ha0_and0;
  wire f_s_cska32_xor1;
  wire f_s_cska32_fa0_xor0;
  wire f_s_cska32_fa0_and0;
  wire f_s_cska32_fa0_xor1;
  wire f_s_cska32_fa0_and1;
  wire f_s_cska32_fa0_or0;
  wire f_s_cska32_xor2;
  wire f_s_cska32_fa1_xor0;
  wire f_s_cska32_fa1_and0;
  wire f_s_cska32_fa1_xor1;
  wire f_s_cska32_fa1_and1;
  wire f_s_cska32_fa1_or0;
  wire f_s_cska32_xor3;
  wire f_s_cska32_fa2_xor0;
  wire f_s_cska32_fa2_and0;
  wire f_s_cska32_fa2_xor1;
  wire f_s_cska32_fa2_and1;
  wire f_s_cska32_fa2_or0;
  wire f_s_cska32_and_propagate00;
  wire f_s_cska32_and_propagate01;
  wire f_s_cska32_and_propagate02;
  wire f_s_cska32_mux2to10_not0;
  wire f_s_cska32_mux2to10_and1;
  wire f_s_cska32_xor4;
  wire f_s_cska32_fa3_xor0;
  wire f_s_cska32_fa3_and0;
  wire f_s_cska32_fa3_xor1;
  wire f_s_cska32_fa3_and1;
  wire f_s_cska32_fa3_or0;
  wire f_s_cska32_xor5;
  wire f_s_cska32_fa4_xor0;
  wire f_s_cska32_fa4_and0;
  wire f_s_cska32_fa4_xor1;
  wire f_s_cska32_fa4_and1;
  wire f_s_cska32_fa4_or0;
  wire f_s_cska32_xor6;
  wire f_s_cska32_fa5_xor0;
  wire f_s_cska32_fa5_and0;
  wire f_s_cska32_fa5_xor1;
  wire f_s_cska32_fa5_and1;
  wire f_s_cska32_fa5_or0;
  wire f_s_cska32_xor7;
  wire f_s_cska32_fa6_xor0;
  wire f_s_cska32_fa6_and0;
  wire f_s_cska32_fa6_xor1;
  wire f_s_cska32_fa6_and1;
  wire f_s_cska32_fa6_or0;
  wire f_s_cska32_and_propagate13;
  wire f_s_cska32_and_propagate14;
  wire f_s_cska32_and_propagate15;
  wire f_s_cska32_mux2to11_and0;
  wire f_s_cska32_mux2to11_not0;
  wire f_s_cska32_mux2to11_and1;
  wire f_s_cska32_mux2to11_xor0;
  wire f_s_cska32_xor8;
  wire f_s_cska32_fa7_xor0;
  wire f_s_cska32_fa7_and0;
  wire f_s_cska32_fa7_xor1;
  wire f_s_cska32_fa7_and1;
  wire f_s_cska32_fa7_or0;
  wire f_s_cska32_xor9;
  wire f_s_cska32_fa8_xor0;
  wire f_s_cska32_fa8_and0;
  wire f_s_cska32_fa8_xor1;
  wire f_s_cska32_fa8_and1;
  wire f_s_cska32_fa8_or0;
  wire f_s_cska32_xor10;
  wire f_s_cska32_fa9_xor0;
  wire f_s_cska32_fa9_and0;
  wire f_s_cska32_fa9_xor1;
  wire f_s_cska32_fa9_and1;
  wire f_s_cska32_fa9_or0;
  wire f_s_cska32_xor11;
  wire f_s_cska32_fa10_xor0;
  wire f_s_cska32_fa10_and0;
  wire f_s_cska32_fa10_xor1;
  wire f_s_cska32_fa10_and1;
  wire f_s_cska32_fa10_or0;
  wire f_s_cska32_and_propagate26;
  wire f_s_cska32_and_propagate27;
  wire f_s_cska32_and_propagate28;
  wire f_s_cska32_mux2to12_and0;
  wire f_s_cska32_mux2to12_not0;
  wire f_s_cska32_mux2to12_and1;
  wire f_s_cska32_mux2to12_xor0;
  wire f_s_cska32_xor12;
  wire f_s_cska32_fa11_xor0;
  wire f_s_cska32_fa11_and0;
  wire f_s_cska32_fa11_xor1;
  wire f_s_cska32_fa11_and1;
  wire f_s_cska32_fa11_or0;
  wire f_s_cska32_xor13;
  wire f_s_cska32_fa12_xor0;
  wire f_s_cska32_fa12_and0;
  wire f_s_cska32_fa12_xor1;
  wire f_s_cska32_fa12_and1;
  wire f_s_cska32_fa12_or0;
  wire f_s_cska32_xor14;
  wire f_s_cska32_fa13_xor0;
  wire f_s_cska32_fa13_and0;
  wire f_s_cska32_fa13_xor1;
  wire f_s_cska32_fa13_and1;
  wire f_s_cska32_fa13_or0;
  wire f_s_cska32_xor15;
  wire f_s_cska32_fa14_xor0;
  wire f_s_cska32_fa14_and0;
  wire f_s_cska32_fa14_xor1;
  wire f_s_cska32_fa14_and1;
  wire f_s_cska32_fa14_or0;
  wire f_s_cska32_and_propagate39;
  wire f_s_cska32_and_propagate310;
  wire f_s_cska32_and_propagate311;
  wire f_s_cska32_mux2to13_and0;
  wire f_s_cska32_mux2to13_not0;
  wire f_s_cska32_mux2to13_and1;
  wire f_s_cska32_mux2to13_xor0;
  wire f_s_cska32_xor16;
  wire f_s_cska32_fa15_xor0;
  wire f_s_cska32_fa15_and0;
  wire f_s_cska32_fa15_xor1;
  wire f_s_cska32_fa15_and1;
  wire f_s_cska32_fa15_or0;
  wire f_s_cska32_xor17;
  wire f_s_cska32_fa16_xor0;
  wire f_s_cska32_fa16_and0;
  wire f_s_cska32_fa16_xor1;
  wire f_s_cska32_fa16_and1;
  wire f_s_cska32_fa16_or0;
  wire f_s_cska32_xor18;
  wire f_s_cska32_fa17_xor0;
  wire f_s_cska32_fa17_and0;
  wire f_s_cska32_fa17_xor1;
  wire f_s_cska32_fa17_and1;
  wire f_s_cska32_fa17_or0;
  wire f_s_cska32_xor19;
  wire f_s_cska32_fa18_xor0;
  wire f_s_cska32_fa18_and0;
  wire f_s_cska32_fa18_xor1;
  wire f_s_cska32_fa18_and1;
  wire f_s_cska32_fa18_or0;
  wire f_s_cska32_and_propagate412;
  wire f_s_cska32_and_propagate413;
  wire f_s_cska32_and_propagate414;
  wire f_s_cska32_mux2to14_and0;
  wire f_s_cska32_mux2to14_not0;
  wire f_s_cska32_mux2to14_and1;
  wire f_s_cska32_mux2to14_xor0;
  wire f_s_cska32_xor20;
  wire f_s_cska32_fa19_xor0;
  wire f_s_cska32_fa19_and0;
  wire f_s_cska32_fa19_xor1;
  wire f_s_cska32_fa19_and1;
  wire f_s_cska32_fa19_or0;
  wire f_s_cska32_xor21;
  wire f_s_cska32_fa20_xor0;
  wire f_s_cska32_fa20_and0;
  wire f_s_cska32_fa20_xor1;
  wire f_s_cska32_fa20_and1;
  wire f_s_cska32_fa20_or0;
  wire f_s_cska32_xor22;
  wire f_s_cska32_fa21_xor0;
  wire f_s_cska32_fa21_and0;
  wire f_s_cska32_fa21_xor1;
  wire f_s_cska32_fa21_and1;
  wire f_s_cska32_fa21_or0;
  wire f_s_cska32_xor23;
  wire f_s_cska32_fa22_xor0;
  wire f_s_cska32_fa22_and0;
  wire f_s_cska32_fa22_xor1;
  wire f_s_cska32_fa22_and1;
  wire f_s_cska32_fa22_or0;
  wire f_s_cska32_and_propagate515;
  wire f_s_cska32_and_propagate516;
  wire f_s_cska32_and_propagate517;
  wire f_s_cska32_mux2to15_and0;
  wire f_s_cska32_mux2to15_not0;
  wire f_s_cska32_mux2to15_and1;
  wire f_s_cska32_mux2to15_xor0;
  wire f_s_cska32_xor24;
  wire f_s_cska32_fa23_xor0;
  wire f_s_cska32_fa23_and0;
  wire f_s_cska32_fa23_xor1;
  wire f_s_cska32_fa23_and1;
  wire f_s_cska32_fa23_or0;
  wire f_s_cska32_xor25;
  wire f_s_cska32_fa24_xor0;
  wire f_s_cska32_fa24_and0;
  wire f_s_cska32_fa24_xor1;
  wire f_s_cska32_fa24_and1;
  wire f_s_cska32_fa24_or0;
  wire f_s_cska32_xor26;
  wire f_s_cska32_fa25_xor0;
  wire f_s_cska32_fa25_and0;
  wire f_s_cska32_fa25_xor1;
  wire f_s_cska32_fa25_and1;
  wire f_s_cska32_fa25_or0;
  wire f_s_cska32_xor27;
  wire f_s_cska32_fa26_xor0;
  wire f_s_cska32_fa26_and0;
  wire f_s_cska32_fa26_xor1;
  wire f_s_cska32_fa26_and1;
  wire f_s_cska32_fa26_or0;
  wire f_s_cska32_and_propagate618;
  wire f_s_cska32_and_propagate619;
  wire f_s_cska32_and_propagate620;
  wire f_s_cska32_mux2to16_and0;
  wire f_s_cska32_mux2to16_not0;
  wire f_s_cska32_mux2to16_and1;
  wire f_s_cska32_mux2to16_xor0;
  wire f_s_cska32_xor28;
  wire f_s_cska32_fa27_xor0;
  wire f_s_cska32_fa27_and0;
  wire f_s_cska32_fa27_xor1;
  wire f_s_cska32_fa27_and1;
  wire f_s_cska32_fa27_or0;
  wire f_s_cska32_xor29;
  wire f_s_cska32_fa28_xor0;
  wire f_s_cska32_fa28_and0;
  wire f_s_cska32_fa28_xor1;
  wire f_s_cska32_fa28_and1;
  wire f_s_cska32_fa28_or0;
  wire f_s_cska32_xor30;
  wire f_s_cska32_fa29_xor0;
  wire f_s_cska32_fa29_and0;
  wire f_s_cska32_fa29_xor1;
  wire f_s_cska32_fa29_and1;
  wire f_s_cska32_fa29_or0;
  wire f_s_cska32_xor31;
  wire f_s_cska32_fa30_xor0;
  wire f_s_cska32_fa30_and0;
  wire f_s_cska32_fa30_xor1;
  wire f_s_cska32_fa30_and1;
  wire f_s_cska32_fa30_or0;
  wire f_s_cska32_and_propagate721;
  wire f_s_cska32_and_propagate722;
  wire f_s_cska32_and_propagate723;
  wire f_s_cska32_mux2to17_and0;
  wire f_s_cska32_mux2to17_not0;
  wire f_s_cska32_mux2to17_and1;
  wire f_s_cska32_mux2to17_xor0;
  wire f_s_cska32_xor32;
  wire f_s_cska32_xor33;

  assign f_s_cska32_xor0 = a[0] ^ b[0];
  assign f_s_cska32_ha0_xor0 = a[0] ^ b[0];
  assign f_s_cska32_ha0_and0 = a[0] & b[0];
  assign f_s_cska32_xor1 = a[1] ^ b[1];
  assign f_s_cska32_fa0_xor0 = a[1] ^ b[1];
  assign f_s_cska32_fa0_and0 = a[1] & b[1];
  assign f_s_cska32_fa0_xor1 = f_s_cska32_fa0_xor0 ^ f_s_cska32_ha0_and0;
  assign f_s_cska32_fa0_and1 = f_s_cska32_fa0_xor0 & f_s_cska32_ha0_and0;
  assign f_s_cska32_fa0_or0 = f_s_cska32_fa0_and0 | f_s_cska32_fa0_and1;
  assign f_s_cska32_xor2 = a[2] ^ b[2];
  assign f_s_cska32_fa1_xor0 = a[2] ^ b[2];
  assign f_s_cska32_fa1_and0 = a[2] & b[2];
  assign f_s_cska32_fa1_xor1 = f_s_cska32_fa1_xor0 ^ f_s_cska32_fa0_or0;
  assign f_s_cska32_fa1_and1 = f_s_cska32_fa1_xor0 & f_s_cska32_fa0_or0;
  assign f_s_cska32_fa1_or0 = f_s_cska32_fa1_and0 | f_s_cska32_fa1_and1;
  assign f_s_cska32_xor3 = a[3] ^ b[3];
  assign f_s_cska32_fa2_xor0 = a[3] ^ b[3];
  assign f_s_cska32_fa2_and0 = a[3] & b[3];
  assign f_s_cska32_fa2_xor1 = f_s_cska32_fa2_xor0 ^ f_s_cska32_fa1_or0;
  assign f_s_cska32_fa2_and1 = f_s_cska32_fa2_xor0 & f_s_cska32_fa1_or0;
  assign f_s_cska32_fa2_or0 = f_s_cska32_fa2_and0 | f_s_cska32_fa2_and1;
  assign f_s_cska32_and_propagate00 = f_s_cska32_xor0 & f_s_cska32_xor2;
  assign f_s_cska32_and_propagate01 = f_s_cska32_xor1 & f_s_cska32_xor3;
  assign f_s_cska32_and_propagate02 = f_s_cska32_and_propagate00 & f_s_cska32_and_propagate01;
  assign f_s_cska32_mux2to10_not0 = ~f_s_cska32_and_propagate02;
  assign f_s_cska32_mux2to10_and1 = f_s_cska32_fa2_or0 & f_s_cska32_mux2to10_not0;
  assign f_s_cska32_xor4 = a[4] ^ b[4];
  assign f_s_cska32_fa3_xor0 = a[4] ^ b[4];
  assign f_s_cska32_fa3_and0 = a[4] & b[4];
  assign f_s_cska32_fa3_xor1 = f_s_cska32_fa3_xor0 ^ f_s_cska32_mux2to10_and1;
  assign f_s_cska32_fa3_and1 = f_s_cska32_fa3_xor0 & f_s_cska32_mux2to10_and1;
  assign f_s_cska32_fa3_or0 = f_s_cska32_fa3_and0 | f_s_cska32_fa3_and1;
  assign f_s_cska32_xor5 = a[5] ^ b[5];
  assign f_s_cska32_fa4_xor0 = a[5] ^ b[5];
  assign f_s_cska32_fa4_and0 = a[5] & b[5];
  assign f_s_cska32_fa4_xor1 = f_s_cska32_fa4_xor0 ^ f_s_cska32_fa3_or0;
  assign f_s_cska32_fa4_and1 = f_s_cska32_fa4_xor0 & f_s_cska32_fa3_or0;
  assign f_s_cska32_fa4_or0 = f_s_cska32_fa4_and0 | f_s_cska32_fa4_and1;
  assign f_s_cska32_xor6 = a[6] ^ b[6];
  assign f_s_cska32_fa5_xor0 = a[6] ^ b[6];
  assign f_s_cska32_fa5_and0 = a[6] & b[6];
  assign f_s_cska32_fa5_xor1 = f_s_cska32_fa5_xor0 ^ f_s_cska32_fa4_or0;
  assign f_s_cska32_fa5_and1 = f_s_cska32_fa5_xor0 & f_s_cska32_fa4_or0;
  assign f_s_cska32_fa5_or0 = f_s_cska32_fa5_and0 | f_s_cska32_fa5_and1;
  assign f_s_cska32_xor7 = a[7] ^ b[7];
  assign f_s_cska32_fa6_xor0 = a[7] ^ b[7];
  assign f_s_cska32_fa6_and0 = a[7] & b[7];
  assign f_s_cska32_fa6_xor1 = f_s_cska32_fa6_xor0 ^ f_s_cska32_fa5_or0;
  assign f_s_cska32_fa6_and1 = f_s_cska32_fa6_xor0 & f_s_cska32_fa5_or0;
  assign f_s_cska32_fa6_or0 = f_s_cska32_fa6_and0 | f_s_cska32_fa6_and1;
  assign f_s_cska32_and_propagate13 = f_s_cska32_xor4 & f_s_cska32_xor6;
  assign f_s_cska32_and_propagate14 = f_s_cska32_xor5 & f_s_cska32_xor7;
  assign f_s_cska32_and_propagate15 = f_s_cska32_and_propagate13 & f_s_cska32_and_propagate14;
  assign f_s_cska32_mux2to11_and0 = f_s_cska32_mux2to10_and1 & f_s_cska32_and_propagate15;
  assign f_s_cska32_mux2to11_not0 = ~f_s_cska32_and_propagate15;
  assign f_s_cska32_mux2to11_and1 = f_s_cska32_fa6_or0 & f_s_cska32_mux2to11_not0;
  assign f_s_cska32_mux2to11_xor0 = f_s_cska32_mux2to11_and0 ^ f_s_cska32_mux2to11_and1;
  assign f_s_cska32_xor8 = a[8] ^ b[8];
  assign f_s_cska32_fa7_xor0 = a[8] ^ b[8];
  assign f_s_cska32_fa7_and0 = a[8] & b[8];
  assign f_s_cska32_fa7_xor1 = f_s_cska32_fa7_xor0 ^ f_s_cska32_mux2to11_xor0;
  assign f_s_cska32_fa7_and1 = f_s_cska32_fa7_xor0 & f_s_cska32_mux2to11_xor0;
  assign f_s_cska32_fa7_or0 = f_s_cska32_fa7_and0 | f_s_cska32_fa7_and1;
  assign f_s_cska32_xor9 = a[9] ^ b[9];
  assign f_s_cska32_fa8_xor0 = a[9] ^ b[9];
  assign f_s_cska32_fa8_and0 = a[9] & b[9];
  assign f_s_cska32_fa8_xor1 = f_s_cska32_fa8_xor0 ^ f_s_cska32_fa7_or0;
  assign f_s_cska32_fa8_and1 = f_s_cska32_fa8_xor0 & f_s_cska32_fa7_or0;
  assign f_s_cska32_fa8_or0 = f_s_cska32_fa8_and0 | f_s_cska32_fa8_and1;
  assign f_s_cska32_xor10 = a[10] ^ b[10];
  assign f_s_cska32_fa9_xor0 = a[10] ^ b[10];
  assign f_s_cska32_fa9_and0 = a[10] & b[10];
  assign f_s_cska32_fa9_xor1 = f_s_cska32_fa9_xor0 ^ f_s_cska32_fa8_or0;
  assign f_s_cska32_fa9_and1 = f_s_cska32_fa9_xor0 & f_s_cska32_fa8_or0;
  assign f_s_cska32_fa9_or0 = f_s_cska32_fa9_and0 | f_s_cska32_fa9_and1;
  assign f_s_cska32_xor11 = a[11] ^ b[11];
  assign f_s_cska32_fa10_xor0 = a[11] ^ b[11];
  assign f_s_cska32_fa10_and0 = a[11] & b[11];
  assign f_s_cska32_fa10_xor1 = f_s_cska32_fa10_xor0 ^ f_s_cska32_fa9_or0;
  assign f_s_cska32_fa10_and1 = f_s_cska32_fa10_xor0 & f_s_cska32_fa9_or0;
  assign f_s_cska32_fa10_or0 = f_s_cska32_fa10_and0 | f_s_cska32_fa10_and1;
  assign f_s_cska32_and_propagate26 = f_s_cska32_xor8 & f_s_cska32_xor10;
  assign f_s_cska32_and_propagate27 = f_s_cska32_xor9 & f_s_cska32_xor11;
  assign f_s_cska32_and_propagate28 = f_s_cska32_and_propagate26 & f_s_cska32_and_propagate27;
  assign f_s_cska32_mux2to12_and0 = f_s_cska32_mux2to11_xor0 & f_s_cska32_and_propagate28;
  assign f_s_cska32_mux2to12_not0 = ~f_s_cska32_and_propagate28;
  assign f_s_cska32_mux2to12_and1 = f_s_cska32_fa10_or0 & f_s_cska32_mux2to12_not0;
  assign f_s_cska32_mux2to12_xor0 = f_s_cska32_mux2to12_and0 ^ f_s_cska32_mux2to12_and1;
  assign f_s_cska32_xor12 = a[12] ^ b[12];
  assign f_s_cska32_fa11_xor0 = a[12] ^ b[12];
  assign f_s_cska32_fa11_and0 = a[12] & b[12];
  assign f_s_cska32_fa11_xor1 = f_s_cska32_fa11_xor0 ^ f_s_cska32_mux2to12_xor0;
  assign f_s_cska32_fa11_and1 = f_s_cska32_fa11_xor0 & f_s_cska32_mux2to12_xor0;
  assign f_s_cska32_fa11_or0 = f_s_cska32_fa11_and0 | f_s_cska32_fa11_and1;
  assign f_s_cska32_xor13 = a[13] ^ b[13];
  assign f_s_cska32_fa12_xor0 = a[13] ^ b[13];
  assign f_s_cska32_fa12_and0 = a[13] & b[13];
  assign f_s_cska32_fa12_xor1 = f_s_cska32_fa12_xor0 ^ f_s_cska32_fa11_or0;
  assign f_s_cska32_fa12_and1 = f_s_cska32_fa12_xor0 & f_s_cska32_fa11_or0;
  assign f_s_cska32_fa12_or0 = f_s_cska32_fa12_and0 | f_s_cska32_fa12_and1;
  assign f_s_cska32_xor14 = a[14] ^ b[14];
  assign f_s_cska32_fa13_xor0 = a[14] ^ b[14];
  assign f_s_cska32_fa13_and0 = a[14] & b[14];
  assign f_s_cska32_fa13_xor1 = f_s_cska32_fa13_xor0 ^ f_s_cska32_fa12_or0;
  assign f_s_cska32_fa13_and1 = f_s_cska32_fa13_xor0 & f_s_cska32_fa12_or0;
  assign f_s_cska32_fa13_or0 = f_s_cska32_fa13_and0 | f_s_cska32_fa13_and1;
  assign f_s_cska32_xor15 = a[15] ^ b[15];
  assign f_s_cska32_fa14_xor0 = a[15] ^ b[15];
  assign f_s_cska32_fa14_and0 = a[15] & b[15];
  assign f_s_cska32_fa14_xor1 = f_s_cska32_fa14_xor0 ^ f_s_cska32_fa13_or0;
  assign f_s_cska32_fa14_and1 = f_s_cska32_fa14_xor0 & f_s_cska32_fa13_or0;
  assign f_s_cska32_fa14_or0 = f_s_cska32_fa14_and0 | f_s_cska32_fa14_and1;
  assign f_s_cska32_and_propagate39 = f_s_cska32_xor12 & f_s_cska32_xor14;
  assign f_s_cska32_and_propagate310 = f_s_cska32_xor13 & f_s_cska32_xor15;
  assign f_s_cska32_and_propagate311 = f_s_cska32_and_propagate39 & f_s_cska32_and_propagate310;
  assign f_s_cska32_mux2to13_and0 = f_s_cska32_mux2to12_xor0 & f_s_cska32_and_propagate311;
  assign f_s_cska32_mux2to13_not0 = ~f_s_cska32_and_propagate311;
  assign f_s_cska32_mux2to13_and1 = f_s_cska32_fa14_or0 & f_s_cska32_mux2to13_not0;
  assign f_s_cska32_mux2to13_xor0 = f_s_cska32_mux2to13_and0 ^ f_s_cska32_mux2to13_and1;
  assign f_s_cska32_xor16 = a[16] ^ b[16];
  assign f_s_cska32_fa15_xor0 = a[16] ^ b[16];
  assign f_s_cska32_fa15_and0 = a[16] & b[16];
  assign f_s_cska32_fa15_xor1 = f_s_cska32_fa15_xor0 ^ f_s_cska32_mux2to13_xor0;
  assign f_s_cska32_fa15_and1 = f_s_cska32_fa15_xor0 & f_s_cska32_mux2to13_xor0;
  assign f_s_cska32_fa15_or0 = f_s_cska32_fa15_and0 | f_s_cska32_fa15_and1;
  assign f_s_cska32_xor17 = a[17] ^ b[17];
  assign f_s_cska32_fa16_xor0 = a[17] ^ b[17];
  assign f_s_cska32_fa16_and0 = a[17] & b[17];
  assign f_s_cska32_fa16_xor1 = f_s_cska32_fa16_xor0 ^ f_s_cska32_fa15_or0;
  assign f_s_cska32_fa16_and1 = f_s_cska32_fa16_xor0 & f_s_cska32_fa15_or0;
  assign f_s_cska32_fa16_or0 = f_s_cska32_fa16_and0 | f_s_cska32_fa16_and1;
  assign f_s_cska32_xor18 = a[18] ^ b[18];
  assign f_s_cska32_fa17_xor0 = a[18] ^ b[18];
  assign f_s_cska32_fa17_and0 = a[18] & b[18];
  assign f_s_cska32_fa17_xor1 = f_s_cska32_fa17_xor0 ^ f_s_cska32_fa16_or0;
  assign f_s_cska32_fa17_and1 = f_s_cska32_fa17_xor0 & f_s_cska32_fa16_or0;
  assign f_s_cska32_fa17_or0 = f_s_cska32_fa17_and0 | f_s_cska32_fa17_and1;
  assign f_s_cska32_xor19 = a[19] ^ b[19];
  assign f_s_cska32_fa18_xor0 = a[19] ^ b[19];
  assign f_s_cska32_fa18_and0 = a[19] & b[19];
  assign f_s_cska32_fa18_xor1 = f_s_cska32_fa18_xor0 ^ f_s_cska32_fa17_or0;
  assign f_s_cska32_fa18_and1 = f_s_cska32_fa18_xor0 & f_s_cska32_fa17_or0;
  assign f_s_cska32_fa18_or0 = f_s_cska32_fa18_and0 | f_s_cska32_fa18_and1;
  assign f_s_cska32_and_propagate412 = f_s_cska32_xor16 & f_s_cska32_xor18;
  assign f_s_cska32_and_propagate413 = f_s_cska32_xor17 & f_s_cska32_xor19;
  assign f_s_cska32_and_propagate414 = f_s_cska32_and_propagate412 & f_s_cska32_and_propagate413;
  assign f_s_cska32_mux2to14_and0 = f_s_cska32_mux2to13_xor0 & f_s_cska32_and_propagate414;
  assign f_s_cska32_mux2to14_not0 = ~f_s_cska32_and_propagate414;
  assign f_s_cska32_mux2to14_and1 = f_s_cska32_fa18_or0 & f_s_cska32_mux2to14_not0;
  assign f_s_cska32_mux2to14_xor0 = f_s_cska32_mux2to14_and0 ^ f_s_cska32_mux2to14_and1;
  assign f_s_cska32_xor20 = a[20] ^ b[20];
  assign f_s_cska32_fa19_xor0 = a[20] ^ b[20];
  assign f_s_cska32_fa19_and0 = a[20] & b[20];
  assign f_s_cska32_fa19_xor1 = f_s_cska32_fa19_xor0 ^ f_s_cska32_mux2to14_xor0;
  assign f_s_cska32_fa19_and1 = f_s_cska32_fa19_xor0 & f_s_cska32_mux2to14_xor0;
  assign f_s_cska32_fa19_or0 = f_s_cska32_fa19_and0 | f_s_cska32_fa19_and1;
  assign f_s_cska32_xor21 = a[21] ^ b[21];
  assign f_s_cska32_fa20_xor0 = a[21] ^ b[21];
  assign f_s_cska32_fa20_and0 = a[21] & b[21];
  assign f_s_cska32_fa20_xor1 = f_s_cska32_fa20_xor0 ^ f_s_cska32_fa19_or0;
  assign f_s_cska32_fa20_and1 = f_s_cska32_fa20_xor0 & f_s_cska32_fa19_or0;
  assign f_s_cska32_fa20_or0 = f_s_cska32_fa20_and0 | f_s_cska32_fa20_and1;
  assign f_s_cska32_xor22 = a[22] ^ b[22];
  assign f_s_cska32_fa21_xor0 = a[22] ^ b[22];
  assign f_s_cska32_fa21_and0 = a[22] & b[22];
  assign f_s_cska32_fa21_xor1 = f_s_cska32_fa21_xor0 ^ f_s_cska32_fa20_or0;
  assign f_s_cska32_fa21_and1 = f_s_cska32_fa21_xor0 & f_s_cska32_fa20_or0;
  assign f_s_cska32_fa21_or0 = f_s_cska32_fa21_and0 | f_s_cska32_fa21_and1;
  assign f_s_cska32_xor23 = a[23] ^ b[23];
  assign f_s_cska32_fa22_xor0 = a[23] ^ b[23];
  assign f_s_cska32_fa22_and0 = a[23] & b[23];
  assign f_s_cska32_fa22_xor1 = f_s_cska32_fa22_xor0 ^ f_s_cska32_fa21_or0;
  assign f_s_cska32_fa22_and1 = f_s_cska32_fa22_xor0 & f_s_cska32_fa21_or0;
  assign f_s_cska32_fa22_or0 = f_s_cska32_fa22_and0 | f_s_cska32_fa22_and1;
  assign f_s_cska32_and_propagate515 = f_s_cska32_xor20 & f_s_cska32_xor22;
  assign f_s_cska32_and_propagate516 = f_s_cska32_xor21 & f_s_cska32_xor23;
  assign f_s_cska32_and_propagate517 = f_s_cska32_and_propagate515 & f_s_cska32_and_propagate516;
  assign f_s_cska32_mux2to15_and0 = f_s_cska32_mux2to14_xor0 & f_s_cska32_and_propagate517;
  assign f_s_cska32_mux2to15_not0 = ~f_s_cska32_and_propagate517;
  assign f_s_cska32_mux2to15_and1 = f_s_cska32_fa22_or0 & f_s_cska32_mux2to15_not0;
  assign f_s_cska32_mux2to15_xor0 = f_s_cska32_mux2to15_and0 ^ f_s_cska32_mux2to15_and1;
  assign f_s_cska32_xor24 = a[24] ^ b[24];
  assign f_s_cska32_fa23_xor0 = a[24] ^ b[24];
  assign f_s_cska32_fa23_and0 = a[24] & b[24];
  assign f_s_cska32_fa23_xor1 = f_s_cska32_fa23_xor0 ^ f_s_cska32_mux2to15_xor0;
  assign f_s_cska32_fa23_and1 = f_s_cska32_fa23_xor0 & f_s_cska32_mux2to15_xor0;
  assign f_s_cska32_fa23_or0 = f_s_cska32_fa23_and0 | f_s_cska32_fa23_and1;
  assign f_s_cska32_xor25 = a[25] ^ b[25];
  assign f_s_cska32_fa24_xor0 = a[25] ^ b[25];
  assign f_s_cska32_fa24_and0 = a[25] & b[25];
  assign f_s_cska32_fa24_xor1 = f_s_cska32_fa24_xor0 ^ f_s_cska32_fa23_or0;
  assign f_s_cska32_fa24_and1 = f_s_cska32_fa24_xor0 & f_s_cska32_fa23_or0;
  assign f_s_cska32_fa24_or0 = f_s_cska32_fa24_and0 | f_s_cska32_fa24_and1;
  assign f_s_cska32_xor26 = a[26] ^ b[26];
  assign f_s_cska32_fa25_xor0 = a[26] ^ b[26];
  assign f_s_cska32_fa25_and0 = a[26] & b[26];
  assign f_s_cska32_fa25_xor1 = f_s_cska32_fa25_xor0 ^ f_s_cska32_fa24_or0;
  assign f_s_cska32_fa25_and1 = f_s_cska32_fa25_xor0 & f_s_cska32_fa24_or0;
  assign f_s_cska32_fa25_or0 = f_s_cska32_fa25_and0 | f_s_cska32_fa25_and1;
  assign f_s_cska32_xor27 = a[27] ^ b[27];
  assign f_s_cska32_fa26_xor0 = a[27] ^ b[27];
  assign f_s_cska32_fa26_and0 = a[27] & b[27];
  assign f_s_cska32_fa26_xor1 = f_s_cska32_fa26_xor0 ^ f_s_cska32_fa25_or0;
  assign f_s_cska32_fa26_and1 = f_s_cska32_fa26_xor0 & f_s_cska32_fa25_or0;
  assign f_s_cska32_fa26_or0 = f_s_cska32_fa26_and0 | f_s_cska32_fa26_and1;
  assign f_s_cska32_and_propagate618 = f_s_cska32_xor24 & f_s_cska32_xor26;
  assign f_s_cska32_and_propagate619 = f_s_cska32_xor25 & f_s_cska32_xor27;
  assign f_s_cska32_and_propagate620 = f_s_cska32_and_propagate618 & f_s_cska32_and_propagate619;
  assign f_s_cska32_mux2to16_and0 = f_s_cska32_mux2to15_xor0 & f_s_cska32_and_propagate620;
  assign f_s_cska32_mux2to16_not0 = ~f_s_cska32_and_propagate620;
  assign f_s_cska32_mux2to16_and1 = f_s_cska32_fa26_or0 & f_s_cska32_mux2to16_not0;
  assign f_s_cska32_mux2to16_xor0 = f_s_cska32_mux2to16_and0 ^ f_s_cska32_mux2to16_and1;
  assign f_s_cska32_xor28 = a[28] ^ b[28];
  assign f_s_cska32_fa27_xor0 = a[28] ^ b[28];
  assign f_s_cska32_fa27_and0 = a[28] & b[28];
  assign f_s_cska32_fa27_xor1 = f_s_cska32_fa27_xor0 ^ f_s_cska32_mux2to16_xor0;
  assign f_s_cska32_fa27_and1 = f_s_cska32_fa27_xor0 & f_s_cska32_mux2to16_xor0;
  assign f_s_cska32_fa27_or0 = f_s_cska32_fa27_and0 | f_s_cska32_fa27_and1;
  assign f_s_cska32_xor29 = a[29] ^ b[29];
  assign f_s_cska32_fa28_xor0 = a[29] ^ b[29];
  assign f_s_cska32_fa28_and0 = a[29] & b[29];
  assign f_s_cska32_fa28_xor1 = f_s_cska32_fa28_xor0 ^ f_s_cska32_fa27_or0;
  assign f_s_cska32_fa28_and1 = f_s_cska32_fa28_xor0 & f_s_cska32_fa27_or0;
  assign f_s_cska32_fa28_or0 = f_s_cska32_fa28_and0 | f_s_cska32_fa28_and1;
  assign f_s_cska32_xor30 = a[30] ^ b[30];
  assign f_s_cska32_fa29_xor0 = a[30] ^ b[30];
  assign f_s_cska32_fa29_and0 = a[30] & b[30];
  assign f_s_cska32_fa29_xor1 = f_s_cska32_fa29_xor0 ^ f_s_cska32_fa28_or0;
  assign f_s_cska32_fa29_and1 = f_s_cska32_fa29_xor0 & f_s_cska32_fa28_or0;
  assign f_s_cska32_fa29_or0 = f_s_cska32_fa29_and0 | f_s_cska32_fa29_and1;
  assign f_s_cska32_xor31 = a[31] ^ b[31];
  assign f_s_cska32_fa30_xor0 = a[31] ^ b[31];
  assign f_s_cska32_fa30_and0 = a[31] & b[31];
  assign f_s_cska32_fa30_xor1 = f_s_cska32_fa30_xor0 ^ f_s_cska32_fa29_or0;
  assign f_s_cska32_fa30_and1 = f_s_cska32_fa30_xor0 & f_s_cska32_fa29_or0;
  assign f_s_cska32_fa30_or0 = f_s_cska32_fa30_and0 | f_s_cska32_fa30_and1;
  assign f_s_cska32_and_propagate721 = f_s_cska32_xor28 & f_s_cska32_xor30;
  assign f_s_cska32_and_propagate722 = f_s_cska32_xor29 & f_s_cska32_xor31;
  assign f_s_cska32_and_propagate723 = f_s_cska32_and_propagate721 & f_s_cska32_and_propagate722;
  assign f_s_cska32_mux2to17_and0 = f_s_cska32_mux2to16_xor0 & f_s_cska32_and_propagate723;
  assign f_s_cska32_mux2to17_not0 = ~f_s_cska32_and_propagate723;
  assign f_s_cska32_mux2to17_and1 = f_s_cska32_fa30_or0 & f_s_cska32_mux2to17_not0;
  assign f_s_cska32_mux2to17_xor0 = f_s_cska32_mux2to17_and0 ^ f_s_cska32_mux2to17_and1;
  assign f_s_cska32_xor32 = a[31] ^ b[31];
  assign f_s_cska32_xor33 = f_s_cska32_xor32 ^ f_s_cska32_mux2to17_xor0;

  assign f_s_cska32_out[0] = f_s_cska32_ha0_xor0;
  assign f_s_cska32_out[1] = f_s_cska32_fa0_xor1;
  assign f_s_cska32_out[2] = f_s_cska32_fa1_xor1;
  assign f_s_cska32_out[3] = f_s_cska32_fa2_xor1;
  assign f_s_cska32_out[4] = f_s_cska32_fa3_xor1;
  assign f_s_cska32_out[5] = f_s_cska32_fa4_xor1;
  assign f_s_cska32_out[6] = f_s_cska32_fa5_xor1;
  assign f_s_cska32_out[7] = f_s_cska32_fa6_xor1;
  assign f_s_cska32_out[8] = f_s_cska32_fa7_xor1;
  assign f_s_cska32_out[9] = f_s_cska32_fa8_xor1;
  assign f_s_cska32_out[10] = f_s_cska32_fa9_xor1;
  assign f_s_cska32_out[11] = f_s_cska32_fa10_xor1;
  assign f_s_cska32_out[12] = f_s_cska32_fa11_xor1;
  assign f_s_cska32_out[13] = f_s_cska32_fa12_xor1;
  assign f_s_cska32_out[14] = f_s_cska32_fa13_xor1;
  assign f_s_cska32_out[15] = f_s_cska32_fa14_xor1;
  assign f_s_cska32_out[16] = f_s_cska32_fa15_xor1;
  assign f_s_cska32_out[17] = f_s_cska32_fa16_xor1;
  assign f_s_cska32_out[18] = f_s_cska32_fa17_xor1;
  assign f_s_cska32_out[19] = f_s_cska32_fa18_xor1;
  assign f_s_cska32_out[20] = f_s_cska32_fa19_xor1;
  assign f_s_cska32_out[21] = f_s_cska32_fa20_xor1;
  assign f_s_cska32_out[22] = f_s_cska32_fa21_xor1;
  assign f_s_cska32_out[23] = f_s_cska32_fa22_xor1;
  assign f_s_cska32_out[24] = f_s_cska32_fa23_xor1;
  assign f_s_cska32_out[25] = f_s_cska32_fa24_xor1;
  assign f_s_cska32_out[26] = f_s_cska32_fa25_xor1;
  assign f_s_cska32_out[27] = f_s_cska32_fa26_xor1;
  assign f_s_cska32_out[28] = f_s_cska32_fa27_xor1;
  assign f_s_cska32_out[29] = f_s_cska32_fa28_xor1;
  assign f_s_cska32_out[30] = f_s_cska32_fa29_xor1;
  assign f_s_cska32_out[31] = f_s_cska32_fa30_xor1;
  assign f_s_cska32_out[32] = f_s_cska32_xor33;
endmodule