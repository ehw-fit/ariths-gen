module u_pg_rca32(input [31:0] a, input [31:0] b, output [32:0] u_pg_rca32_out);
  wire u_pg_rca32_pg_fa0_xor0;
  wire u_pg_rca32_pg_fa0_and0;
  wire u_pg_rca32_pg_fa1_xor0;
  wire u_pg_rca32_pg_fa1_and0;
  wire u_pg_rca32_pg_fa1_xor1;
  wire u_pg_rca32_and1;
  wire u_pg_rca32_or1;
  wire u_pg_rca32_pg_fa2_xor0;
  wire u_pg_rca32_pg_fa2_and0;
  wire u_pg_rca32_pg_fa2_xor1;
  wire u_pg_rca32_and2;
  wire u_pg_rca32_or2;
  wire u_pg_rca32_pg_fa3_xor0;
  wire u_pg_rca32_pg_fa3_and0;
  wire u_pg_rca32_pg_fa3_xor1;
  wire u_pg_rca32_and3;
  wire u_pg_rca32_or3;
  wire u_pg_rca32_pg_fa4_xor0;
  wire u_pg_rca32_pg_fa4_and0;
  wire u_pg_rca32_pg_fa4_xor1;
  wire u_pg_rca32_and4;
  wire u_pg_rca32_or4;
  wire u_pg_rca32_pg_fa5_xor0;
  wire u_pg_rca32_pg_fa5_and0;
  wire u_pg_rca32_pg_fa5_xor1;
  wire u_pg_rca32_and5;
  wire u_pg_rca32_or5;
  wire u_pg_rca32_pg_fa6_xor0;
  wire u_pg_rca32_pg_fa6_and0;
  wire u_pg_rca32_pg_fa6_xor1;
  wire u_pg_rca32_and6;
  wire u_pg_rca32_or6;
  wire u_pg_rca32_pg_fa7_xor0;
  wire u_pg_rca32_pg_fa7_and0;
  wire u_pg_rca32_pg_fa7_xor1;
  wire u_pg_rca32_and7;
  wire u_pg_rca32_or7;
  wire u_pg_rca32_pg_fa8_xor0;
  wire u_pg_rca32_pg_fa8_and0;
  wire u_pg_rca32_pg_fa8_xor1;
  wire u_pg_rca32_and8;
  wire u_pg_rca32_or8;
  wire u_pg_rca32_pg_fa9_xor0;
  wire u_pg_rca32_pg_fa9_and0;
  wire u_pg_rca32_pg_fa9_xor1;
  wire u_pg_rca32_and9;
  wire u_pg_rca32_or9;
  wire u_pg_rca32_pg_fa10_xor0;
  wire u_pg_rca32_pg_fa10_and0;
  wire u_pg_rca32_pg_fa10_xor1;
  wire u_pg_rca32_and10;
  wire u_pg_rca32_or10;
  wire u_pg_rca32_pg_fa11_xor0;
  wire u_pg_rca32_pg_fa11_and0;
  wire u_pg_rca32_pg_fa11_xor1;
  wire u_pg_rca32_and11;
  wire u_pg_rca32_or11;
  wire u_pg_rca32_pg_fa12_xor0;
  wire u_pg_rca32_pg_fa12_and0;
  wire u_pg_rca32_pg_fa12_xor1;
  wire u_pg_rca32_and12;
  wire u_pg_rca32_or12;
  wire u_pg_rca32_pg_fa13_xor0;
  wire u_pg_rca32_pg_fa13_and0;
  wire u_pg_rca32_pg_fa13_xor1;
  wire u_pg_rca32_and13;
  wire u_pg_rca32_or13;
  wire u_pg_rca32_pg_fa14_xor0;
  wire u_pg_rca32_pg_fa14_and0;
  wire u_pg_rca32_pg_fa14_xor1;
  wire u_pg_rca32_and14;
  wire u_pg_rca32_or14;
  wire u_pg_rca32_pg_fa15_xor0;
  wire u_pg_rca32_pg_fa15_and0;
  wire u_pg_rca32_pg_fa15_xor1;
  wire u_pg_rca32_and15;
  wire u_pg_rca32_or15;
  wire u_pg_rca32_pg_fa16_xor0;
  wire u_pg_rca32_pg_fa16_and0;
  wire u_pg_rca32_pg_fa16_xor1;
  wire u_pg_rca32_and16;
  wire u_pg_rca32_or16;
  wire u_pg_rca32_pg_fa17_xor0;
  wire u_pg_rca32_pg_fa17_and0;
  wire u_pg_rca32_pg_fa17_xor1;
  wire u_pg_rca32_and17;
  wire u_pg_rca32_or17;
  wire u_pg_rca32_pg_fa18_xor0;
  wire u_pg_rca32_pg_fa18_and0;
  wire u_pg_rca32_pg_fa18_xor1;
  wire u_pg_rca32_and18;
  wire u_pg_rca32_or18;
  wire u_pg_rca32_pg_fa19_xor0;
  wire u_pg_rca32_pg_fa19_and0;
  wire u_pg_rca32_pg_fa19_xor1;
  wire u_pg_rca32_and19;
  wire u_pg_rca32_or19;
  wire u_pg_rca32_pg_fa20_xor0;
  wire u_pg_rca32_pg_fa20_and0;
  wire u_pg_rca32_pg_fa20_xor1;
  wire u_pg_rca32_and20;
  wire u_pg_rca32_or20;
  wire u_pg_rca32_pg_fa21_xor0;
  wire u_pg_rca32_pg_fa21_and0;
  wire u_pg_rca32_pg_fa21_xor1;
  wire u_pg_rca32_and21;
  wire u_pg_rca32_or21;
  wire u_pg_rca32_pg_fa22_xor0;
  wire u_pg_rca32_pg_fa22_and0;
  wire u_pg_rca32_pg_fa22_xor1;
  wire u_pg_rca32_and22;
  wire u_pg_rca32_or22;
  wire u_pg_rca32_pg_fa23_xor0;
  wire u_pg_rca32_pg_fa23_and0;
  wire u_pg_rca32_pg_fa23_xor1;
  wire u_pg_rca32_and23;
  wire u_pg_rca32_or23;
  wire u_pg_rca32_pg_fa24_xor0;
  wire u_pg_rca32_pg_fa24_and0;
  wire u_pg_rca32_pg_fa24_xor1;
  wire u_pg_rca32_and24;
  wire u_pg_rca32_or24;
  wire u_pg_rca32_pg_fa25_xor0;
  wire u_pg_rca32_pg_fa25_and0;
  wire u_pg_rca32_pg_fa25_xor1;
  wire u_pg_rca32_and25;
  wire u_pg_rca32_or25;
  wire u_pg_rca32_pg_fa26_xor0;
  wire u_pg_rca32_pg_fa26_and0;
  wire u_pg_rca32_pg_fa26_xor1;
  wire u_pg_rca32_and26;
  wire u_pg_rca32_or26;
  wire u_pg_rca32_pg_fa27_xor0;
  wire u_pg_rca32_pg_fa27_and0;
  wire u_pg_rca32_pg_fa27_xor1;
  wire u_pg_rca32_and27;
  wire u_pg_rca32_or27;
  wire u_pg_rca32_pg_fa28_xor0;
  wire u_pg_rca32_pg_fa28_and0;
  wire u_pg_rca32_pg_fa28_xor1;
  wire u_pg_rca32_and28;
  wire u_pg_rca32_or28;
  wire u_pg_rca32_pg_fa29_xor0;
  wire u_pg_rca32_pg_fa29_and0;
  wire u_pg_rca32_pg_fa29_xor1;
  wire u_pg_rca32_and29;
  wire u_pg_rca32_or29;
  wire u_pg_rca32_pg_fa30_xor0;
  wire u_pg_rca32_pg_fa30_and0;
  wire u_pg_rca32_pg_fa30_xor1;
  wire u_pg_rca32_and30;
  wire u_pg_rca32_or30;
  wire u_pg_rca32_pg_fa31_xor0;
  wire u_pg_rca32_pg_fa31_and0;
  wire u_pg_rca32_pg_fa31_xor1;
  wire u_pg_rca32_and31;
  wire u_pg_rca32_or31;

  assign u_pg_rca32_pg_fa0_xor0 = a[0] ^ b[0];
  assign u_pg_rca32_pg_fa0_and0 = a[0] & b[0];
  assign u_pg_rca32_pg_fa1_xor0 = a[1] ^ b[1];
  assign u_pg_rca32_pg_fa1_and0 = a[1] & b[1];
  assign u_pg_rca32_pg_fa1_xor1 = u_pg_rca32_pg_fa1_xor0 ^ u_pg_rca32_pg_fa0_and0;
  assign u_pg_rca32_and1 = u_pg_rca32_pg_fa0_and0 & u_pg_rca32_pg_fa1_xor0;
  assign u_pg_rca32_or1 = u_pg_rca32_and1 | u_pg_rca32_pg_fa1_and0;
  assign u_pg_rca32_pg_fa2_xor0 = a[2] ^ b[2];
  assign u_pg_rca32_pg_fa2_and0 = a[2] & b[2];
  assign u_pg_rca32_pg_fa2_xor1 = u_pg_rca32_pg_fa2_xor0 ^ u_pg_rca32_or1;
  assign u_pg_rca32_and2 = u_pg_rca32_or1 & u_pg_rca32_pg_fa2_xor0;
  assign u_pg_rca32_or2 = u_pg_rca32_and2 | u_pg_rca32_pg_fa2_and0;
  assign u_pg_rca32_pg_fa3_xor0 = a[3] ^ b[3];
  assign u_pg_rca32_pg_fa3_and0 = a[3] & b[3];
  assign u_pg_rca32_pg_fa3_xor1 = u_pg_rca32_pg_fa3_xor0 ^ u_pg_rca32_or2;
  assign u_pg_rca32_and3 = u_pg_rca32_or2 & u_pg_rca32_pg_fa3_xor0;
  assign u_pg_rca32_or3 = u_pg_rca32_and3 | u_pg_rca32_pg_fa3_and0;
  assign u_pg_rca32_pg_fa4_xor0 = a[4] ^ b[4];
  assign u_pg_rca32_pg_fa4_and0 = a[4] & b[4];
  assign u_pg_rca32_pg_fa4_xor1 = u_pg_rca32_pg_fa4_xor0 ^ u_pg_rca32_or3;
  assign u_pg_rca32_and4 = u_pg_rca32_or3 & u_pg_rca32_pg_fa4_xor0;
  assign u_pg_rca32_or4 = u_pg_rca32_and4 | u_pg_rca32_pg_fa4_and0;
  assign u_pg_rca32_pg_fa5_xor0 = a[5] ^ b[5];
  assign u_pg_rca32_pg_fa5_and0 = a[5] & b[5];
  assign u_pg_rca32_pg_fa5_xor1 = u_pg_rca32_pg_fa5_xor0 ^ u_pg_rca32_or4;
  assign u_pg_rca32_and5 = u_pg_rca32_or4 & u_pg_rca32_pg_fa5_xor0;
  assign u_pg_rca32_or5 = u_pg_rca32_and5 | u_pg_rca32_pg_fa5_and0;
  assign u_pg_rca32_pg_fa6_xor0 = a[6] ^ b[6];
  assign u_pg_rca32_pg_fa6_and0 = a[6] & b[6];
  assign u_pg_rca32_pg_fa6_xor1 = u_pg_rca32_pg_fa6_xor0 ^ u_pg_rca32_or5;
  assign u_pg_rca32_and6 = u_pg_rca32_or5 & u_pg_rca32_pg_fa6_xor0;
  assign u_pg_rca32_or6 = u_pg_rca32_and6 | u_pg_rca32_pg_fa6_and0;
  assign u_pg_rca32_pg_fa7_xor0 = a[7] ^ b[7];
  assign u_pg_rca32_pg_fa7_and0 = a[7] & b[7];
  assign u_pg_rca32_pg_fa7_xor1 = u_pg_rca32_pg_fa7_xor0 ^ u_pg_rca32_or6;
  assign u_pg_rca32_and7 = u_pg_rca32_or6 & u_pg_rca32_pg_fa7_xor0;
  assign u_pg_rca32_or7 = u_pg_rca32_and7 | u_pg_rca32_pg_fa7_and0;
  assign u_pg_rca32_pg_fa8_xor0 = a[8] ^ b[8];
  assign u_pg_rca32_pg_fa8_and0 = a[8] & b[8];
  assign u_pg_rca32_pg_fa8_xor1 = u_pg_rca32_pg_fa8_xor0 ^ u_pg_rca32_or7;
  assign u_pg_rca32_and8 = u_pg_rca32_or7 & u_pg_rca32_pg_fa8_xor0;
  assign u_pg_rca32_or8 = u_pg_rca32_and8 | u_pg_rca32_pg_fa8_and0;
  assign u_pg_rca32_pg_fa9_xor0 = a[9] ^ b[9];
  assign u_pg_rca32_pg_fa9_and0 = a[9] & b[9];
  assign u_pg_rca32_pg_fa9_xor1 = u_pg_rca32_pg_fa9_xor0 ^ u_pg_rca32_or8;
  assign u_pg_rca32_and9 = u_pg_rca32_or8 & u_pg_rca32_pg_fa9_xor0;
  assign u_pg_rca32_or9 = u_pg_rca32_and9 | u_pg_rca32_pg_fa9_and0;
  assign u_pg_rca32_pg_fa10_xor0 = a[10] ^ b[10];
  assign u_pg_rca32_pg_fa10_and0 = a[10] & b[10];
  assign u_pg_rca32_pg_fa10_xor1 = u_pg_rca32_pg_fa10_xor0 ^ u_pg_rca32_or9;
  assign u_pg_rca32_and10 = u_pg_rca32_or9 & u_pg_rca32_pg_fa10_xor0;
  assign u_pg_rca32_or10 = u_pg_rca32_and10 | u_pg_rca32_pg_fa10_and0;
  assign u_pg_rca32_pg_fa11_xor0 = a[11] ^ b[11];
  assign u_pg_rca32_pg_fa11_and0 = a[11] & b[11];
  assign u_pg_rca32_pg_fa11_xor1 = u_pg_rca32_pg_fa11_xor0 ^ u_pg_rca32_or10;
  assign u_pg_rca32_and11 = u_pg_rca32_or10 & u_pg_rca32_pg_fa11_xor0;
  assign u_pg_rca32_or11 = u_pg_rca32_and11 | u_pg_rca32_pg_fa11_and0;
  assign u_pg_rca32_pg_fa12_xor0 = a[12] ^ b[12];
  assign u_pg_rca32_pg_fa12_and0 = a[12] & b[12];
  assign u_pg_rca32_pg_fa12_xor1 = u_pg_rca32_pg_fa12_xor0 ^ u_pg_rca32_or11;
  assign u_pg_rca32_and12 = u_pg_rca32_or11 & u_pg_rca32_pg_fa12_xor0;
  assign u_pg_rca32_or12 = u_pg_rca32_and12 | u_pg_rca32_pg_fa12_and0;
  assign u_pg_rca32_pg_fa13_xor0 = a[13] ^ b[13];
  assign u_pg_rca32_pg_fa13_and0 = a[13] & b[13];
  assign u_pg_rca32_pg_fa13_xor1 = u_pg_rca32_pg_fa13_xor0 ^ u_pg_rca32_or12;
  assign u_pg_rca32_and13 = u_pg_rca32_or12 & u_pg_rca32_pg_fa13_xor0;
  assign u_pg_rca32_or13 = u_pg_rca32_and13 | u_pg_rca32_pg_fa13_and0;
  assign u_pg_rca32_pg_fa14_xor0 = a[14] ^ b[14];
  assign u_pg_rca32_pg_fa14_and0 = a[14] & b[14];
  assign u_pg_rca32_pg_fa14_xor1 = u_pg_rca32_pg_fa14_xor0 ^ u_pg_rca32_or13;
  assign u_pg_rca32_and14 = u_pg_rca32_or13 & u_pg_rca32_pg_fa14_xor0;
  assign u_pg_rca32_or14 = u_pg_rca32_and14 | u_pg_rca32_pg_fa14_and0;
  assign u_pg_rca32_pg_fa15_xor0 = a[15] ^ b[15];
  assign u_pg_rca32_pg_fa15_and0 = a[15] & b[15];
  assign u_pg_rca32_pg_fa15_xor1 = u_pg_rca32_pg_fa15_xor0 ^ u_pg_rca32_or14;
  assign u_pg_rca32_and15 = u_pg_rca32_or14 & u_pg_rca32_pg_fa15_xor0;
  assign u_pg_rca32_or15 = u_pg_rca32_and15 | u_pg_rca32_pg_fa15_and0;
  assign u_pg_rca32_pg_fa16_xor0 = a[16] ^ b[16];
  assign u_pg_rca32_pg_fa16_and0 = a[16] & b[16];
  assign u_pg_rca32_pg_fa16_xor1 = u_pg_rca32_pg_fa16_xor0 ^ u_pg_rca32_or15;
  assign u_pg_rca32_and16 = u_pg_rca32_or15 & u_pg_rca32_pg_fa16_xor0;
  assign u_pg_rca32_or16 = u_pg_rca32_and16 | u_pg_rca32_pg_fa16_and0;
  assign u_pg_rca32_pg_fa17_xor0 = a[17] ^ b[17];
  assign u_pg_rca32_pg_fa17_and0 = a[17] & b[17];
  assign u_pg_rca32_pg_fa17_xor1 = u_pg_rca32_pg_fa17_xor0 ^ u_pg_rca32_or16;
  assign u_pg_rca32_and17 = u_pg_rca32_or16 & u_pg_rca32_pg_fa17_xor0;
  assign u_pg_rca32_or17 = u_pg_rca32_and17 | u_pg_rca32_pg_fa17_and0;
  assign u_pg_rca32_pg_fa18_xor0 = a[18] ^ b[18];
  assign u_pg_rca32_pg_fa18_and0 = a[18] & b[18];
  assign u_pg_rca32_pg_fa18_xor1 = u_pg_rca32_pg_fa18_xor0 ^ u_pg_rca32_or17;
  assign u_pg_rca32_and18 = u_pg_rca32_or17 & u_pg_rca32_pg_fa18_xor0;
  assign u_pg_rca32_or18 = u_pg_rca32_and18 | u_pg_rca32_pg_fa18_and0;
  assign u_pg_rca32_pg_fa19_xor0 = a[19] ^ b[19];
  assign u_pg_rca32_pg_fa19_and0 = a[19] & b[19];
  assign u_pg_rca32_pg_fa19_xor1 = u_pg_rca32_pg_fa19_xor0 ^ u_pg_rca32_or18;
  assign u_pg_rca32_and19 = u_pg_rca32_or18 & u_pg_rca32_pg_fa19_xor0;
  assign u_pg_rca32_or19 = u_pg_rca32_and19 | u_pg_rca32_pg_fa19_and0;
  assign u_pg_rca32_pg_fa20_xor0 = a[20] ^ b[20];
  assign u_pg_rca32_pg_fa20_and0 = a[20] & b[20];
  assign u_pg_rca32_pg_fa20_xor1 = u_pg_rca32_pg_fa20_xor0 ^ u_pg_rca32_or19;
  assign u_pg_rca32_and20 = u_pg_rca32_or19 & u_pg_rca32_pg_fa20_xor0;
  assign u_pg_rca32_or20 = u_pg_rca32_and20 | u_pg_rca32_pg_fa20_and0;
  assign u_pg_rca32_pg_fa21_xor0 = a[21] ^ b[21];
  assign u_pg_rca32_pg_fa21_and0 = a[21] & b[21];
  assign u_pg_rca32_pg_fa21_xor1 = u_pg_rca32_pg_fa21_xor0 ^ u_pg_rca32_or20;
  assign u_pg_rca32_and21 = u_pg_rca32_or20 & u_pg_rca32_pg_fa21_xor0;
  assign u_pg_rca32_or21 = u_pg_rca32_and21 | u_pg_rca32_pg_fa21_and0;
  assign u_pg_rca32_pg_fa22_xor0 = a[22] ^ b[22];
  assign u_pg_rca32_pg_fa22_and0 = a[22] & b[22];
  assign u_pg_rca32_pg_fa22_xor1 = u_pg_rca32_pg_fa22_xor0 ^ u_pg_rca32_or21;
  assign u_pg_rca32_and22 = u_pg_rca32_or21 & u_pg_rca32_pg_fa22_xor0;
  assign u_pg_rca32_or22 = u_pg_rca32_and22 | u_pg_rca32_pg_fa22_and0;
  assign u_pg_rca32_pg_fa23_xor0 = a[23] ^ b[23];
  assign u_pg_rca32_pg_fa23_and0 = a[23] & b[23];
  assign u_pg_rca32_pg_fa23_xor1 = u_pg_rca32_pg_fa23_xor0 ^ u_pg_rca32_or22;
  assign u_pg_rca32_and23 = u_pg_rca32_or22 & u_pg_rca32_pg_fa23_xor0;
  assign u_pg_rca32_or23 = u_pg_rca32_and23 | u_pg_rca32_pg_fa23_and0;
  assign u_pg_rca32_pg_fa24_xor0 = a[24] ^ b[24];
  assign u_pg_rca32_pg_fa24_and0 = a[24] & b[24];
  assign u_pg_rca32_pg_fa24_xor1 = u_pg_rca32_pg_fa24_xor0 ^ u_pg_rca32_or23;
  assign u_pg_rca32_and24 = u_pg_rca32_or23 & u_pg_rca32_pg_fa24_xor0;
  assign u_pg_rca32_or24 = u_pg_rca32_and24 | u_pg_rca32_pg_fa24_and0;
  assign u_pg_rca32_pg_fa25_xor0 = a[25] ^ b[25];
  assign u_pg_rca32_pg_fa25_and0 = a[25] & b[25];
  assign u_pg_rca32_pg_fa25_xor1 = u_pg_rca32_pg_fa25_xor0 ^ u_pg_rca32_or24;
  assign u_pg_rca32_and25 = u_pg_rca32_or24 & u_pg_rca32_pg_fa25_xor0;
  assign u_pg_rca32_or25 = u_pg_rca32_and25 | u_pg_rca32_pg_fa25_and0;
  assign u_pg_rca32_pg_fa26_xor0 = a[26] ^ b[26];
  assign u_pg_rca32_pg_fa26_and0 = a[26] & b[26];
  assign u_pg_rca32_pg_fa26_xor1 = u_pg_rca32_pg_fa26_xor0 ^ u_pg_rca32_or25;
  assign u_pg_rca32_and26 = u_pg_rca32_or25 & u_pg_rca32_pg_fa26_xor0;
  assign u_pg_rca32_or26 = u_pg_rca32_and26 | u_pg_rca32_pg_fa26_and0;
  assign u_pg_rca32_pg_fa27_xor0 = a[27] ^ b[27];
  assign u_pg_rca32_pg_fa27_and0 = a[27] & b[27];
  assign u_pg_rca32_pg_fa27_xor1 = u_pg_rca32_pg_fa27_xor0 ^ u_pg_rca32_or26;
  assign u_pg_rca32_and27 = u_pg_rca32_or26 & u_pg_rca32_pg_fa27_xor0;
  assign u_pg_rca32_or27 = u_pg_rca32_and27 | u_pg_rca32_pg_fa27_and0;
  assign u_pg_rca32_pg_fa28_xor0 = a[28] ^ b[28];
  assign u_pg_rca32_pg_fa28_and0 = a[28] & b[28];
  assign u_pg_rca32_pg_fa28_xor1 = u_pg_rca32_pg_fa28_xor0 ^ u_pg_rca32_or27;
  assign u_pg_rca32_and28 = u_pg_rca32_or27 & u_pg_rca32_pg_fa28_xor0;
  assign u_pg_rca32_or28 = u_pg_rca32_and28 | u_pg_rca32_pg_fa28_and0;
  assign u_pg_rca32_pg_fa29_xor0 = a[29] ^ b[29];
  assign u_pg_rca32_pg_fa29_and0 = a[29] & b[29];
  assign u_pg_rca32_pg_fa29_xor1 = u_pg_rca32_pg_fa29_xor0 ^ u_pg_rca32_or28;
  assign u_pg_rca32_and29 = u_pg_rca32_or28 & u_pg_rca32_pg_fa29_xor0;
  assign u_pg_rca32_or29 = u_pg_rca32_and29 | u_pg_rca32_pg_fa29_and0;
  assign u_pg_rca32_pg_fa30_xor0 = a[30] ^ b[30];
  assign u_pg_rca32_pg_fa30_and0 = a[30] & b[30];
  assign u_pg_rca32_pg_fa30_xor1 = u_pg_rca32_pg_fa30_xor0 ^ u_pg_rca32_or29;
  assign u_pg_rca32_and30 = u_pg_rca32_or29 & u_pg_rca32_pg_fa30_xor0;
  assign u_pg_rca32_or30 = u_pg_rca32_and30 | u_pg_rca32_pg_fa30_and0;
  assign u_pg_rca32_pg_fa31_xor0 = a[31] ^ b[31];
  assign u_pg_rca32_pg_fa31_and0 = a[31] & b[31];
  assign u_pg_rca32_pg_fa31_xor1 = u_pg_rca32_pg_fa31_xor0 ^ u_pg_rca32_or30;
  assign u_pg_rca32_and31 = u_pg_rca32_or30 & u_pg_rca32_pg_fa31_xor0;
  assign u_pg_rca32_or31 = u_pg_rca32_and31 | u_pg_rca32_pg_fa31_and0;

  assign u_pg_rca32_out[0] = u_pg_rca32_pg_fa0_xor0;
  assign u_pg_rca32_out[1] = u_pg_rca32_pg_fa1_xor1;
  assign u_pg_rca32_out[2] = u_pg_rca32_pg_fa2_xor1;
  assign u_pg_rca32_out[3] = u_pg_rca32_pg_fa3_xor1;
  assign u_pg_rca32_out[4] = u_pg_rca32_pg_fa4_xor1;
  assign u_pg_rca32_out[5] = u_pg_rca32_pg_fa5_xor1;
  assign u_pg_rca32_out[6] = u_pg_rca32_pg_fa6_xor1;
  assign u_pg_rca32_out[7] = u_pg_rca32_pg_fa7_xor1;
  assign u_pg_rca32_out[8] = u_pg_rca32_pg_fa8_xor1;
  assign u_pg_rca32_out[9] = u_pg_rca32_pg_fa9_xor1;
  assign u_pg_rca32_out[10] = u_pg_rca32_pg_fa10_xor1;
  assign u_pg_rca32_out[11] = u_pg_rca32_pg_fa11_xor1;
  assign u_pg_rca32_out[12] = u_pg_rca32_pg_fa12_xor1;
  assign u_pg_rca32_out[13] = u_pg_rca32_pg_fa13_xor1;
  assign u_pg_rca32_out[14] = u_pg_rca32_pg_fa14_xor1;
  assign u_pg_rca32_out[15] = u_pg_rca32_pg_fa15_xor1;
  assign u_pg_rca32_out[16] = u_pg_rca32_pg_fa16_xor1;
  assign u_pg_rca32_out[17] = u_pg_rca32_pg_fa17_xor1;
  assign u_pg_rca32_out[18] = u_pg_rca32_pg_fa18_xor1;
  assign u_pg_rca32_out[19] = u_pg_rca32_pg_fa19_xor1;
  assign u_pg_rca32_out[20] = u_pg_rca32_pg_fa20_xor1;
  assign u_pg_rca32_out[21] = u_pg_rca32_pg_fa21_xor1;
  assign u_pg_rca32_out[22] = u_pg_rca32_pg_fa22_xor1;
  assign u_pg_rca32_out[23] = u_pg_rca32_pg_fa23_xor1;
  assign u_pg_rca32_out[24] = u_pg_rca32_pg_fa24_xor1;
  assign u_pg_rca32_out[25] = u_pg_rca32_pg_fa25_xor1;
  assign u_pg_rca32_out[26] = u_pg_rca32_pg_fa26_xor1;
  assign u_pg_rca32_out[27] = u_pg_rca32_pg_fa27_xor1;
  assign u_pg_rca32_out[28] = u_pg_rca32_pg_fa28_xor1;
  assign u_pg_rca32_out[29] = u_pg_rca32_pg_fa29_xor1;
  assign u_pg_rca32_out[30] = u_pg_rca32_pg_fa30_xor1;
  assign u_pg_rca32_out[31] = u_pg_rca32_pg_fa31_xor1;
  assign u_pg_rca32_out[32] = u_pg_rca32_or31;
endmodule