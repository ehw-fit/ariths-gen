module s_CSAwallace_rca24(input [23:0] a, input [23:0] b, output [47:0] s_CSAwallace_rca24_out);
  wire s_CSAwallace_rca24_and_0_0;
  wire s_CSAwallace_rca24_and_1_0;
  wire s_CSAwallace_rca24_and_2_0;
  wire s_CSAwallace_rca24_and_3_0;
  wire s_CSAwallace_rca24_and_4_0;
  wire s_CSAwallace_rca24_and_5_0;
  wire s_CSAwallace_rca24_and_6_0;
  wire s_CSAwallace_rca24_and_7_0;
  wire s_CSAwallace_rca24_and_8_0;
  wire s_CSAwallace_rca24_and_9_0;
  wire s_CSAwallace_rca24_and_10_0;
  wire s_CSAwallace_rca24_and_11_0;
  wire s_CSAwallace_rca24_and_12_0;
  wire s_CSAwallace_rca24_and_13_0;
  wire s_CSAwallace_rca24_and_14_0;
  wire s_CSAwallace_rca24_and_15_0;
  wire s_CSAwallace_rca24_and_16_0;
  wire s_CSAwallace_rca24_and_17_0;
  wire s_CSAwallace_rca24_and_18_0;
  wire s_CSAwallace_rca24_and_19_0;
  wire s_CSAwallace_rca24_and_20_0;
  wire s_CSAwallace_rca24_and_21_0;
  wire s_CSAwallace_rca24_and_22_0;
  wire s_CSAwallace_rca24_nand_23_0;
  wire s_CSAwallace_rca24_and_0_1;
  wire s_CSAwallace_rca24_and_1_1;
  wire s_CSAwallace_rca24_and_2_1;
  wire s_CSAwallace_rca24_and_3_1;
  wire s_CSAwallace_rca24_and_4_1;
  wire s_CSAwallace_rca24_and_5_1;
  wire s_CSAwallace_rca24_and_6_1;
  wire s_CSAwallace_rca24_and_7_1;
  wire s_CSAwallace_rca24_and_8_1;
  wire s_CSAwallace_rca24_and_9_1;
  wire s_CSAwallace_rca24_and_10_1;
  wire s_CSAwallace_rca24_and_11_1;
  wire s_CSAwallace_rca24_and_12_1;
  wire s_CSAwallace_rca24_and_13_1;
  wire s_CSAwallace_rca24_and_14_1;
  wire s_CSAwallace_rca24_and_15_1;
  wire s_CSAwallace_rca24_and_16_1;
  wire s_CSAwallace_rca24_and_17_1;
  wire s_CSAwallace_rca24_and_18_1;
  wire s_CSAwallace_rca24_and_19_1;
  wire s_CSAwallace_rca24_and_20_1;
  wire s_CSAwallace_rca24_and_21_1;
  wire s_CSAwallace_rca24_and_22_1;
  wire s_CSAwallace_rca24_nand_23_1;
  wire s_CSAwallace_rca24_and_0_2;
  wire s_CSAwallace_rca24_and_1_2;
  wire s_CSAwallace_rca24_and_2_2;
  wire s_CSAwallace_rca24_and_3_2;
  wire s_CSAwallace_rca24_and_4_2;
  wire s_CSAwallace_rca24_and_5_2;
  wire s_CSAwallace_rca24_and_6_2;
  wire s_CSAwallace_rca24_and_7_2;
  wire s_CSAwallace_rca24_and_8_2;
  wire s_CSAwallace_rca24_and_9_2;
  wire s_CSAwallace_rca24_and_10_2;
  wire s_CSAwallace_rca24_and_11_2;
  wire s_CSAwallace_rca24_and_12_2;
  wire s_CSAwallace_rca24_and_13_2;
  wire s_CSAwallace_rca24_and_14_2;
  wire s_CSAwallace_rca24_and_15_2;
  wire s_CSAwallace_rca24_and_16_2;
  wire s_CSAwallace_rca24_and_17_2;
  wire s_CSAwallace_rca24_and_18_2;
  wire s_CSAwallace_rca24_and_19_2;
  wire s_CSAwallace_rca24_and_20_2;
  wire s_CSAwallace_rca24_and_21_2;
  wire s_CSAwallace_rca24_and_22_2;
  wire s_CSAwallace_rca24_nand_23_2;
  wire s_CSAwallace_rca24_and_0_3;
  wire s_CSAwallace_rca24_and_1_3;
  wire s_CSAwallace_rca24_and_2_3;
  wire s_CSAwallace_rca24_and_3_3;
  wire s_CSAwallace_rca24_and_4_3;
  wire s_CSAwallace_rca24_and_5_3;
  wire s_CSAwallace_rca24_and_6_3;
  wire s_CSAwallace_rca24_and_7_3;
  wire s_CSAwallace_rca24_and_8_3;
  wire s_CSAwallace_rca24_and_9_3;
  wire s_CSAwallace_rca24_and_10_3;
  wire s_CSAwallace_rca24_and_11_3;
  wire s_CSAwallace_rca24_and_12_3;
  wire s_CSAwallace_rca24_and_13_3;
  wire s_CSAwallace_rca24_and_14_3;
  wire s_CSAwallace_rca24_and_15_3;
  wire s_CSAwallace_rca24_and_16_3;
  wire s_CSAwallace_rca24_and_17_3;
  wire s_CSAwallace_rca24_and_18_3;
  wire s_CSAwallace_rca24_and_19_3;
  wire s_CSAwallace_rca24_and_20_3;
  wire s_CSAwallace_rca24_and_21_3;
  wire s_CSAwallace_rca24_and_22_3;
  wire s_CSAwallace_rca24_nand_23_3;
  wire s_CSAwallace_rca24_and_0_4;
  wire s_CSAwallace_rca24_and_1_4;
  wire s_CSAwallace_rca24_and_2_4;
  wire s_CSAwallace_rca24_and_3_4;
  wire s_CSAwallace_rca24_and_4_4;
  wire s_CSAwallace_rca24_and_5_4;
  wire s_CSAwallace_rca24_and_6_4;
  wire s_CSAwallace_rca24_and_7_4;
  wire s_CSAwallace_rca24_and_8_4;
  wire s_CSAwallace_rca24_and_9_4;
  wire s_CSAwallace_rca24_and_10_4;
  wire s_CSAwallace_rca24_and_11_4;
  wire s_CSAwallace_rca24_and_12_4;
  wire s_CSAwallace_rca24_and_13_4;
  wire s_CSAwallace_rca24_and_14_4;
  wire s_CSAwallace_rca24_and_15_4;
  wire s_CSAwallace_rca24_and_16_4;
  wire s_CSAwallace_rca24_and_17_4;
  wire s_CSAwallace_rca24_and_18_4;
  wire s_CSAwallace_rca24_and_19_4;
  wire s_CSAwallace_rca24_and_20_4;
  wire s_CSAwallace_rca24_and_21_4;
  wire s_CSAwallace_rca24_and_22_4;
  wire s_CSAwallace_rca24_nand_23_4;
  wire s_CSAwallace_rca24_and_0_5;
  wire s_CSAwallace_rca24_and_1_5;
  wire s_CSAwallace_rca24_and_2_5;
  wire s_CSAwallace_rca24_and_3_5;
  wire s_CSAwallace_rca24_and_4_5;
  wire s_CSAwallace_rca24_and_5_5;
  wire s_CSAwallace_rca24_and_6_5;
  wire s_CSAwallace_rca24_and_7_5;
  wire s_CSAwallace_rca24_and_8_5;
  wire s_CSAwallace_rca24_and_9_5;
  wire s_CSAwallace_rca24_and_10_5;
  wire s_CSAwallace_rca24_and_11_5;
  wire s_CSAwallace_rca24_and_12_5;
  wire s_CSAwallace_rca24_and_13_5;
  wire s_CSAwallace_rca24_and_14_5;
  wire s_CSAwallace_rca24_and_15_5;
  wire s_CSAwallace_rca24_and_16_5;
  wire s_CSAwallace_rca24_and_17_5;
  wire s_CSAwallace_rca24_and_18_5;
  wire s_CSAwallace_rca24_and_19_5;
  wire s_CSAwallace_rca24_and_20_5;
  wire s_CSAwallace_rca24_and_21_5;
  wire s_CSAwallace_rca24_and_22_5;
  wire s_CSAwallace_rca24_nand_23_5;
  wire s_CSAwallace_rca24_and_0_6;
  wire s_CSAwallace_rca24_and_1_6;
  wire s_CSAwallace_rca24_and_2_6;
  wire s_CSAwallace_rca24_and_3_6;
  wire s_CSAwallace_rca24_and_4_6;
  wire s_CSAwallace_rca24_and_5_6;
  wire s_CSAwallace_rca24_and_6_6;
  wire s_CSAwallace_rca24_and_7_6;
  wire s_CSAwallace_rca24_and_8_6;
  wire s_CSAwallace_rca24_and_9_6;
  wire s_CSAwallace_rca24_and_10_6;
  wire s_CSAwallace_rca24_and_11_6;
  wire s_CSAwallace_rca24_and_12_6;
  wire s_CSAwallace_rca24_and_13_6;
  wire s_CSAwallace_rca24_and_14_6;
  wire s_CSAwallace_rca24_and_15_6;
  wire s_CSAwallace_rca24_and_16_6;
  wire s_CSAwallace_rca24_and_17_6;
  wire s_CSAwallace_rca24_and_18_6;
  wire s_CSAwallace_rca24_and_19_6;
  wire s_CSAwallace_rca24_and_20_6;
  wire s_CSAwallace_rca24_and_21_6;
  wire s_CSAwallace_rca24_and_22_6;
  wire s_CSAwallace_rca24_nand_23_6;
  wire s_CSAwallace_rca24_and_0_7;
  wire s_CSAwallace_rca24_and_1_7;
  wire s_CSAwallace_rca24_and_2_7;
  wire s_CSAwallace_rca24_and_3_7;
  wire s_CSAwallace_rca24_and_4_7;
  wire s_CSAwallace_rca24_and_5_7;
  wire s_CSAwallace_rca24_and_6_7;
  wire s_CSAwallace_rca24_and_7_7;
  wire s_CSAwallace_rca24_and_8_7;
  wire s_CSAwallace_rca24_and_9_7;
  wire s_CSAwallace_rca24_and_10_7;
  wire s_CSAwallace_rca24_and_11_7;
  wire s_CSAwallace_rca24_and_12_7;
  wire s_CSAwallace_rca24_and_13_7;
  wire s_CSAwallace_rca24_and_14_7;
  wire s_CSAwallace_rca24_and_15_7;
  wire s_CSAwallace_rca24_and_16_7;
  wire s_CSAwallace_rca24_and_17_7;
  wire s_CSAwallace_rca24_and_18_7;
  wire s_CSAwallace_rca24_and_19_7;
  wire s_CSAwallace_rca24_and_20_7;
  wire s_CSAwallace_rca24_and_21_7;
  wire s_CSAwallace_rca24_and_22_7;
  wire s_CSAwallace_rca24_nand_23_7;
  wire s_CSAwallace_rca24_and_0_8;
  wire s_CSAwallace_rca24_and_1_8;
  wire s_CSAwallace_rca24_and_2_8;
  wire s_CSAwallace_rca24_and_3_8;
  wire s_CSAwallace_rca24_and_4_8;
  wire s_CSAwallace_rca24_and_5_8;
  wire s_CSAwallace_rca24_and_6_8;
  wire s_CSAwallace_rca24_and_7_8;
  wire s_CSAwallace_rca24_and_8_8;
  wire s_CSAwallace_rca24_and_9_8;
  wire s_CSAwallace_rca24_and_10_8;
  wire s_CSAwallace_rca24_and_11_8;
  wire s_CSAwallace_rca24_and_12_8;
  wire s_CSAwallace_rca24_and_13_8;
  wire s_CSAwallace_rca24_and_14_8;
  wire s_CSAwallace_rca24_and_15_8;
  wire s_CSAwallace_rca24_and_16_8;
  wire s_CSAwallace_rca24_and_17_8;
  wire s_CSAwallace_rca24_and_18_8;
  wire s_CSAwallace_rca24_and_19_8;
  wire s_CSAwallace_rca24_and_20_8;
  wire s_CSAwallace_rca24_and_21_8;
  wire s_CSAwallace_rca24_and_22_8;
  wire s_CSAwallace_rca24_nand_23_8;
  wire s_CSAwallace_rca24_and_0_9;
  wire s_CSAwallace_rca24_and_1_9;
  wire s_CSAwallace_rca24_and_2_9;
  wire s_CSAwallace_rca24_and_3_9;
  wire s_CSAwallace_rca24_and_4_9;
  wire s_CSAwallace_rca24_and_5_9;
  wire s_CSAwallace_rca24_and_6_9;
  wire s_CSAwallace_rca24_and_7_9;
  wire s_CSAwallace_rca24_and_8_9;
  wire s_CSAwallace_rca24_and_9_9;
  wire s_CSAwallace_rca24_and_10_9;
  wire s_CSAwallace_rca24_and_11_9;
  wire s_CSAwallace_rca24_and_12_9;
  wire s_CSAwallace_rca24_and_13_9;
  wire s_CSAwallace_rca24_and_14_9;
  wire s_CSAwallace_rca24_and_15_9;
  wire s_CSAwallace_rca24_and_16_9;
  wire s_CSAwallace_rca24_and_17_9;
  wire s_CSAwallace_rca24_and_18_9;
  wire s_CSAwallace_rca24_and_19_9;
  wire s_CSAwallace_rca24_and_20_9;
  wire s_CSAwallace_rca24_and_21_9;
  wire s_CSAwallace_rca24_and_22_9;
  wire s_CSAwallace_rca24_nand_23_9;
  wire s_CSAwallace_rca24_and_0_10;
  wire s_CSAwallace_rca24_and_1_10;
  wire s_CSAwallace_rca24_and_2_10;
  wire s_CSAwallace_rca24_and_3_10;
  wire s_CSAwallace_rca24_and_4_10;
  wire s_CSAwallace_rca24_and_5_10;
  wire s_CSAwallace_rca24_and_6_10;
  wire s_CSAwallace_rca24_and_7_10;
  wire s_CSAwallace_rca24_and_8_10;
  wire s_CSAwallace_rca24_and_9_10;
  wire s_CSAwallace_rca24_and_10_10;
  wire s_CSAwallace_rca24_and_11_10;
  wire s_CSAwallace_rca24_and_12_10;
  wire s_CSAwallace_rca24_and_13_10;
  wire s_CSAwallace_rca24_and_14_10;
  wire s_CSAwallace_rca24_and_15_10;
  wire s_CSAwallace_rca24_and_16_10;
  wire s_CSAwallace_rca24_and_17_10;
  wire s_CSAwallace_rca24_and_18_10;
  wire s_CSAwallace_rca24_and_19_10;
  wire s_CSAwallace_rca24_and_20_10;
  wire s_CSAwallace_rca24_and_21_10;
  wire s_CSAwallace_rca24_and_22_10;
  wire s_CSAwallace_rca24_nand_23_10;
  wire s_CSAwallace_rca24_and_0_11;
  wire s_CSAwallace_rca24_and_1_11;
  wire s_CSAwallace_rca24_and_2_11;
  wire s_CSAwallace_rca24_and_3_11;
  wire s_CSAwallace_rca24_and_4_11;
  wire s_CSAwallace_rca24_and_5_11;
  wire s_CSAwallace_rca24_and_6_11;
  wire s_CSAwallace_rca24_and_7_11;
  wire s_CSAwallace_rca24_and_8_11;
  wire s_CSAwallace_rca24_and_9_11;
  wire s_CSAwallace_rca24_and_10_11;
  wire s_CSAwallace_rca24_and_11_11;
  wire s_CSAwallace_rca24_and_12_11;
  wire s_CSAwallace_rca24_and_13_11;
  wire s_CSAwallace_rca24_and_14_11;
  wire s_CSAwallace_rca24_and_15_11;
  wire s_CSAwallace_rca24_and_16_11;
  wire s_CSAwallace_rca24_and_17_11;
  wire s_CSAwallace_rca24_and_18_11;
  wire s_CSAwallace_rca24_and_19_11;
  wire s_CSAwallace_rca24_and_20_11;
  wire s_CSAwallace_rca24_and_21_11;
  wire s_CSAwallace_rca24_and_22_11;
  wire s_CSAwallace_rca24_nand_23_11;
  wire s_CSAwallace_rca24_and_0_12;
  wire s_CSAwallace_rca24_and_1_12;
  wire s_CSAwallace_rca24_and_2_12;
  wire s_CSAwallace_rca24_and_3_12;
  wire s_CSAwallace_rca24_and_4_12;
  wire s_CSAwallace_rca24_and_5_12;
  wire s_CSAwallace_rca24_and_6_12;
  wire s_CSAwallace_rca24_and_7_12;
  wire s_CSAwallace_rca24_and_8_12;
  wire s_CSAwallace_rca24_and_9_12;
  wire s_CSAwallace_rca24_and_10_12;
  wire s_CSAwallace_rca24_and_11_12;
  wire s_CSAwallace_rca24_and_12_12;
  wire s_CSAwallace_rca24_and_13_12;
  wire s_CSAwallace_rca24_and_14_12;
  wire s_CSAwallace_rca24_and_15_12;
  wire s_CSAwallace_rca24_and_16_12;
  wire s_CSAwallace_rca24_and_17_12;
  wire s_CSAwallace_rca24_and_18_12;
  wire s_CSAwallace_rca24_and_19_12;
  wire s_CSAwallace_rca24_and_20_12;
  wire s_CSAwallace_rca24_and_21_12;
  wire s_CSAwallace_rca24_and_22_12;
  wire s_CSAwallace_rca24_nand_23_12;
  wire s_CSAwallace_rca24_and_0_13;
  wire s_CSAwallace_rca24_and_1_13;
  wire s_CSAwallace_rca24_and_2_13;
  wire s_CSAwallace_rca24_and_3_13;
  wire s_CSAwallace_rca24_and_4_13;
  wire s_CSAwallace_rca24_and_5_13;
  wire s_CSAwallace_rca24_and_6_13;
  wire s_CSAwallace_rca24_and_7_13;
  wire s_CSAwallace_rca24_and_8_13;
  wire s_CSAwallace_rca24_and_9_13;
  wire s_CSAwallace_rca24_and_10_13;
  wire s_CSAwallace_rca24_and_11_13;
  wire s_CSAwallace_rca24_and_12_13;
  wire s_CSAwallace_rca24_and_13_13;
  wire s_CSAwallace_rca24_and_14_13;
  wire s_CSAwallace_rca24_and_15_13;
  wire s_CSAwallace_rca24_and_16_13;
  wire s_CSAwallace_rca24_and_17_13;
  wire s_CSAwallace_rca24_and_18_13;
  wire s_CSAwallace_rca24_and_19_13;
  wire s_CSAwallace_rca24_and_20_13;
  wire s_CSAwallace_rca24_and_21_13;
  wire s_CSAwallace_rca24_and_22_13;
  wire s_CSAwallace_rca24_nand_23_13;
  wire s_CSAwallace_rca24_and_0_14;
  wire s_CSAwallace_rca24_and_1_14;
  wire s_CSAwallace_rca24_and_2_14;
  wire s_CSAwallace_rca24_and_3_14;
  wire s_CSAwallace_rca24_and_4_14;
  wire s_CSAwallace_rca24_and_5_14;
  wire s_CSAwallace_rca24_and_6_14;
  wire s_CSAwallace_rca24_and_7_14;
  wire s_CSAwallace_rca24_and_8_14;
  wire s_CSAwallace_rca24_and_9_14;
  wire s_CSAwallace_rca24_and_10_14;
  wire s_CSAwallace_rca24_and_11_14;
  wire s_CSAwallace_rca24_and_12_14;
  wire s_CSAwallace_rca24_and_13_14;
  wire s_CSAwallace_rca24_and_14_14;
  wire s_CSAwallace_rca24_and_15_14;
  wire s_CSAwallace_rca24_and_16_14;
  wire s_CSAwallace_rca24_and_17_14;
  wire s_CSAwallace_rca24_and_18_14;
  wire s_CSAwallace_rca24_and_19_14;
  wire s_CSAwallace_rca24_and_20_14;
  wire s_CSAwallace_rca24_and_21_14;
  wire s_CSAwallace_rca24_and_22_14;
  wire s_CSAwallace_rca24_nand_23_14;
  wire s_CSAwallace_rca24_and_0_15;
  wire s_CSAwallace_rca24_and_1_15;
  wire s_CSAwallace_rca24_and_2_15;
  wire s_CSAwallace_rca24_and_3_15;
  wire s_CSAwallace_rca24_and_4_15;
  wire s_CSAwallace_rca24_and_5_15;
  wire s_CSAwallace_rca24_and_6_15;
  wire s_CSAwallace_rca24_and_7_15;
  wire s_CSAwallace_rca24_and_8_15;
  wire s_CSAwallace_rca24_and_9_15;
  wire s_CSAwallace_rca24_and_10_15;
  wire s_CSAwallace_rca24_and_11_15;
  wire s_CSAwallace_rca24_and_12_15;
  wire s_CSAwallace_rca24_and_13_15;
  wire s_CSAwallace_rca24_and_14_15;
  wire s_CSAwallace_rca24_and_15_15;
  wire s_CSAwallace_rca24_and_16_15;
  wire s_CSAwallace_rca24_and_17_15;
  wire s_CSAwallace_rca24_and_18_15;
  wire s_CSAwallace_rca24_and_19_15;
  wire s_CSAwallace_rca24_and_20_15;
  wire s_CSAwallace_rca24_and_21_15;
  wire s_CSAwallace_rca24_and_22_15;
  wire s_CSAwallace_rca24_nand_23_15;
  wire s_CSAwallace_rca24_and_0_16;
  wire s_CSAwallace_rca24_and_1_16;
  wire s_CSAwallace_rca24_and_2_16;
  wire s_CSAwallace_rca24_and_3_16;
  wire s_CSAwallace_rca24_and_4_16;
  wire s_CSAwallace_rca24_and_5_16;
  wire s_CSAwallace_rca24_and_6_16;
  wire s_CSAwallace_rca24_and_7_16;
  wire s_CSAwallace_rca24_and_8_16;
  wire s_CSAwallace_rca24_and_9_16;
  wire s_CSAwallace_rca24_and_10_16;
  wire s_CSAwallace_rca24_and_11_16;
  wire s_CSAwallace_rca24_and_12_16;
  wire s_CSAwallace_rca24_and_13_16;
  wire s_CSAwallace_rca24_and_14_16;
  wire s_CSAwallace_rca24_and_15_16;
  wire s_CSAwallace_rca24_and_16_16;
  wire s_CSAwallace_rca24_and_17_16;
  wire s_CSAwallace_rca24_and_18_16;
  wire s_CSAwallace_rca24_and_19_16;
  wire s_CSAwallace_rca24_and_20_16;
  wire s_CSAwallace_rca24_and_21_16;
  wire s_CSAwallace_rca24_and_22_16;
  wire s_CSAwallace_rca24_nand_23_16;
  wire s_CSAwallace_rca24_and_0_17;
  wire s_CSAwallace_rca24_and_1_17;
  wire s_CSAwallace_rca24_and_2_17;
  wire s_CSAwallace_rca24_and_3_17;
  wire s_CSAwallace_rca24_and_4_17;
  wire s_CSAwallace_rca24_and_5_17;
  wire s_CSAwallace_rca24_and_6_17;
  wire s_CSAwallace_rca24_and_7_17;
  wire s_CSAwallace_rca24_and_8_17;
  wire s_CSAwallace_rca24_and_9_17;
  wire s_CSAwallace_rca24_and_10_17;
  wire s_CSAwallace_rca24_and_11_17;
  wire s_CSAwallace_rca24_and_12_17;
  wire s_CSAwallace_rca24_and_13_17;
  wire s_CSAwallace_rca24_and_14_17;
  wire s_CSAwallace_rca24_and_15_17;
  wire s_CSAwallace_rca24_and_16_17;
  wire s_CSAwallace_rca24_and_17_17;
  wire s_CSAwallace_rca24_and_18_17;
  wire s_CSAwallace_rca24_and_19_17;
  wire s_CSAwallace_rca24_and_20_17;
  wire s_CSAwallace_rca24_and_21_17;
  wire s_CSAwallace_rca24_and_22_17;
  wire s_CSAwallace_rca24_nand_23_17;
  wire s_CSAwallace_rca24_and_0_18;
  wire s_CSAwallace_rca24_and_1_18;
  wire s_CSAwallace_rca24_and_2_18;
  wire s_CSAwallace_rca24_and_3_18;
  wire s_CSAwallace_rca24_and_4_18;
  wire s_CSAwallace_rca24_and_5_18;
  wire s_CSAwallace_rca24_and_6_18;
  wire s_CSAwallace_rca24_and_7_18;
  wire s_CSAwallace_rca24_and_8_18;
  wire s_CSAwallace_rca24_and_9_18;
  wire s_CSAwallace_rca24_and_10_18;
  wire s_CSAwallace_rca24_and_11_18;
  wire s_CSAwallace_rca24_and_12_18;
  wire s_CSAwallace_rca24_and_13_18;
  wire s_CSAwallace_rca24_and_14_18;
  wire s_CSAwallace_rca24_and_15_18;
  wire s_CSAwallace_rca24_and_16_18;
  wire s_CSAwallace_rca24_and_17_18;
  wire s_CSAwallace_rca24_and_18_18;
  wire s_CSAwallace_rca24_and_19_18;
  wire s_CSAwallace_rca24_and_20_18;
  wire s_CSAwallace_rca24_and_21_18;
  wire s_CSAwallace_rca24_and_22_18;
  wire s_CSAwallace_rca24_nand_23_18;
  wire s_CSAwallace_rca24_and_0_19;
  wire s_CSAwallace_rca24_and_1_19;
  wire s_CSAwallace_rca24_and_2_19;
  wire s_CSAwallace_rca24_and_3_19;
  wire s_CSAwallace_rca24_and_4_19;
  wire s_CSAwallace_rca24_and_5_19;
  wire s_CSAwallace_rca24_and_6_19;
  wire s_CSAwallace_rca24_and_7_19;
  wire s_CSAwallace_rca24_and_8_19;
  wire s_CSAwallace_rca24_and_9_19;
  wire s_CSAwallace_rca24_and_10_19;
  wire s_CSAwallace_rca24_and_11_19;
  wire s_CSAwallace_rca24_and_12_19;
  wire s_CSAwallace_rca24_and_13_19;
  wire s_CSAwallace_rca24_and_14_19;
  wire s_CSAwallace_rca24_and_15_19;
  wire s_CSAwallace_rca24_and_16_19;
  wire s_CSAwallace_rca24_and_17_19;
  wire s_CSAwallace_rca24_and_18_19;
  wire s_CSAwallace_rca24_and_19_19;
  wire s_CSAwallace_rca24_and_20_19;
  wire s_CSAwallace_rca24_and_21_19;
  wire s_CSAwallace_rca24_and_22_19;
  wire s_CSAwallace_rca24_nand_23_19;
  wire s_CSAwallace_rca24_and_0_20;
  wire s_CSAwallace_rca24_and_1_20;
  wire s_CSAwallace_rca24_and_2_20;
  wire s_CSAwallace_rca24_and_3_20;
  wire s_CSAwallace_rca24_and_4_20;
  wire s_CSAwallace_rca24_and_5_20;
  wire s_CSAwallace_rca24_and_6_20;
  wire s_CSAwallace_rca24_and_7_20;
  wire s_CSAwallace_rca24_and_8_20;
  wire s_CSAwallace_rca24_and_9_20;
  wire s_CSAwallace_rca24_and_10_20;
  wire s_CSAwallace_rca24_and_11_20;
  wire s_CSAwallace_rca24_and_12_20;
  wire s_CSAwallace_rca24_and_13_20;
  wire s_CSAwallace_rca24_and_14_20;
  wire s_CSAwallace_rca24_and_15_20;
  wire s_CSAwallace_rca24_and_16_20;
  wire s_CSAwallace_rca24_and_17_20;
  wire s_CSAwallace_rca24_and_18_20;
  wire s_CSAwallace_rca24_and_19_20;
  wire s_CSAwallace_rca24_and_20_20;
  wire s_CSAwallace_rca24_and_21_20;
  wire s_CSAwallace_rca24_and_22_20;
  wire s_CSAwallace_rca24_nand_23_20;
  wire s_CSAwallace_rca24_and_0_21;
  wire s_CSAwallace_rca24_and_1_21;
  wire s_CSAwallace_rca24_and_2_21;
  wire s_CSAwallace_rca24_and_3_21;
  wire s_CSAwallace_rca24_and_4_21;
  wire s_CSAwallace_rca24_and_5_21;
  wire s_CSAwallace_rca24_and_6_21;
  wire s_CSAwallace_rca24_and_7_21;
  wire s_CSAwallace_rca24_and_8_21;
  wire s_CSAwallace_rca24_and_9_21;
  wire s_CSAwallace_rca24_and_10_21;
  wire s_CSAwallace_rca24_and_11_21;
  wire s_CSAwallace_rca24_and_12_21;
  wire s_CSAwallace_rca24_and_13_21;
  wire s_CSAwallace_rca24_and_14_21;
  wire s_CSAwallace_rca24_and_15_21;
  wire s_CSAwallace_rca24_and_16_21;
  wire s_CSAwallace_rca24_and_17_21;
  wire s_CSAwallace_rca24_and_18_21;
  wire s_CSAwallace_rca24_and_19_21;
  wire s_CSAwallace_rca24_and_20_21;
  wire s_CSAwallace_rca24_and_21_21;
  wire s_CSAwallace_rca24_and_22_21;
  wire s_CSAwallace_rca24_nand_23_21;
  wire s_CSAwallace_rca24_and_0_22;
  wire s_CSAwallace_rca24_and_1_22;
  wire s_CSAwallace_rca24_and_2_22;
  wire s_CSAwallace_rca24_and_3_22;
  wire s_CSAwallace_rca24_and_4_22;
  wire s_CSAwallace_rca24_and_5_22;
  wire s_CSAwallace_rca24_and_6_22;
  wire s_CSAwallace_rca24_and_7_22;
  wire s_CSAwallace_rca24_and_8_22;
  wire s_CSAwallace_rca24_and_9_22;
  wire s_CSAwallace_rca24_and_10_22;
  wire s_CSAwallace_rca24_and_11_22;
  wire s_CSAwallace_rca24_and_12_22;
  wire s_CSAwallace_rca24_and_13_22;
  wire s_CSAwallace_rca24_and_14_22;
  wire s_CSAwallace_rca24_and_15_22;
  wire s_CSAwallace_rca24_and_16_22;
  wire s_CSAwallace_rca24_and_17_22;
  wire s_CSAwallace_rca24_and_18_22;
  wire s_CSAwallace_rca24_and_19_22;
  wire s_CSAwallace_rca24_and_20_22;
  wire s_CSAwallace_rca24_and_21_22;
  wire s_CSAwallace_rca24_and_22_22;
  wire s_CSAwallace_rca24_nand_23_22;
  wire s_CSAwallace_rca24_nand_0_23;
  wire s_CSAwallace_rca24_nand_1_23;
  wire s_CSAwallace_rca24_nand_2_23;
  wire s_CSAwallace_rca24_nand_3_23;
  wire s_CSAwallace_rca24_nand_4_23;
  wire s_CSAwallace_rca24_nand_5_23;
  wire s_CSAwallace_rca24_nand_6_23;
  wire s_CSAwallace_rca24_nand_7_23;
  wire s_CSAwallace_rca24_nand_8_23;
  wire s_CSAwallace_rca24_nand_9_23;
  wire s_CSAwallace_rca24_nand_10_23;
  wire s_CSAwallace_rca24_nand_11_23;
  wire s_CSAwallace_rca24_nand_12_23;
  wire s_CSAwallace_rca24_nand_13_23;
  wire s_CSAwallace_rca24_nand_14_23;
  wire s_CSAwallace_rca24_nand_15_23;
  wire s_CSAwallace_rca24_nand_16_23;
  wire s_CSAwallace_rca24_nand_17_23;
  wire s_CSAwallace_rca24_nand_18_23;
  wire s_CSAwallace_rca24_nand_19_23;
  wire s_CSAwallace_rca24_nand_20_23;
  wire s_CSAwallace_rca24_nand_21_23;
  wire s_CSAwallace_rca24_nand_22_23;
  wire s_CSAwallace_rca24_and_23_23;
  wire s_CSAwallace_rca24_csa0_csa_component_fa1_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa1_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa2_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa2_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa2_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa2_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa2_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa3_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa3_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa3_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa3_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa3_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa4_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa4_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa4_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa4_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa4_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa5_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa5_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa5_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa5_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa5_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa6_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa6_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa6_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa6_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa6_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa7_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa7_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa7_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa8_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa8_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa8_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa9_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa9_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa9_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa10_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa10_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa10_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa11_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa11_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa11_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa0_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa0_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa4_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa4_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa5_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa5_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa5_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa5_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa5_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa6_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa6_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa6_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa6_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa6_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa7_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa7_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa7_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa8_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa8_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa8_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa9_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa9_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa9_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa10_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa10_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa10_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa11_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa11_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa11_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa1_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa1_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa8_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa8_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa8_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa9_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa9_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa9_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa10_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa10_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa10_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa11_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa11_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa11_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa2_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa2_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa11_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa11_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa11_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa3_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa3_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa4_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa4_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa38_and0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa5_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa5_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa38_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa39_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa40_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa40_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa40_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa40_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa40_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa41_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa41_and0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa41_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa41_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa41_or0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa42_xor0;
  wire s_CSAwallace_rca24_csa6_csa_component_fa42_xor1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa42_and1;
  wire s_CSAwallace_rca24_csa6_csa_component_fa42_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa38_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa39_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa40_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa40_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa40_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa40_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa40_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa41_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa41_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa41_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa41_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa41_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa42_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa42_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa42_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa42_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa42_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa43_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa43_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa43_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa43_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa43_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa44_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa44_and0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa44_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa44_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa44_or0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa45_xor0;
  wire s_CSAwallace_rca24_csa7_csa_component_fa45_xor1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa45_and1;
  wire s_CSAwallace_rca24_csa7_csa_component_fa45_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa2_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa2_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa3_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa3_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa3_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa3_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa3_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa4_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa4_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa4_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa4_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa4_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa5_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa5_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa5_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa5_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa5_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa6_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa6_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa6_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa6_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa6_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa7_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa7_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa7_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa8_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa8_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa8_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa9_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa9_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa9_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa10_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa10_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa10_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa11_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa11_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa11_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa8_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa8_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa6_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa6_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa8_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa8_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa8_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa9_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa9_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa9_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa10_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa10_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa10_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa11_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa11_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa11_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa9_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa9_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa10_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa10_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa40_xor0;
  wire s_CSAwallace_rca24_csa11_csa_component_fa40_xor1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa40_and1;
  wire s_CSAwallace_rca24_csa11_csa_component_fa40_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa38_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa39_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa40_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa40_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa40_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa40_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa40_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa41_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa41_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa41_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa41_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa41_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa42_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa42_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa42_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa42_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa42_or0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa43_xor0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa43_and0;
  wire s_CSAwallace_rca24_csa12_csa_component_fa43_xor1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa43_and1;
  wire s_CSAwallace_rca24_csa12_csa_component_fa43_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa3_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa3_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa4_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa4_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa5_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa5_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa5_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa5_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa5_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa6_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa6_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa6_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa6_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa6_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa7_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa7_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa7_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa8_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa8_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa8_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa9_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa9_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa9_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa10_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa10_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa10_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa11_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa11_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa11_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa13_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa13_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa14_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa14_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa38_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa39_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa40_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa40_and0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa40_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa40_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa40_or0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa41_xor0;
  wire s_CSAwallace_rca24_csa15_csa_component_fa41_xor1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa41_and1;
  wire s_CSAwallace_rca24_csa15_csa_component_fa41_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa4_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa4_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa5_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa5_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa6_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa6_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa7_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa7_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa7_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa8_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa8_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa8_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa9_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa9_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa9_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa10_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa10_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa10_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa11_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa11_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa11_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa16_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa16_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa38_and0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa40_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa40_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa40_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa40_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa41_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa41_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa41_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa41_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa42_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa42_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa42_and1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa42_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa43_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa43_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa43_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa44_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa44_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa44_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa45_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa45_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa45_or0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa46_xor0;
  wire s_CSAwallace_rca24_csa17_csa_component_fa46_xor1;
  wire s_CSAwallace_rca24_csa17_csa_component_fa46_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa5_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa5_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa6_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa6_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa10_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa10_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa10_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa11_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa11_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa11_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa12_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa12_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa12_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa13_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa13_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa13_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa14_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa14_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa14_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa18_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa18_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa38_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa39_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa40_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa40_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa40_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa40_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa40_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa41_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa41_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa41_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa41_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa41_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa42_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa42_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa42_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa42_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa42_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa43_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa43_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa43_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa43_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa43_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa44_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa44_and0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa44_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa44_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa44_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa45_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa45_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa45_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa45_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa46_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa46_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa46_and1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa46_or0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa47_xor0;
  wire s_CSAwallace_rca24_csa19_csa_component_fa47_xor1;
  wire s_CSAwallace_rca24_csa19_csa_component_fa47_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa6_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa6_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa15_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa15_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa15_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa16_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa16_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa16_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa17_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa17_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa17_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa18_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa18_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa18_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa19_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa19_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa19_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa20_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa20_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa20_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa21_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa21_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa21_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa38_and0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa40_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa40_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa40_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa40_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa41_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa41_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa41_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa41_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa42_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa42_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa42_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa42_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa43_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa43_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa43_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa43_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa44_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa44_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa44_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa44_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa45_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa45_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa45_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa45_or0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa46_xor0;
  wire s_CSAwallace_rca24_csa20_csa_component_fa46_xor1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa46_and1;
  wire s_CSAwallace_rca24_csa20_csa_component_fa46_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa7_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa7_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa8_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa8_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa9_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa9_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa10_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa10_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa11_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa11_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa12_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa12_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa13_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa13_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa14_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa14_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa15_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa15_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa16_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa16_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa17_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa17_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa18_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa18_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa19_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa19_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa20_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa20_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa21_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa21_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa22_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa22_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa22_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa22_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa22_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa23_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa23_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa23_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa23_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa23_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa24_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa24_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa24_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa24_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa24_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa25_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa25_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa25_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa25_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa25_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa26_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa26_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa26_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa26_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa26_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa27_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa27_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa27_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa27_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa27_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa28_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa28_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa28_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa28_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa28_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa29_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa29_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa29_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa29_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa29_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa30_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa30_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa30_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa30_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa30_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa31_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa31_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa31_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa31_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa31_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa32_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa32_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa32_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa32_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa32_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa33_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa33_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa33_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa33_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa33_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa34_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa34_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa34_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa34_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa34_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa35_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa35_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa35_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa35_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa35_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa36_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa36_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa36_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa36_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa36_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa37_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa37_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa37_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa37_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa37_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa38_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa38_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa38_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa38_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa38_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa39_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa39_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa39_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa39_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa39_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa40_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa40_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa40_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa40_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa40_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa41_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa41_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa41_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa41_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa41_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa42_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa42_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa42_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa42_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa42_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa43_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa43_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa43_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa43_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa43_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa44_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa44_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa44_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa44_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa44_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa45_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa45_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa45_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa45_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa45_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa46_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa46_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa46_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa46_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa46_or0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa47_xor0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa47_and0;
  wire s_CSAwallace_rca24_csa21_csa_component_fa47_xor1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa47_and1;
  wire s_CSAwallace_rca24_csa21_csa_component_fa47_or0;
  wire s_CSAwallace_rca24_u_rca48_fa8_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa8_and0;
  wire s_CSAwallace_rca24_u_rca48_fa9_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa9_and0;
  wire s_CSAwallace_rca24_u_rca48_fa9_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa9_and1;
  wire s_CSAwallace_rca24_u_rca48_fa9_or0;
  wire s_CSAwallace_rca24_u_rca48_fa10_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa10_and0;
  wire s_CSAwallace_rca24_u_rca48_fa10_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa10_and1;
  wire s_CSAwallace_rca24_u_rca48_fa10_or0;
  wire s_CSAwallace_rca24_u_rca48_fa11_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa11_and0;
  wire s_CSAwallace_rca24_u_rca48_fa11_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa11_and1;
  wire s_CSAwallace_rca24_u_rca48_fa11_or0;
  wire s_CSAwallace_rca24_u_rca48_fa12_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa12_and0;
  wire s_CSAwallace_rca24_u_rca48_fa12_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa12_and1;
  wire s_CSAwallace_rca24_u_rca48_fa12_or0;
  wire s_CSAwallace_rca24_u_rca48_fa13_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa13_and0;
  wire s_CSAwallace_rca24_u_rca48_fa13_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa13_and1;
  wire s_CSAwallace_rca24_u_rca48_fa13_or0;
  wire s_CSAwallace_rca24_u_rca48_fa14_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa14_and0;
  wire s_CSAwallace_rca24_u_rca48_fa14_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa14_and1;
  wire s_CSAwallace_rca24_u_rca48_fa14_or0;
  wire s_CSAwallace_rca24_u_rca48_fa15_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa15_and0;
  wire s_CSAwallace_rca24_u_rca48_fa15_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa15_and1;
  wire s_CSAwallace_rca24_u_rca48_fa15_or0;
  wire s_CSAwallace_rca24_u_rca48_fa16_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa16_and0;
  wire s_CSAwallace_rca24_u_rca48_fa16_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa16_and1;
  wire s_CSAwallace_rca24_u_rca48_fa16_or0;
  wire s_CSAwallace_rca24_u_rca48_fa17_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa17_and0;
  wire s_CSAwallace_rca24_u_rca48_fa17_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa17_and1;
  wire s_CSAwallace_rca24_u_rca48_fa17_or0;
  wire s_CSAwallace_rca24_u_rca48_fa18_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa18_and0;
  wire s_CSAwallace_rca24_u_rca48_fa18_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa18_and1;
  wire s_CSAwallace_rca24_u_rca48_fa18_or0;
  wire s_CSAwallace_rca24_u_rca48_fa19_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa19_and0;
  wire s_CSAwallace_rca24_u_rca48_fa19_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa19_and1;
  wire s_CSAwallace_rca24_u_rca48_fa19_or0;
  wire s_CSAwallace_rca24_u_rca48_fa20_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa20_and0;
  wire s_CSAwallace_rca24_u_rca48_fa20_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa20_and1;
  wire s_CSAwallace_rca24_u_rca48_fa20_or0;
  wire s_CSAwallace_rca24_u_rca48_fa21_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa21_and0;
  wire s_CSAwallace_rca24_u_rca48_fa21_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa21_and1;
  wire s_CSAwallace_rca24_u_rca48_fa21_or0;
  wire s_CSAwallace_rca24_u_rca48_fa22_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa22_and0;
  wire s_CSAwallace_rca24_u_rca48_fa22_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa22_and1;
  wire s_CSAwallace_rca24_u_rca48_fa22_or0;
  wire s_CSAwallace_rca24_u_rca48_fa23_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa23_and0;
  wire s_CSAwallace_rca24_u_rca48_fa23_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa23_and1;
  wire s_CSAwallace_rca24_u_rca48_fa23_or0;
  wire s_CSAwallace_rca24_u_rca48_fa24_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa24_and0;
  wire s_CSAwallace_rca24_u_rca48_fa24_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa24_and1;
  wire s_CSAwallace_rca24_u_rca48_fa24_or0;
  wire s_CSAwallace_rca24_u_rca48_fa25_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa25_and0;
  wire s_CSAwallace_rca24_u_rca48_fa25_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa25_and1;
  wire s_CSAwallace_rca24_u_rca48_fa25_or0;
  wire s_CSAwallace_rca24_u_rca48_fa26_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa26_and0;
  wire s_CSAwallace_rca24_u_rca48_fa26_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa26_and1;
  wire s_CSAwallace_rca24_u_rca48_fa26_or0;
  wire s_CSAwallace_rca24_u_rca48_fa27_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa27_and0;
  wire s_CSAwallace_rca24_u_rca48_fa27_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa27_and1;
  wire s_CSAwallace_rca24_u_rca48_fa27_or0;
  wire s_CSAwallace_rca24_u_rca48_fa28_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa28_and0;
  wire s_CSAwallace_rca24_u_rca48_fa28_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa28_and1;
  wire s_CSAwallace_rca24_u_rca48_fa28_or0;
  wire s_CSAwallace_rca24_u_rca48_fa29_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa29_and0;
  wire s_CSAwallace_rca24_u_rca48_fa29_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa29_and1;
  wire s_CSAwallace_rca24_u_rca48_fa29_or0;
  wire s_CSAwallace_rca24_u_rca48_fa30_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa30_and0;
  wire s_CSAwallace_rca24_u_rca48_fa30_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa30_and1;
  wire s_CSAwallace_rca24_u_rca48_fa30_or0;
  wire s_CSAwallace_rca24_u_rca48_fa31_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa31_and0;
  wire s_CSAwallace_rca24_u_rca48_fa31_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa31_and1;
  wire s_CSAwallace_rca24_u_rca48_fa31_or0;
  wire s_CSAwallace_rca24_u_rca48_fa32_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa32_and0;
  wire s_CSAwallace_rca24_u_rca48_fa32_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa32_and1;
  wire s_CSAwallace_rca24_u_rca48_fa32_or0;
  wire s_CSAwallace_rca24_u_rca48_fa33_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa33_and0;
  wire s_CSAwallace_rca24_u_rca48_fa33_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa33_and1;
  wire s_CSAwallace_rca24_u_rca48_fa33_or0;
  wire s_CSAwallace_rca24_u_rca48_fa34_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa34_and0;
  wire s_CSAwallace_rca24_u_rca48_fa34_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa34_and1;
  wire s_CSAwallace_rca24_u_rca48_fa34_or0;
  wire s_CSAwallace_rca24_u_rca48_fa35_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa35_and0;
  wire s_CSAwallace_rca24_u_rca48_fa35_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa35_and1;
  wire s_CSAwallace_rca24_u_rca48_fa35_or0;
  wire s_CSAwallace_rca24_u_rca48_fa36_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa36_and0;
  wire s_CSAwallace_rca24_u_rca48_fa36_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa36_and1;
  wire s_CSAwallace_rca24_u_rca48_fa36_or0;
  wire s_CSAwallace_rca24_u_rca48_fa37_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa37_and0;
  wire s_CSAwallace_rca24_u_rca48_fa37_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa37_and1;
  wire s_CSAwallace_rca24_u_rca48_fa37_or0;
  wire s_CSAwallace_rca24_u_rca48_fa38_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa38_and0;
  wire s_CSAwallace_rca24_u_rca48_fa38_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa38_and1;
  wire s_CSAwallace_rca24_u_rca48_fa38_or0;
  wire s_CSAwallace_rca24_u_rca48_fa39_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa39_and0;
  wire s_CSAwallace_rca24_u_rca48_fa39_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa39_and1;
  wire s_CSAwallace_rca24_u_rca48_fa39_or0;
  wire s_CSAwallace_rca24_u_rca48_fa40_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa40_and0;
  wire s_CSAwallace_rca24_u_rca48_fa40_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa40_and1;
  wire s_CSAwallace_rca24_u_rca48_fa40_or0;
  wire s_CSAwallace_rca24_u_rca48_fa41_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa41_and0;
  wire s_CSAwallace_rca24_u_rca48_fa41_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa41_and1;
  wire s_CSAwallace_rca24_u_rca48_fa41_or0;
  wire s_CSAwallace_rca24_u_rca48_fa42_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa42_and0;
  wire s_CSAwallace_rca24_u_rca48_fa42_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa42_and1;
  wire s_CSAwallace_rca24_u_rca48_fa42_or0;
  wire s_CSAwallace_rca24_u_rca48_fa43_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa43_and0;
  wire s_CSAwallace_rca24_u_rca48_fa43_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa43_and1;
  wire s_CSAwallace_rca24_u_rca48_fa43_or0;
  wire s_CSAwallace_rca24_u_rca48_fa44_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa44_and0;
  wire s_CSAwallace_rca24_u_rca48_fa44_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa44_and1;
  wire s_CSAwallace_rca24_u_rca48_fa44_or0;
  wire s_CSAwallace_rca24_u_rca48_fa45_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa45_and0;
  wire s_CSAwallace_rca24_u_rca48_fa45_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa45_and1;
  wire s_CSAwallace_rca24_u_rca48_fa45_or0;
  wire s_CSAwallace_rca24_u_rca48_fa46_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa46_and0;
  wire s_CSAwallace_rca24_u_rca48_fa46_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa46_and1;
  wire s_CSAwallace_rca24_u_rca48_fa46_or0;
  wire s_CSAwallace_rca24_u_rca48_fa47_xor0;
  wire s_CSAwallace_rca24_u_rca48_fa47_and0;
  wire s_CSAwallace_rca24_u_rca48_fa47_xor1;
  wire s_CSAwallace_rca24_u_rca48_fa47_and1;
  wire s_CSAwallace_rca24_u_rca48_fa47_or0;
  wire s_CSAwallace_rca24_xor0;

  assign s_CSAwallace_rca24_and_0_0 = a[0] & b[0];
  assign s_CSAwallace_rca24_and_1_0 = a[1] & b[0];
  assign s_CSAwallace_rca24_and_2_0 = a[2] & b[0];
  assign s_CSAwallace_rca24_and_3_0 = a[3] & b[0];
  assign s_CSAwallace_rca24_and_4_0 = a[4] & b[0];
  assign s_CSAwallace_rca24_and_5_0 = a[5] & b[0];
  assign s_CSAwallace_rca24_and_6_0 = a[6] & b[0];
  assign s_CSAwallace_rca24_and_7_0 = a[7] & b[0];
  assign s_CSAwallace_rca24_and_8_0 = a[8] & b[0];
  assign s_CSAwallace_rca24_and_9_0 = a[9] & b[0];
  assign s_CSAwallace_rca24_and_10_0 = a[10] & b[0];
  assign s_CSAwallace_rca24_and_11_0 = a[11] & b[0];
  assign s_CSAwallace_rca24_and_12_0 = a[12] & b[0];
  assign s_CSAwallace_rca24_and_13_0 = a[13] & b[0];
  assign s_CSAwallace_rca24_and_14_0 = a[14] & b[0];
  assign s_CSAwallace_rca24_and_15_0 = a[15] & b[0];
  assign s_CSAwallace_rca24_and_16_0 = a[16] & b[0];
  assign s_CSAwallace_rca24_and_17_0 = a[17] & b[0];
  assign s_CSAwallace_rca24_and_18_0 = a[18] & b[0];
  assign s_CSAwallace_rca24_and_19_0 = a[19] & b[0];
  assign s_CSAwallace_rca24_and_20_0 = a[20] & b[0];
  assign s_CSAwallace_rca24_and_21_0 = a[21] & b[0];
  assign s_CSAwallace_rca24_and_22_0 = a[22] & b[0];
  assign s_CSAwallace_rca24_nand_23_0 = ~(a[23] & b[0]);
  assign s_CSAwallace_rca24_and_0_1 = a[0] & b[1];
  assign s_CSAwallace_rca24_and_1_1 = a[1] & b[1];
  assign s_CSAwallace_rca24_and_2_1 = a[2] & b[1];
  assign s_CSAwallace_rca24_and_3_1 = a[3] & b[1];
  assign s_CSAwallace_rca24_and_4_1 = a[4] & b[1];
  assign s_CSAwallace_rca24_and_5_1 = a[5] & b[1];
  assign s_CSAwallace_rca24_and_6_1 = a[6] & b[1];
  assign s_CSAwallace_rca24_and_7_1 = a[7] & b[1];
  assign s_CSAwallace_rca24_and_8_1 = a[8] & b[1];
  assign s_CSAwallace_rca24_and_9_1 = a[9] & b[1];
  assign s_CSAwallace_rca24_and_10_1 = a[10] & b[1];
  assign s_CSAwallace_rca24_and_11_1 = a[11] & b[1];
  assign s_CSAwallace_rca24_and_12_1 = a[12] & b[1];
  assign s_CSAwallace_rca24_and_13_1 = a[13] & b[1];
  assign s_CSAwallace_rca24_and_14_1 = a[14] & b[1];
  assign s_CSAwallace_rca24_and_15_1 = a[15] & b[1];
  assign s_CSAwallace_rca24_and_16_1 = a[16] & b[1];
  assign s_CSAwallace_rca24_and_17_1 = a[17] & b[1];
  assign s_CSAwallace_rca24_and_18_1 = a[18] & b[1];
  assign s_CSAwallace_rca24_and_19_1 = a[19] & b[1];
  assign s_CSAwallace_rca24_and_20_1 = a[20] & b[1];
  assign s_CSAwallace_rca24_and_21_1 = a[21] & b[1];
  assign s_CSAwallace_rca24_and_22_1 = a[22] & b[1];
  assign s_CSAwallace_rca24_nand_23_1 = ~(a[23] & b[1]);
  assign s_CSAwallace_rca24_and_0_2 = a[0] & b[2];
  assign s_CSAwallace_rca24_and_1_2 = a[1] & b[2];
  assign s_CSAwallace_rca24_and_2_2 = a[2] & b[2];
  assign s_CSAwallace_rca24_and_3_2 = a[3] & b[2];
  assign s_CSAwallace_rca24_and_4_2 = a[4] & b[2];
  assign s_CSAwallace_rca24_and_5_2 = a[5] & b[2];
  assign s_CSAwallace_rca24_and_6_2 = a[6] & b[2];
  assign s_CSAwallace_rca24_and_7_2 = a[7] & b[2];
  assign s_CSAwallace_rca24_and_8_2 = a[8] & b[2];
  assign s_CSAwallace_rca24_and_9_2 = a[9] & b[2];
  assign s_CSAwallace_rca24_and_10_2 = a[10] & b[2];
  assign s_CSAwallace_rca24_and_11_2 = a[11] & b[2];
  assign s_CSAwallace_rca24_and_12_2 = a[12] & b[2];
  assign s_CSAwallace_rca24_and_13_2 = a[13] & b[2];
  assign s_CSAwallace_rca24_and_14_2 = a[14] & b[2];
  assign s_CSAwallace_rca24_and_15_2 = a[15] & b[2];
  assign s_CSAwallace_rca24_and_16_2 = a[16] & b[2];
  assign s_CSAwallace_rca24_and_17_2 = a[17] & b[2];
  assign s_CSAwallace_rca24_and_18_2 = a[18] & b[2];
  assign s_CSAwallace_rca24_and_19_2 = a[19] & b[2];
  assign s_CSAwallace_rca24_and_20_2 = a[20] & b[2];
  assign s_CSAwallace_rca24_and_21_2 = a[21] & b[2];
  assign s_CSAwallace_rca24_and_22_2 = a[22] & b[2];
  assign s_CSAwallace_rca24_nand_23_2 = ~(a[23] & b[2]);
  assign s_CSAwallace_rca24_and_0_3 = a[0] & b[3];
  assign s_CSAwallace_rca24_and_1_3 = a[1] & b[3];
  assign s_CSAwallace_rca24_and_2_3 = a[2] & b[3];
  assign s_CSAwallace_rca24_and_3_3 = a[3] & b[3];
  assign s_CSAwallace_rca24_and_4_3 = a[4] & b[3];
  assign s_CSAwallace_rca24_and_5_3 = a[5] & b[3];
  assign s_CSAwallace_rca24_and_6_3 = a[6] & b[3];
  assign s_CSAwallace_rca24_and_7_3 = a[7] & b[3];
  assign s_CSAwallace_rca24_and_8_3 = a[8] & b[3];
  assign s_CSAwallace_rca24_and_9_3 = a[9] & b[3];
  assign s_CSAwallace_rca24_and_10_3 = a[10] & b[3];
  assign s_CSAwallace_rca24_and_11_3 = a[11] & b[3];
  assign s_CSAwallace_rca24_and_12_3 = a[12] & b[3];
  assign s_CSAwallace_rca24_and_13_3 = a[13] & b[3];
  assign s_CSAwallace_rca24_and_14_3 = a[14] & b[3];
  assign s_CSAwallace_rca24_and_15_3 = a[15] & b[3];
  assign s_CSAwallace_rca24_and_16_3 = a[16] & b[3];
  assign s_CSAwallace_rca24_and_17_3 = a[17] & b[3];
  assign s_CSAwallace_rca24_and_18_3 = a[18] & b[3];
  assign s_CSAwallace_rca24_and_19_3 = a[19] & b[3];
  assign s_CSAwallace_rca24_and_20_3 = a[20] & b[3];
  assign s_CSAwallace_rca24_and_21_3 = a[21] & b[3];
  assign s_CSAwallace_rca24_and_22_3 = a[22] & b[3];
  assign s_CSAwallace_rca24_nand_23_3 = ~(a[23] & b[3]);
  assign s_CSAwallace_rca24_and_0_4 = a[0] & b[4];
  assign s_CSAwallace_rca24_and_1_4 = a[1] & b[4];
  assign s_CSAwallace_rca24_and_2_4 = a[2] & b[4];
  assign s_CSAwallace_rca24_and_3_4 = a[3] & b[4];
  assign s_CSAwallace_rca24_and_4_4 = a[4] & b[4];
  assign s_CSAwallace_rca24_and_5_4 = a[5] & b[4];
  assign s_CSAwallace_rca24_and_6_4 = a[6] & b[4];
  assign s_CSAwallace_rca24_and_7_4 = a[7] & b[4];
  assign s_CSAwallace_rca24_and_8_4 = a[8] & b[4];
  assign s_CSAwallace_rca24_and_9_4 = a[9] & b[4];
  assign s_CSAwallace_rca24_and_10_4 = a[10] & b[4];
  assign s_CSAwallace_rca24_and_11_4 = a[11] & b[4];
  assign s_CSAwallace_rca24_and_12_4 = a[12] & b[4];
  assign s_CSAwallace_rca24_and_13_4 = a[13] & b[4];
  assign s_CSAwallace_rca24_and_14_4 = a[14] & b[4];
  assign s_CSAwallace_rca24_and_15_4 = a[15] & b[4];
  assign s_CSAwallace_rca24_and_16_4 = a[16] & b[4];
  assign s_CSAwallace_rca24_and_17_4 = a[17] & b[4];
  assign s_CSAwallace_rca24_and_18_4 = a[18] & b[4];
  assign s_CSAwallace_rca24_and_19_4 = a[19] & b[4];
  assign s_CSAwallace_rca24_and_20_4 = a[20] & b[4];
  assign s_CSAwallace_rca24_and_21_4 = a[21] & b[4];
  assign s_CSAwallace_rca24_and_22_4 = a[22] & b[4];
  assign s_CSAwallace_rca24_nand_23_4 = ~(a[23] & b[4]);
  assign s_CSAwallace_rca24_and_0_5 = a[0] & b[5];
  assign s_CSAwallace_rca24_and_1_5 = a[1] & b[5];
  assign s_CSAwallace_rca24_and_2_5 = a[2] & b[5];
  assign s_CSAwallace_rca24_and_3_5 = a[3] & b[5];
  assign s_CSAwallace_rca24_and_4_5 = a[4] & b[5];
  assign s_CSAwallace_rca24_and_5_5 = a[5] & b[5];
  assign s_CSAwallace_rca24_and_6_5 = a[6] & b[5];
  assign s_CSAwallace_rca24_and_7_5 = a[7] & b[5];
  assign s_CSAwallace_rca24_and_8_5 = a[8] & b[5];
  assign s_CSAwallace_rca24_and_9_5 = a[9] & b[5];
  assign s_CSAwallace_rca24_and_10_5 = a[10] & b[5];
  assign s_CSAwallace_rca24_and_11_5 = a[11] & b[5];
  assign s_CSAwallace_rca24_and_12_5 = a[12] & b[5];
  assign s_CSAwallace_rca24_and_13_5 = a[13] & b[5];
  assign s_CSAwallace_rca24_and_14_5 = a[14] & b[5];
  assign s_CSAwallace_rca24_and_15_5 = a[15] & b[5];
  assign s_CSAwallace_rca24_and_16_5 = a[16] & b[5];
  assign s_CSAwallace_rca24_and_17_5 = a[17] & b[5];
  assign s_CSAwallace_rca24_and_18_5 = a[18] & b[5];
  assign s_CSAwallace_rca24_and_19_5 = a[19] & b[5];
  assign s_CSAwallace_rca24_and_20_5 = a[20] & b[5];
  assign s_CSAwallace_rca24_and_21_5 = a[21] & b[5];
  assign s_CSAwallace_rca24_and_22_5 = a[22] & b[5];
  assign s_CSAwallace_rca24_nand_23_5 = ~(a[23] & b[5]);
  assign s_CSAwallace_rca24_and_0_6 = a[0] & b[6];
  assign s_CSAwallace_rca24_and_1_6 = a[1] & b[6];
  assign s_CSAwallace_rca24_and_2_6 = a[2] & b[6];
  assign s_CSAwallace_rca24_and_3_6 = a[3] & b[6];
  assign s_CSAwallace_rca24_and_4_6 = a[4] & b[6];
  assign s_CSAwallace_rca24_and_5_6 = a[5] & b[6];
  assign s_CSAwallace_rca24_and_6_6 = a[6] & b[6];
  assign s_CSAwallace_rca24_and_7_6 = a[7] & b[6];
  assign s_CSAwallace_rca24_and_8_6 = a[8] & b[6];
  assign s_CSAwallace_rca24_and_9_6 = a[9] & b[6];
  assign s_CSAwallace_rca24_and_10_6 = a[10] & b[6];
  assign s_CSAwallace_rca24_and_11_6 = a[11] & b[6];
  assign s_CSAwallace_rca24_and_12_6 = a[12] & b[6];
  assign s_CSAwallace_rca24_and_13_6 = a[13] & b[6];
  assign s_CSAwallace_rca24_and_14_6 = a[14] & b[6];
  assign s_CSAwallace_rca24_and_15_6 = a[15] & b[6];
  assign s_CSAwallace_rca24_and_16_6 = a[16] & b[6];
  assign s_CSAwallace_rca24_and_17_6 = a[17] & b[6];
  assign s_CSAwallace_rca24_and_18_6 = a[18] & b[6];
  assign s_CSAwallace_rca24_and_19_6 = a[19] & b[6];
  assign s_CSAwallace_rca24_and_20_6 = a[20] & b[6];
  assign s_CSAwallace_rca24_and_21_6 = a[21] & b[6];
  assign s_CSAwallace_rca24_and_22_6 = a[22] & b[6];
  assign s_CSAwallace_rca24_nand_23_6 = ~(a[23] & b[6]);
  assign s_CSAwallace_rca24_and_0_7 = a[0] & b[7];
  assign s_CSAwallace_rca24_and_1_7 = a[1] & b[7];
  assign s_CSAwallace_rca24_and_2_7 = a[2] & b[7];
  assign s_CSAwallace_rca24_and_3_7 = a[3] & b[7];
  assign s_CSAwallace_rca24_and_4_7 = a[4] & b[7];
  assign s_CSAwallace_rca24_and_5_7 = a[5] & b[7];
  assign s_CSAwallace_rca24_and_6_7 = a[6] & b[7];
  assign s_CSAwallace_rca24_and_7_7 = a[7] & b[7];
  assign s_CSAwallace_rca24_and_8_7 = a[8] & b[7];
  assign s_CSAwallace_rca24_and_9_7 = a[9] & b[7];
  assign s_CSAwallace_rca24_and_10_7 = a[10] & b[7];
  assign s_CSAwallace_rca24_and_11_7 = a[11] & b[7];
  assign s_CSAwallace_rca24_and_12_7 = a[12] & b[7];
  assign s_CSAwallace_rca24_and_13_7 = a[13] & b[7];
  assign s_CSAwallace_rca24_and_14_7 = a[14] & b[7];
  assign s_CSAwallace_rca24_and_15_7 = a[15] & b[7];
  assign s_CSAwallace_rca24_and_16_7 = a[16] & b[7];
  assign s_CSAwallace_rca24_and_17_7 = a[17] & b[7];
  assign s_CSAwallace_rca24_and_18_7 = a[18] & b[7];
  assign s_CSAwallace_rca24_and_19_7 = a[19] & b[7];
  assign s_CSAwallace_rca24_and_20_7 = a[20] & b[7];
  assign s_CSAwallace_rca24_and_21_7 = a[21] & b[7];
  assign s_CSAwallace_rca24_and_22_7 = a[22] & b[7];
  assign s_CSAwallace_rca24_nand_23_7 = ~(a[23] & b[7]);
  assign s_CSAwallace_rca24_and_0_8 = a[0] & b[8];
  assign s_CSAwallace_rca24_and_1_8 = a[1] & b[8];
  assign s_CSAwallace_rca24_and_2_8 = a[2] & b[8];
  assign s_CSAwallace_rca24_and_3_8 = a[3] & b[8];
  assign s_CSAwallace_rca24_and_4_8 = a[4] & b[8];
  assign s_CSAwallace_rca24_and_5_8 = a[5] & b[8];
  assign s_CSAwallace_rca24_and_6_8 = a[6] & b[8];
  assign s_CSAwallace_rca24_and_7_8 = a[7] & b[8];
  assign s_CSAwallace_rca24_and_8_8 = a[8] & b[8];
  assign s_CSAwallace_rca24_and_9_8 = a[9] & b[8];
  assign s_CSAwallace_rca24_and_10_8 = a[10] & b[8];
  assign s_CSAwallace_rca24_and_11_8 = a[11] & b[8];
  assign s_CSAwallace_rca24_and_12_8 = a[12] & b[8];
  assign s_CSAwallace_rca24_and_13_8 = a[13] & b[8];
  assign s_CSAwallace_rca24_and_14_8 = a[14] & b[8];
  assign s_CSAwallace_rca24_and_15_8 = a[15] & b[8];
  assign s_CSAwallace_rca24_and_16_8 = a[16] & b[8];
  assign s_CSAwallace_rca24_and_17_8 = a[17] & b[8];
  assign s_CSAwallace_rca24_and_18_8 = a[18] & b[8];
  assign s_CSAwallace_rca24_and_19_8 = a[19] & b[8];
  assign s_CSAwallace_rca24_and_20_8 = a[20] & b[8];
  assign s_CSAwallace_rca24_and_21_8 = a[21] & b[8];
  assign s_CSAwallace_rca24_and_22_8 = a[22] & b[8];
  assign s_CSAwallace_rca24_nand_23_8 = ~(a[23] & b[8]);
  assign s_CSAwallace_rca24_and_0_9 = a[0] & b[9];
  assign s_CSAwallace_rca24_and_1_9 = a[1] & b[9];
  assign s_CSAwallace_rca24_and_2_9 = a[2] & b[9];
  assign s_CSAwallace_rca24_and_3_9 = a[3] & b[9];
  assign s_CSAwallace_rca24_and_4_9 = a[4] & b[9];
  assign s_CSAwallace_rca24_and_5_9 = a[5] & b[9];
  assign s_CSAwallace_rca24_and_6_9 = a[6] & b[9];
  assign s_CSAwallace_rca24_and_7_9 = a[7] & b[9];
  assign s_CSAwallace_rca24_and_8_9 = a[8] & b[9];
  assign s_CSAwallace_rca24_and_9_9 = a[9] & b[9];
  assign s_CSAwallace_rca24_and_10_9 = a[10] & b[9];
  assign s_CSAwallace_rca24_and_11_9 = a[11] & b[9];
  assign s_CSAwallace_rca24_and_12_9 = a[12] & b[9];
  assign s_CSAwallace_rca24_and_13_9 = a[13] & b[9];
  assign s_CSAwallace_rca24_and_14_9 = a[14] & b[9];
  assign s_CSAwallace_rca24_and_15_9 = a[15] & b[9];
  assign s_CSAwallace_rca24_and_16_9 = a[16] & b[9];
  assign s_CSAwallace_rca24_and_17_9 = a[17] & b[9];
  assign s_CSAwallace_rca24_and_18_9 = a[18] & b[9];
  assign s_CSAwallace_rca24_and_19_9 = a[19] & b[9];
  assign s_CSAwallace_rca24_and_20_9 = a[20] & b[9];
  assign s_CSAwallace_rca24_and_21_9 = a[21] & b[9];
  assign s_CSAwallace_rca24_and_22_9 = a[22] & b[9];
  assign s_CSAwallace_rca24_nand_23_9 = ~(a[23] & b[9]);
  assign s_CSAwallace_rca24_and_0_10 = a[0] & b[10];
  assign s_CSAwallace_rca24_and_1_10 = a[1] & b[10];
  assign s_CSAwallace_rca24_and_2_10 = a[2] & b[10];
  assign s_CSAwallace_rca24_and_3_10 = a[3] & b[10];
  assign s_CSAwallace_rca24_and_4_10 = a[4] & b[10];
  assign s_CSAwallace_rca24_and_5_10 = a[5] & b[10];
  assign s_CSAwallace_rca24_and_6_10 = a[6] & b[10];
  assign s_CSAwallace_rca24_and_7_10 = a[7] & b[10];
  assign s_CSAwallace_rca24_and_8_10 = a[8] & b[10];
  assign s_CSAwallace_rca24_and_9_10 = a[9] & b[10];
  assign s_CSAwallace_rca24_and_10_10 = a[10] & b[10];
  assign s_CSAwallace_rca24_and_11_10 = a[11] & b[10];
  assign s_CSAwallace_rca24_and_12_10 = a[12] & b[10];
  assign s_CSAwallace_rca24_and_13_10 = a[13] & b[10];
  assign s_CSAwallace_rca24_and_14_10 = a[14] & b[10];
  assign s_CSAwallace_rca24_and_15_10 = a[15] & b[10];
  assign s_CSAwallace_rca24_and_16_10 = a[16] & b[10];
  assign s_CSAwallace_rca24_and_17_10 = a[17] & b[10];
  assign s_CSAwallace_rca24_and_18_10 = a[18] & b[10];
  assign s_CSAwallace_rca24_and_19_10 = a[19] & b[10];
  assign s_CSAwallace_rca24_and_20_10 = a[20] & b[10];
  assign s_CSAwallace_rca24_and_21_10 = a[21] & b[10];
  assign s_CSAwallace_rca24_and_22_10 = a[22] & b[10];
  assign s_CSAwallace_rca24_nand_23_10 = ~(a[23] & b[10]);
  assign s_CSAwallace_rca24_and_0_11 = a[0] & b[11];
  assign s_CSAwallace_rca24_and_1_11 = a[1] & b[11];
  assign s_CSAwallace_rca24_and_2_11 = a[2] & b[11];
  assign s_CSAwallace_rca24_and_3_11 = a[3] & b[11];
  assign s_CSAwallace_rca24_and_4_11 = a[4] & b[11];
  assign s_CSAwallace_rca24_and_5_11 = a[5] & b[11];
  assign s_CSAwallace_rca24_and_6_11 = a[6] & b[11];
  assign s_CSAwallace_rca24_and_7_11 = a[7] & b[11];
  assign s_CSAwallace_rca24_and_8_11 = a[8] & b[11];
  assign s_CSAwallace_rca24_and_9_11 = a[9] & b[11];
  assign s_CSAwallace_rca24_and_10_11 = a[10] & b[11];
  assign s_CSAwallace_rca24_and_11_11 = a[11] & b[11];
  assign s_CSAwallace_rca24_and_12_11 = a[12] & b[11];
  assign s_CSAwallace_rca24_and_13_11 = a[13] & b[11];
  assign s_CSAwallace_rca24_and_14_11 = a[14] & b[11];
  assign s_CSAwallace_rca24_and_15_11 = a[15] & b[11];
  assign s_CSAwallace_rca24_and_16_11 = a[16] & b[11];
  assign s_CSAwallace_rca24_and_17_11 = a[17] & b[11];
  assign s_CSAwallace_rca24_and_18_11 = a[18] & b[11];
  assign s_CSAwallace_rca24_and_19_11 = a[19] & b[11];
  assign s_CSAwallace_rca24_and_20_11 = a[20] & b[11];
  assign s_CSAwallace_rca24_and_21_11 = a[21] & b[11];
  assign s_CSAwallace_rca24_and_22_11 = a[22] & b[11];
  assign s_CSAwallace_rca24_nand_23_11 = ~(a[23] & b[11]);
  assign s_CSAwallace_rca24_and_0_12 = a[0] & b[12];
  assign s_CSAwallace_rca24_and_1_12 = a[1] & b[12];
  assign s_CSAwallace_rca24_and_2_12 = a[2] & b[12];
  assign s_CSAwallace_rca24_and_3_12 = a[3] & b[12];
  assign s_CSAwallace_rca24_and_4_12 = a[4] & b[12];
  assign s_CSAwallace_rca24_and_5_12 = a[5] & b[12];
  assign s_CSAwallace_rca24_and_6_12 = a[6] & b[12];
  assign s_CSAwallace_rca24_and_7_12 = a[7] & b[12];
  assign s_CSAwallace_rca24_and_8_12 = a[8] & b[12];
  assign s_CSAwallace_rca24_and_9_12 = a[9] & b[12];
  assign s_CSAwallace_rca24_and_10_12 = a[10] & b[12];
  assign s_CSAwallace_rca24_and_11_12 = a[11] & b[12];
  assign s_CSAwallace_rca24_and_12_12 = a[12] & b[12];
  assign s_CSAwallace_rca24_and_13_12 = a[13] & b[12];
  assign s_CSAwallace_rca24_and_14_12 = a[14] & b[12];
  assign s_CSAwallace_rca24_and_15_12 = a[15] & b[12];
  assign s_CSAwallace_rca24_and_16_12 = a[16] & b[12];
  assign s_CSAwallace_rca24_and_17_12 = a[17] & b[12];
  assign s_CSAwallace_rca24_and_18_12 = a[18] & b[12];
  assign s_CSAwallace_rca24_and_19_12 = a[19] & b[12];
  assign s_CSAwallace_rca24_and_20_12 = a[20] & b[12];
  assign s_CSAwallace_rca24_and_21_12 = a[21] & b[12];
  assign s_CSAwallace_rca24_and_22_12 = a[22] & b[12];
  assign s_CSAwallace_rca24_nand_23_12 = ~(a[23] & b[12]);
  assign s_CSAwallace_rca24_and_0_13 = a[0] & b[13];
  assign s_CSAwallace_rca24_and_1_13 = a[1] & b[13];
  assign s_CSAwallace_rca24_and_2_13 = a[2] & b[13];
  assign s_CSAwallace_rca24_and_3_13 = a[3] & b[13];
  assign s_CSAwallace_rca24_and_4_13 = a[4] & b[13];
  assign s_CSAwallace_rca24_and_5_13 = a[5] & b[13];
  assign s_CSAwallace_rca24_and_6_13 = a[6] & b[13];
  assign s_CSAwallace_rca24_and_7_13 = a[7] & b[13];
  assign s_CSAwallace_rca24_and_8_13 = a[8] & b[13];
  assign s_CSAwallace_rca24_and_9_13 = a[9] & b[13];
  assign s_CSAwallace_rca24_and_10_13 = a[10] & b[13];
  assign s_CSAwallace_rca24_and_11_13 = a[11] & b[13];
  assign s_CSAwallace_rca24_and_12_13 = a[12] & b[13];
  assign s_CSAwallace_rca24_and_13_13 = a[13] & b[13];
  assign s_CSAwallace_rca24_and_14_13 = a[14] & b[13];
  assign s_CSAwallace_rca24_and_15_13 = a[15] & b[13];
  assign s_CSAwallace_rca24_and_16_13 = a[16] & b[13];
  assign s_CSAwallace_rca24_and_17_13 = a[17] & b[13];
  assign s_CSAwallace_rca24_and_18_13 = a[18] & b[13];
  assign s_CSAwallace_rca24_and_19_13 = a[19] & b[13];
  assign s_CSAwallace_rca24_and_20_13 = a[20] & b[13];
  assign s_CSAwallace_rca24_and_21_13 = a[21] & b[13];
  assign s_CSAwallace_rca24_and_22_13 = a[22] & b[13];
  assign s_CSAwallace_rca24_nand_23_13 = ~(a[23] & b[13]);
  assign s_CSAwallace_rca24_and_0_14 = a[0] & b[14];
  assign s_CSAwallace_rca24_and_1_14 = a[1] & b[14];
  assign s_CSAwallace_rca24_and_2_14 = a[2] & b[14];
  assign s_CSAwallace_rca24_and_3_14 = a[3] & b[14];
  assign s_CSAwallace_rca24_and_4_14 = a[4] & b[14];
  assign s_CSAwallace_rca24_and_5_14 = a[5] & b[14];
  assign s_CSAwallace_rca24_and_6_14 = a[6] & b[14];
  assign s_CSAwallace_rca24_and_7_14 = a[7] & b[14];
  assign s_CSAwallace_rca24_and_8_14 = a[8] & b[14];
  assign s_CSAwallace_rca24_and_9_14 = a[9] & b[14];
  assign s_CSAwallace_rca24_and_10_14 = a[10] & b[14];
  assign s_CSAwallace_rca24_and_11_14 = a[11] & b[14];
  assign s_CSAwallace_rca24_and_12_14 = a[12] & b[14];
  assign s_CSAwallace_rca24_and_13_14 = a[13] & b[14];
  assign s_CSAwallace_rca24_and_14_14 = a[14] & b[14];
  assign s_CSAwallace_rca24_and_15_14 = a[15] & b[14];
  assign s_CSAwallace_rca24_and_16_14 = a[16] & b[14];
  assign s_CSAwallace_rca24_and_17_14 = a[17] & b[14];
  assign s_CSAwallace_rca24_and_18_14 = a[18] & b[14];
  assign s_CSAwallace_rca24_and_19_14 = a[19] & b[14];
  assign s_CSAwallace_rca24_and_20_14 = a[20] & b[14];
  assign s_CSAwallace_rca24_and_21_14 = a[21] & b[14];
  assign s_CSAwallace_rca24_and_22_14 = a[22] & b[14];
  assign s_CSAwallace_rca24_nand_23_14 = ~(a[23] & b[14]);
  assign s_CSAwallace_rca24_and_0_15 = a[0] & b[15];
  assign s_CSAwallace_rca24_and_1_15 = a[1] & b[15];
  assign s_CSAwallace_rca24_and_2_15 = a[2] & b[15];
  assign s_CSAwallace_rca24_and_3_15 = a[3] & b[15];
  assign s_CSAwallace_rca24_and_4_15 = a[4] & b[15];
  assign s_CSAwallace_rca24_and_5_15 = a[5] & b[15];
  assign s_CSAwallace_rca24_and_6_15 = a[6] & b[15];
  assign s_CSAwallace_rca24_and_7_15 = a[7] & b[15];
  assign s_CSAwallace_rca24_and_8_15 = a[8] & b[15];
  assign s_CSAwallace_rca24_and_9_15 = a[9] & b[15];
  assign s_CSAwallace_rca24_and_10_15 = a[10] & b[15];
  assign s_CSAwallace_rca24_and_11_15 = a[11] & b[15];
  assign s_CSAwallace_rca24_and_12_15 = a[12] & b[15];
  assign s_CSAwallace_rca24_and_13_15 = a[13] & b[15];
  assign s_CSAwallace_rca24_and_14_15 = a[14] & b[15];
  assign s_CSAwallace_rca24_and_15_15 = a[15] & b[15];
  assign s_CSAwallace_rca24_and_16_15 = a[16] & b[15];
  assign s_CSAwallace_rca24_and_17_15 = a[17] & b[15];
  assign s_CSAwallace_rca24_and_18_15 = a[18] & b[15];
  assign s_CSAwallace_rca24_and_19_15 = a[19] & b[15];
  assign s_CSAwallace_rca24_and_20_15 = a[20] & b[15];
  assign s_CSAwallace_rca24_and_21_15 = a[21] & b[15];
  assign s_CSAwallace_rca24_and_22_15 = a[22] & b[15];
  assign s_CSAwallace_rca24_nand_23_15 = ~(a[23] & b[15]);
  assign s_CSAwallace_rca24_and_0_16 = a[0] & b[16];
  assign s_CSAwallace_rca24_and_1_16 = a[1] & b[16];
  assign s_CSAwallace_rca24_and_2_16 = a[2] & b[16];
  assign s_CSAwallace_rca24_and_3_16 = a[3] & b[16];
  assign s_CSAwallace_rca24_and_4_16 = a[4] & b[16];
  assign s_CSAwallace_rca24_and_5_16 = a[5] & b[16];
  assign s_CSAwallace_rca24_and_6_16 = a[6] & b[16];
  assign s_CSAwallace_rca24_and_7_16 = a[7] & b[16];
  assign s_CSAwallace_rca24_and_8_16 = a[8] & b[16];
  assign s_CSAwallace_rca24_and_9_16 = a[9] & b[16];
  assign s_CSAwallace_rca24_and_10_16 = a[10] & b[16];
  assign s_CSAwallace_rca24_and_11_16 = a[11] & b[16];
  assign s_CSAwallace_rca24_and_12_16 = a[12] & b[16];
  assign s_CSAwallace_rca24_and_13_16 = a[13] & b[16];
  assign s_CSAwallace_rca24_and_14_16 = a[14] & b[16];
  assign s_CSAwallace_rca24_and_15_16 = a[15] & b[16];
  assign s_CSAwallace_rca24_and_16_16 = a[16] & b[16];
  assign s_CSAwallace_rca24_and_17_16 = a[17] & b[16];
  assign s_CSAwallace_rca24_and_18_16 = a[18] & b[16];
  assign s_CSAwallace_rca24_and_19_16 = a[19] & b[16];
  assign s_CSAwallace_rca24_and_20_16 = a[20] & b[16];
  assign s_CSAwallace_rca24_and_21_16 = a[21] & b[16];
  assign s_CSAwallace_rca24_and_22_16 = a[22] & b[16];
  assign s_CSAwallace_rca24_nand_23_16 = ~(a[23] & b[16]);
  assign s_CSAwallace_rca24_and_0_17 = a[0] & b[17];
  assign s_CSAwallace_rca24_and_1_17 = a[1] & b[17];
  assign s_CSAwallace_rca24_and_2_17 = a[2] & b[17];
  assign s_CSAwallace_rca24_and_3_17 = a[3] & b[17];
  assign s_CSAwallace_rca24_and_4_17 = a[4] & b[17];
  assign s_CSAwallace_rca24_and_5_17 = a[5] & b[17];
  assign s_CSAwallace_rca24_and_6_17 = a[6] & b[17];
  assign s_CSAwallace_rca24_and_7_17 = a[7] & b[17];
  assign s_CSAwallace_rca24_and_8_17 = a[8] & b[17];
  assign s_CSAwallace_rca24_and_9_17 = a[9] & b[17];
  assign s_CSAwallace_rca24_and_10_17 = a[10] & b[17];
  assign s_CSAwallace_rca24_and_11_17 = a[11] & b[17];
  assign s_CSAwallace_rca24_and_12_17 = a[12] & b[17];
  assign s_CSAwallace_rca24_and_13_17 = a[13] & b[17];
  assign s_CSAwallace_rca24_and_14_17 = a[14] & b[17];
  assign s_CSAwallace_rca24_and_15_17 = a[15] & b[17];
  assign s_CSAwallace_rca24_and_16_17 = a[16] & b[17];
  assign s_CSAwallace_rca24_and_17_17 = a[17] & b[17];
  assign s_CSAwallace_rca24_and_18_17 = a[18] & b[17];
  assign s_CSAwallace_rca24_and_19_17 = a[19] & b[17];
  assign s_CSAwallace_rca24_and_20_17 = a[20] & b[17];
  assign s_CSAwallace_rca24_and_21_17 = a[21] & b[17];
  assign s_CSAwallace_rca24_and_22_17 = a[22] & b[17];
  assign s_CSAwallace_rca24_nand_23_17 = ~(a[23] & b[17]);
  assign s_CSAwallace_rca24_and_0_18 = a[0] & b[18];
  assign s_CSAwallace_rca24_and_1_18 = a[1] & b[18];
  assign s_CSAwallace_rca24_and_2_18 = a[2] & b[18];
  assign s_CSAwallace_rca24_and_3_18 = a[3] & b[18];
  assign s_CSAwallace_rca24_and_4_18 = a[4] & b[18];
  assign s_CSAwallace_rca24_and_5_18 = a[5] & b[18];
  assign s_CSAwallace_rca24_and_6_18 = a[6] & b[18];
  assign s_CSAwallace_rca24_and_7_18 = a[7] & b[18];
  assign s_CSAwallace_rca24_and_8_18 = a[8] & b[18];
  assign s_CSAwallace_rca24_and_9_18 = a[9] & b[18];
  assign s_CSAwallace_rca24_and_10_18 = a[10] & b[18];
  assign s_CSAwallace_rca24_and_11_18 = a[11] & b[18];
  assign s_CSAwallace_rca24_and_12_18 = a[12] & b[18];
  assign s_CSAwallace_rca24_and_13_18 = a[13] & b[18];
  assign s_CSAwallace_rca24_and_14_18 = a[14] & b[18];
  assign s_CSAwallace_rca24_and_15_18 = a[15] & b[18];
  assign s_CSAwallace_rca24_and_16_18 = a[16] & b[18];
  assign s_CSAwallace_rca24_and_17_18 = a[17] & b[18];
  assign s_CSAwallace_rca24_and_18_18 = a[18] & b[18];
  assign s_CSAwallace_rca24_and_19_18 = a[19] & b[18];
  assign s_CSAwallace_rca24_and_20_18 = a[20] & b[18];
  assign s_CSAwallace_rca24_and_21_18 = a[21] & b[18];
  assign s_CSAwallace_rca24_and_22_18 = a[22] & b[18];
  assign s_CSAwallace_rca24_nand_23_18 = ~(a[23] & b[18]);
  assign s_CSAwallace_rca24_and_0_19 = a[0] & b[19];
  assign s_CSAwallace_rca24_and_1_19 = a[1] & b[19];
  assign s_CSAwallace_rca24_and_2_19 = a[2] & b[19];
  assign s_CSAwallace_rca24_and_3_19 = a[3] & b[19];
  assign s_CSAwallace_rca24_and_4_19 = a[4] & b[19];
  assign s_CSAwallace_rca24_and_5_19 = a[5] & b[19];
  assign s_CSAwallace_rca24_and_6_19 = a[6] & b[19];
  assign s_CSAwallace_rca24_and_7_19 = a[7] & b[19];
  assign s_CSAwallace_rca24_and_8_19 = a[8] & b[19];
  assign s_CSAwallace_rca24_and_9_19 = a[9] & b[19];
  assign s_CSAwallace_rca24_and_10_19 = a[10] & b[19];
  assign s_CSAwallace_rca24_and_11_19 = a[11] & b[19];
  assign s_CSAwallace_rca24_and_12_19 = a[12] & b[19];
  assign s_CSAwallace_rca24_and_13_19 = a[13] & b[19];
  assign s_CSAwallace_rca24_and_14_19 = a[14] & b[19];
  assign s_CSAwallace_rca24_and_15_19 = a[15] & b[19];
  assign s_CSAwallace_rca24_and_16_19 = a[16] & b[19];
  assign s_CSAwallace_rca24_and_17_19 = a[17] & b[19];
  assign s_CSAwallace_rca24_and_18_19 = a[18] & b[19];
  assign s_CSAwallace_rca24_and_19_19 = a[19] & b[19];
  assign s_CSAwallace_rca24_and_20_19 = a[20] & b[19];
  assign s_CSAwallace_rca24_and_21_19 = a[21] & b[19];
  assign s_CSAwallace_rca24_and_22_19 = a[22] & b[19];
  assign s_CSAwallace_rca24_nand_23_19 = ~(a[23] & b[19]);
  assign s_CSAwallace_rca24_and_0_20 = a[0] & b[20];
  assign s_CSAwallace_rca24_and_1_20 = a[1] & b[20];
  assign s_CSAwallace_rca24_and_2_20 = a[2] & b[20];
  assign s_CSAwallace_rca24_and_3_20 = a[3] & b[20];
  assign s_CSAwallace_rca24_and_4_20 = a[4] & b[20];
  assign s_CSAwallace_rca24_and_5_20 = a[5] & b[20];
  assign s_CSAwallace_rca24_and_6_20 = a[6] & b[20];
  assign s_CSAwallace_rca24_and_7_20 = a[7] & b[20];
  assign s_CSAwallace_rca24_and_8_20 = a[8] & b[20];
  assign s_CSAwallace_rca24_and_9_20 = a[9] & b[20];
  assign s_CSAwallace_rca24_and_10_20 = a[10] & b[20];
  assign s_CSAwallace_rca24_and_11_20 = a[11] & b[20];
  assign s_CSAwallace_rca24_and_12_20 = a[12] & b[20];
  assign s_CSAwallace_rca24_and_13_20 = a[13] & b[20];
  assign s_CSAwallace_rca24_and_14_20 = a[14] & b[20];
  assign s_CSAwallace_rca24_and_15_20 = a[15] & b[20];
  assign s_CSAwallace_rca24_and_16_20 = a[16] & b[20];
  assign s_CSAwallace_rca24_and_17_20 = a[17] & b[20];
  assign s_CSAwallace_rca24_and_18_20 = a[18] & b[20];
  assign s_CSAwallace_rca24_and_19_20 = a[19] & b[20];
  assign s_CSAwallace_rca24_and_20_20 = a[20] & b[20];
  assign s_CSAwallace_rca24_and_21_20 = a[21] & b[20];
  assign s_CSAwallace_rca24_and_22_20 = a[22] & b[20];
  assign s_CSAwallace_rca24_nand_23_20 = ~(a[23] & b[20]);
  assign s_CSAwallace_rca24_and_0_21 = a[0] & b[21];
  assign s_CSAwallace_rca24_and_1_21 = a[1] & b[21];
  assign s_CSAwallace_rca24_and_2_21 = a[2] & b[21];
  assign s_CSAwallace_rca24_and_3_21 = a[3] & b[21];
  assign s_CSAwallace_rca24_and_4_21 = a[4] & b[21];
  assign s_CSAwallace_rca24_and_5_21 = a[5] & b[21];
  assign s_CSAwallace_rca24_and_6_21 = a[6] & b[21];
  assign s_CSAwallace_rca24_and_7_21 = a[7] & b[21];
  assign s_CSAwallace_rca24_and_8_21 = a[8] & b[21];
  assign s_CSAwallace_rca24_and_9_21 = a[9] & b[21];
  assign s_CSAwallace_rca24_and_10_21 = a[10] & b[21];
  assign s_CSAwallace_rca24_and_11_21 = a[11] & b[21];
  assign s_CSAwallace_rca24_and_12_21 = a[12] & b[21];
  assign s_CSAwallace_rca24_and_13_21 = a[13] & b[21];
  assign s_CSAwallace_rca24_and_14_21 = a[14] & b[21];
  assign s_CSAwallace_rca24_and_15_21 = a[15] & b[21];
  assign s_CSAwallace_rca24_and_16_21 = a[16] & b[21];
  assign s_CSAwallace_rca24_and_17_21 = a[17] & b[21];
  assign s_CSAwallace_rca24_and_18_21 = a[18] & b[21];
  assign s_CSAwallace_rca24_and_19_21 = a[19] & b[21];
  assign s_CSAwallace_rca24_and_20_21 = a[20] & b[21];
  assign s_CSAwallace_rca24_and_21_21 = a[21] & b[21];
  assign s_CSAwallace_rca24_and_22_21 = a[22] & b[21];
  assign s_CSAwallace_rca24_nand_23_21 = ~(a[23] & b[21]);
  assign s_CSAwallace_rca24_and_0_22 = a[0] & b[22];
  assign s_CSAwallace_rca24_and_1_22 = a[1] & b[22];
  assign s_CSAwallace_rca24_and_2_22 = a[2] & b[22];
  assign s_CSAwallace_rca24_and_3_22 = a[3] & b[22];
  assign s_CSAwallace_rca24_and_4_22 = a[4] & b[22];
  assign s_CSAwallace_rca24_and_5_22 = a[5] & b[22];
  assign s_CSAwallace_rca24_and_6_22 = a[6] & b[22];
  assign s_CSAwallace_rca24_and_7_22 = a[7] & b[22];
  assign s_CSAwallace_rca24_and_8_22 = a[8] & b[22];
  assign s_CSAwallace_rca24_and_9_22 = a[9] & b[22];
  assign s_CSAwallace_rca24_and_10_22 = a[10] & b[22];
  assign s_CSAwallace_rca24_and_11_22 = a[11] & b[22];
  assign s_CSAwallace_rca24_and_12_22 = a[12] & b[22];
  assign s_CSAwallace_rca24_and_13_22 = a[13] & b[22];
  assign s_CSAwallace_rca24_and_14_22 = a[14] & b[22];
  assign s_CSAwallace_rca24_and_15_22 = a[15] & b[22];
  assign s_CSAwallace_rca24_and_16_22 = a[16] & b[22];
  assign s_CSAwallace_rca24_and_17_22 = a[17] & b[22];
  assign s_CSAwallace_rca24_and_18_22 = a[18] & b[22];
  assign s_CSAwallace_rca24_and_19_22 = a[19] & b[22];
  assign s_CSAwallace_rca24_and_20_22 = a[20] & b[22];
  assign s_CSAwallace_rca24_and_21_22 = a[21] & b[22];
  assign s_CSAwallace_rca24_and_22_22 = a[22] & b[22];
  assign s_CSAwallace_rca24_nand_23_22 = ~(a[23] & b[22]);
  assign s_CSAwallace_rca24_nand_0_23 = ~(a[0] & b[23]);
  assign s_CSAwallace_rca24_nand_1_23 = ~(a[1] & b[23]);
  assign s_CSAwallace_rca24_nand_2_23 = ~(a[2] & b[23]);
  assign s_CSAwallace_rca24_nand_3_23 = ~(a[3] & b[23]);
  assign s_CSAwallace_rca24_nand_4_23 = ~(a[4] & b[23]);
  assign s_CSAwallace_rca24_nand_5_23 = ~(a[5] & b[23]);
  assign s_CSAwallace_rca24_nand_6_23 = ~(a[6] & b[23]);
  assign s_CSAwallace_rca24_nand_7_23 = ~(a[7] & b[23]);
  assign s_CSAwallace_rca24_nand_8_23 = ~(a[8] & b[23]);
  assign s_CSAwallace_rca24_nand_9_23 = ~(a[9] & b[23]);
  assign s_CSAwallace_rca24_nand_10_23 = ~(a[10] & b[23]);
  assign s_CSAwallace_rca24_nand_11_23 = ~(a[11] & b[23]);
  assign s_CSAwallace_rca24_nand_12_23 = ~(a[12] & b[23]);
  assign s_CSAwallace_rca24_nand_13_23 = ~(a[13] & b[23]);
  assign s_CSAwallace_rca24_nand_14_23 = ~(a[14] & b[23]);
  assign s_CSAwallace_rca24_nand_15_23 = ~(a[15] & b[23]);
  assign s_CSAwallace_rca24_nand_16_23 = ~(a[16] & b[23]);
  assign s_CSAwallace_rca24_nand_17_23 = ~(a[17] & b[23]);
  assign s_CSAwallace_rca24_nand_18_23 = ~(a[18] & b[23]);
  assign s_CSAwallace_rca24_nand_19_23 = ~(a[19] & b[23]);
  assign s_CSAwallace_rca24_nand_20_23 = ~(a[20] & b[23]);
  assign s_CSAwallace_rca24_nand_21_23 = ~(a[21] & b[23]);
  assign s_CSAwallace_rca24_nand_22_23 = ~(a[22] & b[23]);
  assign s_CSAwallace_rca24_and_23_23 = a[23] & b[23];
  assign s_CSAwallace_rca24_csa0_csa_component_fa1_xor0 = s_CSAwallace_rca24_and_1_0 ^ s_CSAwallace_rca24_and_0_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa1_and0 = s_CSAwallace_rca24_and_1_0 & s_CSAwallace_rca24_and_0_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa2_xor0 = s_CSAwallace_rca24_and_2_0 ^ s_CSAwallace_rca24_and_1_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa2_and0 = s_CSAwallace_rca24_and_2_0 & s_CSAwallace_rca24_and_1_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa2_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa2_xor0 ^ s_CSAwallace_rca24_and_0_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa2_and1 = s_CSAwallace_rca24_csa0_csa_component_fa2_xor0 & s_CSAwallace_rca24_and_0_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa2_or0 = s_CSAwallace_rca24_csa0_csa_component_fa2_and0 | s_CSAwallace_rca24_csa0_csa_component_fa2_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa3_xor0 = s_CSAwallace_rca24_and_3_0 ^ s_CSAwallace_rca24_and_2_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa3_and0 = s_CSAwallace_rca24_and_3_0 & s_CSAwallace_rca24_and_2_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa3_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa3_xor0 ^ s_CSAwallace_rca24_and_1_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa3_and1 = s_CSAwallace_rca24_csa0_csa_component_fa3_xor0 & s_CSAwallace_rca24_and_1_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa3_or0 = s_CSAwallace_rca24_csa0_csa_component_fa3_and0 | s_CSAwallace_rca24_csa0_csa_component_fa3_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa4_xor0 = s_CSAwallace_rca24_and_4_0 ^ s_CSAwallace_rca24_and_3_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa4_and0 = s_CSAwallace_rca24_and_4_0 & s_CSAwallace_rca24_and_3_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa4_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa4_xor0 ^ s_CSAwallace_rca24_and_2_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa4_and1 = s_CSAwallace_rca24_csa0_csa_component_fa4_xor0 & s_CSAwallace_rca24_and_2_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa4_or0 = s_CSAwallace_rca24_csa0_csa_component_fa4_and0 | s_CSAwallace_rca24_csa0_csa_component_fa4_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa5_xor0 = s_CSAwallace_rca24_and_5_0 ^ s_CSAwallace_rca24_and_4_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa5_and0 = s_CSAwallace_rca24_and_5_0 & s_CSAwallace_rca24_and_4_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa5_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa5_xor0 ^ s_CSAwallace_rca24_and_3_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa5_and1 = s_CSAwallace_rca24_csa0_csa_component_fa5_xor0 & s_CSAwallace_rca24_and_3_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa5_or0 = s_CSAwallace_rca24_csa0_csa_component_fa5_and0 | s_CSAwallace_rca24_csa0_csa_component_fa5_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa6_xor0 = s_CSAwallace_rca24_and_6_0 ^ s_CSAwallace_rca24_and_5_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa6_and0 = s_CSAwallace_rca24_and_6_0 & s_CSAwallace_rca24_and_5_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa6_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa6_xor0 ^ s_CSAwallace_rca24_and_4_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa6_and1 = s_CSAwallace_rca24_csa0_csa_component_fa6_xor0 & s_CSAwallace_rca24_and_4_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa6_or0 = s_CSAwallace_rca24_csa0_csa_component_fa6_and0 | s_CSAwallace_rca24_csa0_csa_component_fa6_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa7_xor0 = s_CSAwallace_rca24_and_7_0 ^ s_CSAwallace_rca24_and_6_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa7_and0 = s_CSAwallace_rca24_and_7_0 & s_CSAwallace_rca24_and_6_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa7_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa7_xor0 ^ s_CSAwallace_rca24_and_5_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa7_and1 = s_CSAwallace_rca24_csa0_csa_component_fa7_xor0 & s_CSAwallace_rca24_and_5_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa7_or0 = s_CSAwallace_rca24_csa0_csa_component_fa7_and0 | s_CSAwallace_rca24_csa0_csa_component_fa7_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa8_xor0 = s_CSAwallace_rca24_and_8_0 ^ s_CSAwallace_rca24_and_7_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa8_and0 = s_CSAwallace_rca24_and_8_0 & s_CSAwallace_rca24_and_7_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa8_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_and_6_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa8_and1 = s_CSAwallace_rca24_csa0_csa_component_fa8_xor0 & s_CSAwallace_rca24_and_6_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa8_or0 = s_CSAwallace_rca24_csa0_csa_component_fa8_and0 | s_CSAwallace_rca24_csa0_csa_component_fa8_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa9_xor0 = s_CSAwallace_rca24_and_9_0 ^ s_CSAwallace_rca24_and_8_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa9_and0 = s_CSAwallace_rca24_and_9_0 & s_CSAwallace_rca24_and_8_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa9_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_and_7_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa9_and1 = s_CSAwallace_rca24_csa0_csa_component_fa9_xor0 & s_CSAwallace_rca24_and_7_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa9_or0 = s_CSAwallace_rca24_csa0_csa_component_fa9_and0 | s_CSAwallace_rca24_csa0_csa_component_fa9_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa10_xor0 = s_CSAwallace_rca24_and_10_0 ^ s_CSAwallace_rca24_and_9_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa10_and0 = s_CSAwallace_rca24_and_10_0 & s_CSAwallace_rca24_and_9_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa10_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_and_8_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa10_and1 = s_CSAwallace_rca24_csa0_csa_component_fa10_xor0 & s_CSAwallace_rca24_and_8_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa10_or0 = s_CSAwallace_rca24_csa0_csa_component_fa10_and0 | s_CSAwallace_rca24_csa0_csa_component_fa10_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa11_xor0 = s_CSAwallace_rca24_and_11_0 ^ s_CSAwallace_rca24_and_10_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa11_and0 = s_CSAwallace_rca24_and_11_0 & s_CSAwallace_rca24_and_10_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa11_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_and_9_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa11_and1 = s_CSAwallace_rca24_csa0_csa_component_fa11_xor0 & s_CSAwallace_rca24_and_9_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa11_or0 = s_CSAwallace_rca24_csa0_csa_component_fa11_and0 | s_CSAwallace_rca24_csa0_csa_component_fa11_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa12_xor0 = s_CSAwallace_rca24_and_12_0 ^ s_CSAwallace_rca24_and_11_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa12_and0 = s_CSAwallace_rca24_and_12_0 & s_CSAwallace_rca24_and_11_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_and_10_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa12_and1 = s_CSAwallace_rca24_csa0_csa_component_fa12_xor0 & s_CSAwallace_rca24_and_10_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa12_or0 = s_CSAwallace_rca24_csa0_csa_component_fa12_and0 | s_CSAwallace_rca24_csa0_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa13_xor0 = s_CSAwallace_rca24_and_13_0 ^ s_CSAwallace_rca24_and_12_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa13_and0 = s_CSAwallace_rca24_and_13_0 & s_CSAwallace_rca24_and_12_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_and_11_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa13_and1 = s_CSAwallace_rca24_csa0_csa_component_fa13_xor0 & s_CSAwallace_rca24_and_11_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa13_or0 = s_CSAwallace_rca24_csa0_csa_component_fa13_and0 | s_CSAwallace_rca24_csa0_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa14_xor0 = s_CSAwallace_rca24_and_14_0 ^ s_CSAwallace_rca24_and_13_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa14_and0 = s_CSAwallace_rca24_and_14_0 & s_CSAwallace_rca24_and_13_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_and_12_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa14_and1 = s_CSAwallace_rca24_csa0_csa_component_fa14_xor0 & s_CSAwallace_rca24_and_12_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa14_or0 = s_CSAwallace_rca24_csa0_csa_component_fa14_and0 | s_CSAwallace_rca24_csa0_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa15_xor0 = s_CSAwallace_rca24_and_15_0 ^ s_CSAwallace_rca24_and_14_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa15_and0 = s_CSAwallace_rca24_and_15_0 & s_CSAwallace_rca24_and_14_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_and_13_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa15_and1 = s_CSAwallace_rca24_csa0_csa_component_fa15_xor0 & s_CSAwallace_rca24_and_13_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa15_or0 = s_CSAwallace_rca24_csa0_csa_component_fa15_and0 | s_CSAwallace_rca24_csa0_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa16_xor0 = s_CSAwallace_rca24_and_16_0 ^ s_CSAwallace_rca24_and_15_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa16_and0 = s_CSAwallace_rca24_and_16_0 & s_CSAwallace_rca24_and_15_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_and_14_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa16_and1 = s_CSAwallace_rca24_csa0_csa_component_fa16_xor0 & s_CSAwallace_rca24_and_14_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa16_or0 = s_CSAwallace_rca24_csa0_csa_component_fa16_and0 | s_CSAwallace_rca24_csa0_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa17_xor0 = s_CSAwallace_rca24_and_17_0 ^ s_CSAwallace_rca24_and_16_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa17_and0 = s_CSAwallace_rca24_and_17_0 & s_CSAwallace_rca24_and_16_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_and_15_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa17_and1 = s_CSAwallace_rca24_csa0_csa_component_fa17_xor0 & s_CSAwallace_rca24_and_15_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa17_or0 = s_CSAwallace_rca24_csa0_csa_component_fa17_and0 | s_CSAwallace_rca24_csa0_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa18_xor0 = s_CSAwallace_rca24_and_18_0 ^ s_CSAwallace_rca24_and_17_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa18_and0 = s_CSAwallace_rca24_and_18_0 & s_CSAwallace_rca24_and_17_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_and_16_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa18_and1 = s_CSAwallace_rca24_csa0_csa_component_fa18_xor0 & s_CSAwallace_rca24_and_16_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa18_or0 = s_CSAwallace_rca24_csa0_csa_component_fa18_and0 | s_CSAwallace_rca24_csa0_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa19_xor0 = s_CSAwallace_rca24_and_19_0 ^ s_CSAwallace_rca24_and_18_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa19_and0 = s_CSAwallace_rca24_and_19_0 & s_CSAwallace_rca24_and_18_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_and_17_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa19_and1 = s_CSAwallace_rca24_csa0_csa_component_fa19_xor0 & s_CSAwallace_rca24_and_17_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa19_or0 = s_CSAwallace_rca24_csa0_csa_component_fa19_and0 | s_CSAwallace_rca24_csa0_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa20_xor0 = s_CSAwallace_rca24_and_20_0 ^ s_CSAwallace_rca24_and_19_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa20_and0 = s_CSAwallace_rca24_and_20_0 & s_CSAwallace_rca24_and_19_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_and_18_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa20_and1 = s_CSAwallace_rca24_csa0_csa_component_fa20_xor0 & s_CSAwallace_rca24_and_18_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa20_or0 = s_CSAwallace_rca24_csa0_csa_component_fa20_and0 | s_CSAwallace_rca24_csa0_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa21_xor0 = s_CSAwallace_rca24_and_21_0 ^ s_CSAwallace_rca24_and_20_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa21_and0 = s_CSAwallace_rca24_and_21_0 & s_CSAwallace_rca24_and_20_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_and_19_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa21_and1 = s_CSAwallace_rca24_csa0_csa_component_fa21_xor0 & s_CSAwallace_rca24_and_19_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa21_or0 = s_CSAwallace_rca24_csa0_csa_component_fa21_and0 | s_CSAwallace_rca24_csa0_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa22_xor0 = s_CSAwallace_rca24_and_22_0 ^ s_CSAwallace_rca24_and_21_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa22_and0 = s_CSAwallace_rca24_and_22_0 & s_CSAwallace_rca24_and_21_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_and_20_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa22_and1 = s_CSAwallace_rca24_csa0_csa_component_fa22_xor0 & s_CSAwallace_rca24_and_20_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa22_or0 = s_CSAwallace_rca24_csa0_csa_component_fa22_and0 | s_CSAwallace_rca24_csa0_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa23_xor0 = s_CSAwallace_rca24_nand_23_0 ^ s_CSAwallace_rca24_and_22_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa23_and0 = s_CSAwallace_rca24_nand_23_0 & s_CSAwallace_rca24_and_22_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_and_21_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa23_and1 = s_CSAwallace_rca24_csa0_csa_component_fa23_xor0 & s_CSAwallace_rca24_and_21_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa23_or0 = s_CSAwallace_rca24_csa0_csa_component_fa23_and0 | s_CSAwallace_rca24_csa0_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa24_xor0 = ~s_CSAwallace_rca24_nand_23_1;
  assign s_CSAwallace_rca24_csa0_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa0_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_and_22_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa24_and1 = s_CSAwallace_rca24_csa0_csa_component_fa24_xor0 & s_CSAwallace_rca24_and_22_2;
  assign s_CSAwallace_rca24_csa0_csa_component_fa24_or0 = s_CSAwallace_rca24_nand_23_1 | s_CSAwallace_rca24_csa0_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa4_xor0 = s_CSAwallace_rca24_and_1_3 ^ s_CSAwallace_rca24_and_0_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa4_and0 = s_CSAwallace_rca24_and_1_3 & s_CSAwallace_rca24_and_0_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa5_xor0 = s_CSAwallace_rca24_and_2_3 ^ s_CSAwallace_rca24_and_1_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa5_and0 = s_CSAwallace_rca24_and_2_3 & s_CSAwallace_rca24_and_1_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa5_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa5_xor0 ^ s_CSAwallace_rca24_and_0_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa5_and1 = s_CSAwallace_rca24_csa1_csa_component_fa5_xor0 & s_CSAwallace_rca24_and_0_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa5_or0 = s_CSAwallace_rca24_csa1_csa_component_fa5_and0 | s_CSAwallace_rca24_csa1_csa_component_fa5_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa6_xor0 = s_CSAwallace_rca24_and_3_3 ^ s_CSAwallace_rca24_and_2_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa6_and0 = s_CSAwallace_rca24_and_3_3 & s_CSAwallace_rca24_and_2_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa6_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa6_xor0 ^ s_CSAwallace_rca24_and_1_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa6_and1 = s_CSAwallace_rca24_csa1_csa_component_fa6_xor0 & s_CSAwallace_rca24_and_1_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa6_or0 = s_CSAwallace_rca24_csa1_csa_component_fa6_and0 | s_CSAwallace_rca24_csa1_csa_component_fa6_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa7_xor0 = s_CSAwallace_rca24_and_4_3 ^ s_CSAwallace_rca24_and_3_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa7_and0 = s_CSAwallace_rca24_and_4_3 & s_CSAwallace_rca24_and_3_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa7_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa7_xor0 ^ s_CSAwallace_rca24_and_2_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa7_and1 = s_CSAwallace_rca24_csa1_csa_component_fa7_xor0 & s_CSAwallace_rca24_and_2_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa7_or0 = s_CSAwallace_rca24_csa1_csa_component_fa7_and0 | s_CSAwallace_rca24_csa1_csa_component_fa7_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa8_xor0 = s_CSAwallace_rca24_and_5_3 ^ s_CSAwallace_rca24_and_4_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa8_and0 = s_CSAwallace_rca24_and_5_3 & s_CSAwallace_rca24_and_4_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa8_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_and_3_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa8_and1 = s_CSAwallace_rca24_csa1_csa_component_fa8_xor0 & s_CSAwallace_rca24_and_3_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa8_or0 = s_CSAwallace_rca24_csa1_csa_component_fa8_and0 | s_CSAwallace_rca24_csa1_csa_component_fa8_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa9_xor0 = s_CSAwallace_rca24_and_6_3 ^ s_CSAwallace_rca24_and_5_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa9_and0 = s_CSAwallace_rca24_and_6_3 & s_CSAwallace_rca24_and_5_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa9_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_and_4_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa9_and1 = s_CSAwallace_rca24_csa1_csa_component_fa9_xor0 & s_CSAwallace_rca24_and_4_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa9_or0 = s_CSAwallace_rca24_csa1_csa_component_fa9_and0 | s_CSAwallace_rca24_csa1_csa_component_fa9_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa10_xor0 = s_CSAwallace_rca24_and_7_3 ^ s_CSAwallace_rca24_and_6_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa10_and0 = s_CSAwallace_rca24_and_7_3 & s_CSAwallace_rca24_and_6_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa10_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_and_5_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa10_and1 = s_CSAwallace_rca24_csa1_csa_component_fa10_xor0 & s_CSAwallace_rca24_and_5_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa10_or0 = s_CSAwallace_rca24_csa1_csa_component_fa10_and0 | s_CSAwallace_rca24_csa1_csa_component_fa10_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa11_xor0 = s_CSAwallace_rca24_and_8_3 ^ s_CSAwallace_rca24_and_7_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa11_and0 = s_CSAwallace_rca24_and_8_3 & s_CSAwallace_rca24_and_7_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa11_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_and_6_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa11_and1 = s_CSAwallace_rca24_csa1_csa_component_fa11_xor0 & s_CSAwallace_rca24_and_6_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa11_or0 = s_CSAwallace_rca24_csa1_csa_component_fa11_and0 | s_CSAwallace_rca24_csa1_csa_component_fa11_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa12_xor0 = s_CSAwallace_rca24_and_9_3 ^ s_CSAwallace_rca24_and_8_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa12_and0 = s_CSAwallace_rca24_and_9_3 & s_CSAwallace_rca24_and_8_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_and_7_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa12_and1 = s_CSAwallace_rca24_csa1_csa_component_fa12_xor0 & s_CSAwallace_rca24_and_7_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa12_or0 = s_CSAwallace_rca24_csa1_csa_component_fa12_and0 | s_CSAwallace_rca24_csa1_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa13_xor0 = s_CSAwallace_rca24_and_10_3 ^ s_CSAwallace_rca24_and_9_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa13_and0 = s_CSAwallace_rca24_and_10_3 & s_CSAwallace_rca24_and_9_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_and_8_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa13_and1 = s_CSAwallace_rca24_csa1_csa_component_fa13_xor0 & s_CSAwallace_rca24_and_8_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa13_or0 = s_CSAwallace_rca24_csa1_csa_component_fa13_and0 | s_CSAwallace_rca24_csa1_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa14_xor0 = s_CSAwallace_rca24_and_11_3 ^ s_CSAwallace_rca24_and_10_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa14_and0 = s_CSAwallace_rca24_and_11_3 & s_CSAwallace_rca24_and_10_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_and_9_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa14_and1 = s_CSAwallace_rca24_csa1_csa_component_fa14_xor0 & s_CSAwallace_rca24_and_9_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa14_or0 = s_CSAwallace_rca24_csa1_csa_component_fa14_and0 | s_CSAwallace_rca24_csa1_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa15_xor0 = s_CSAwallace_rca24_and_12_3 ^ s_CSAwallace_rca24_and_11_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa15_and0 = s_CSAwallace_rca24_and_12_3 & s_CSAwallace_rca24_and_11_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_and_10_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa15_and1 = s_CSAwallace_rca24_csa1_csa_component_fa15_xor0 & s_CSAwallace_rca24_and_10_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa15_or0 = s_CSAwallace_rca24_csa1_csa_component_fa15_and0 | s_CSAwallace_rca24_csa1_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa16_xor0 = s_CSAwallace_rca24_and_13_3 ^ s_CSAwallace_rca24_and_12_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa16_and0 = s_CSAwallace_rca24_and_13_3 & s_CSAwallace_rca24_and_12_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_and_11_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa16_and1 = s_CSAwallace_rca24_csa1_csa_component_fa16_xor0 & s_CSAwallace_rca24_and_11_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa16_or0 = s_CSAwallace_rca24_csa1_csa_component_fa16_and0 | s_CSAwallace_rca24_csa1_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa17_xor0 = s_CSAwallace_rca24_and_14_3 ^ s_CSAwallace_rca24_and_13_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa17_and0 = s_CSAwallace_rca24_and_14_3 & s_CSAwallace_rca24_and_13_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_and_12_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa17_and1 = s_CSAwallace_rca24_csa1_csa_component_fa17_xor0 & s_CSAwallace_rca24_and_12_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa17_or0 = s_CSAwallace_rca24_csa1_csa_component_fa17_and0 | s_CSAwallace_rca24_csa1_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa18_xor0 = s_CSAwallace_rca24_and_15_3 ^ s_CSAwallace_rca24_and_14_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa18_and0 = s_CSAwallace_rca24_and_15_3 & s_CSAwallace_rca24_and_14_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_and_13_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa18_and1 = s_CSAwallace_rca24_csa1_csa_component_fa18_xor0 & s_CSAwallace_rca24_and_13_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa18_or0 = s_CSAwallace_rca24_csa1_csa_component_fa18_and0 | s_CSAwallace_rca24_csa1_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa19_xor0 = s_CSAwallace_rca24_and_16_3 ^ s_CSAwallace_rca24_and_15_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa19_and0 = s_CSAwallace_rca24_and_16_3 & s_CSAwallace_rca24_and_15_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_and_14_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa19_and1 = s_CSAwallace_rca24_csa1_csa_component_fa19_xor0 & s_CSAwallace_rca24_and_14_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa19_or0 = s_CSAwallace_rca24_csa1_csa_component_fa19_and0 | s_CSAwallace_rca24_csa1_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa20_xor0 = s_CSAwallace_rca24_and_17_3 ^ s_CSAwallace_rca24_and_16_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa20_and0 = s_CSAwallace_rca24_and_17_3 & s_CSAwallace_rca24_and_16_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_and_15_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa20_and1 = s_CSAwallace_rca24_csa1_csa_component_fa20_xor0 & s_CSAwallace_rca24_and_15_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa20_or0 = s_CSAwallace_rca24_csa1_csa_component_fa20_and0 | s_CSAwallace_rca24_csa1_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa21_xor0 = s_CSAwallace_rca24_and_18_3 ^ s_CSAwallace_rca24_and_17_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa21_and0 = s_CSAwallace_rca24_and_18_3 & s_CSAwallace_rca24_and_17_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_and_16_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa21_and1 = s_CSAwallace_rca24_csa1_csa_component_fa21_xor0 & s_CSAwallace_rca24_and_16_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa21_or0 = s_CSAwallace_rca24_csa1_csa_component_fa21_and0 | s_CSAwallace_rca24_csa1_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa22_xor0 = s_CSAwallace_rca24_and_19_3 ^ s_CSAwallace_rca24_and_18_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa22_and0 = s_CSAwallace_rca24_and_19_3 & s_CSAwallace_rca24_and_18_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_and_17_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa22_and1 = s_CSAwallace_rca24_csa1_csa_component_fa22_xor0 & s_CSAwallace_rca24_and_17_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa22_or0 = s_CSAwallace_rca24_csa1_csa_component_fa22_and0 | s_CSAwallace_rca24_csa1_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa23_xor0 = s_CSAwallace_rca24_and_20_3 ^ s_CSAwallace_rca24_and_19_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa23_and0 = s_CSAwallace_rca24_and_20_3 & s_CSAwallace_rca24_and_19_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_and_18_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa23_and1 = s_CSAwallace_rca24_csa1_csa_component_fa23_xor0 & s_CSAwallace_rca24_and_18_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa23_or0 = s_CSAwallace_rca24_csa1_csa_component_fa23_and0 | s_CSAwallace_rca24_csa1_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa24_xor0 = s_CSAwallace_rca24_and_21_3 ^ s_CSAwallace_rca24_and_20_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa24_and0 = s_CSAwallace_rca24_and_21_3 & s_CSAwallace_rca24_and_20_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_and_19_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa24_and1 = s_CSAwallace_rca24_csa1_csa_component_fa24_xor0 & s_CSAwallace_rca24_and_19_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa24_or0 = s_CSAwallace_rca24_csa1_csa_component_fa24_and0 | s_CSAwallace_rca24_csa1_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa25_xor0 = s_CSAwallace_rca24_and_22_3 ^ s_CSAwallace_rca24_and_21_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa25_and0 = s_CSAwallace_rca24_and_22_3 & s_CSAwallace_rca24_and_21_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_and_20_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa25_and1 = s_CSAwallace_rca24_csa1_csa_component_fa25_xor0 & s_CSAwallace_rca24_and_20_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa25_or0 = s_CSAwallace_rca24_csa1_csa_component_fa25_and0 | s_CSAwallace_rca24_csa1_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa26_xor0 = s_CSAwallace_rca24_nand_23_3 ^ s_CSAwallace_rca24_and_22_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa26_and0 = s_CSAwallace_rca24_nand_23_3 & s_CSAwallace_rca24_and_22_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_and_21_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa26_and1 = s_CSAwallace_rca24_csa1_csa_component_fa26_xor0 & s_CSAwallace_rca24_and_21_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa26_or0 = s_CSAwallace_rca24_csa1_csa_component_fa26_and0 | s_CSAwallace_rca24_csa1_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa1_csa_component_fa27_xor0 = ~s_CSAwallace_rca24_nand_23_4;
  assign s_CSAwallace_rca24_csa1_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa1_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_and_22_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa27_and1 = s_CSAwallace_rca24_csa1_csa_component_fa27_xor0 & s_CSAwallace_rca24_and_22_5;
  assign s_CSAwallace_rca24_csa1_csa_component_fa27_or0 = s_CSAwallace_rca24_nand_23_4 | s_CSAwallace_rca24_csa1_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa7_xor0 = s_CSAwallace_rca24_and_1_6 ^ s_CSAwallace_rca24_and_0_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa7_and0 = s_CSAwallace_rca24_and_1_6 & s_CSAwallace_rca24_and_0_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa8_xor0 = s_CSAwallace_rca24_and_2_6 ^ s_CSAwallace_rca24_and_1_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa8_and0 = s_CSAwallace_rca24_and_2_6 & s_CSAwallace_rca24_and_1_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa8_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_and_0_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa8_and1 = s_CSAwallace_rca24_csa2_csa_component_fa8_xor0 & s_CSAwallace_rca24_and_0_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa8_or0 = s_CSAwallace_rca24_csa2_csa_component_fa8_and0 | s_CSAwallace_rca24_csa2_csa_component_fa8_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa9_xor0 = s_CSAwallace_rca24_and_3_6 ^ s_CSAwallace_rca24_and_2_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa9_and0 = s_CSAwallace_rca24_and_3_6 & s_CSAwallace_rca24_and_2_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa9_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_and_1_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa9_and1 = s_CSAwallace_rca24_csa2_csa_component_fa9_xor0 & s_CSAwallace_rca24_and_1_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa9_or0 = s_CSAwallace_rca24_csa2_csa_component_fa9_and0 | s_CSAwallace_rca24_csa2_csa_component_fa9_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa10_xor0 = s_CSAwallace_rca24_and_4_6 ^ s_CSAwallace_rca24_and_3_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa10_and0 = s_CSAwallace_rca24_and_4_6 & s_CSAwallace_rca24_and_3_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa10_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_and_2_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa10_and1 = s_CSAwallace_rca24_csa2_csa_component_fa10_xor0 & s_CSAwallace_rca24_and_2_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa10_or0 = s_CSAwallace_rca24_csa2_csa_component_fa10_and0 | s_CSAwallace_rca24_csa2_csa_component_fa10_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa11_xor0 = s_CSAwallace_rca24_and_5_6 ^ s_CSAwallace_rca24_and_4_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa11_and0 = s_CSAwallace_rca24_and_5_6 & s_CSAwallace_rca24_and_4_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa11_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_and_3_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa11_and1 = s_CSAwallace_rca24_csa2_csa_component_fa11_xor0 & s_CSAwallace_rca24_and_3_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa11_or0 = s_CSAwallace_rca24_csa2_csa_component_fa11_and0 | s_CSAwallace_rca24_csa2_csa_component_fa11_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa12_xor0 = s_CSAwallace_rca24_and_6_6 ^ s_CSAwallace_rca24_and_5_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa12_and0 = s_CSAwallace_rca24_and_6_6 & s_CSAwallace_rca24_and_5_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_and_4_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa12_and1 = s_CSAwallace_rca24_csa2_csa_component_fa12_xor0 & s_CSAwallace_rca24_and_4_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa12_or0 = s_CSAwallace_rca24_csa2_csa_component_fa12_and0 | s_CSAwallace_rca24_csa2_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa13_xor0 = s_CSAwallace_rca24_and_7_6 ^ s_CSAwallace_rca24_and_6_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa13_and0 = s_CSAwallace_rca24_and_7_6 & s_CSAwallace_rca24_and_6_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_and_5_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa13_and1 = s_CSAwallace_rca24_csa2_csa_component_fa13_xor0 & s_CSAwallace_rca24_and_5_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa13_or0 = s_CSAwallace_rca24_csa2_csa_component_fa13_and0 | s_CSAwallace_rca24_csa2_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa14_xor0 = s_CSAwallace_rca24_and_8_6 ^ s_CSAwallace_rca24_and_7_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa14_and0 = s_CSAwallace_rca24_and_8_6 & s_CSAwallace_rca24_and_7_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_and_6_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa14_and1 = s_CSAwallace_rca24_csa2_csa_component_fa14_xor0 & s_CSAwallace_rca24_and_6_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa14_or0 = s_CSAwallace_rca24_csa2_csa_component_fa14_and0 | s_CSAwallace_rca24_csa2_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa15_xor0 = s_CSAwallace_rca24_and_9_6 ^ s_CSAwallace_rca24_and_8_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa15_and0 = s_CSAwallace_rca24_and_9_6 & s_CSAwallace_rca24_and_8_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_and_7_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa15_and1 = s_CSAwallace_rca24_csa2_csa_component_fa15_xor0 & s_CSAwallace_rca24_and_7_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa15_or0 = s_CSAwallace_rca24_csa2_csa_component_fa15_and0 | s_CSAwallace_rca24_csa2_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa16_xor0 = s_CSAwallace_rca24_and_10_6 ^ s_CSAwallace_rca24_and_9_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa16_and0 = s_CSAwallace_rca24_and_10_6 & s_CSAwallace_rca24_and_9_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_and_8_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa16_and1 = s_CSAwallace_rca24_csa2_csa_component_fa16_xor0 & s_CSAwallace_rca24_and_8_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa16_or0 = s_CSAwallace_rca24_csa2_csa_component_fa16_and0 | s_CSAwallace_rca24_csa2_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa17_xor0 = s_CSAwallace_rca24_and_11_6 ^ s_CSAwallace_rca24_and_10_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa17_and0 = s_CSAwallace_rca24_and_11_6 & s_CSAwallace_rca24_and_10_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_and_9_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa17_and1 = s_CSAwallace_rca24_csa2_csa_component_fa17_xor0 & s_CSAwallace_rca24_and_9_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa17_or0 = s_CSAwallace_rca24_csa2_csa_component_fa17_and0 | s_CSAwallace_rca24_csa2_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa18_xor0 = s_CSAwallace_rca24_and_12_6 ^ s_CSAwallace_rca24_and_11_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa18_and0 = s_CSAwallace_rca24_and_12_6 & s_CSAwallace_rca24_and_11_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_and_10_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa18_and1 = s_CSAwallace_rca24_csa2_csa_component_fa18_xor0 & s_CSAwallace_rca24_and_10_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa18_or0 = s_CSAwallace_rca24_csa2_csa_component_fa18_and0 | s_CSAwallace_rca24_csa2_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa19_xor0 = s_CSAwallace_rca24_and_13_6 ^ s_CSAwallace_rca24_and_12_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa19_and0 = s_CSAwallace_rca24_and_13_6 & s_CSAwallace_rca24_and_12_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_and_11_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa19_and1 = s_CSAwallace_rca24_csa2_csa_component_fa19_xor0 & s_CSAwallace_rca24_and_11_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa19_or0 = s_CSAwallace_rca24_csa2_csa_component_fa19_and0 | s_CSAwallace_rca24_csa2_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa20_xor0 = s_CSAwallace_rca24_and_14_6 ^ s_CSAwallace_rca24_and_13_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa20_and0 = s_CSAwallace_rca24_and_14_6 & s_CSAwallace_rca24_and_13_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_and_12_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa20_and1 = s_CSAwallace_rca24_csa2_csa_component_fa20_xor0 & s_CSAwallace_rca24_and_12_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa20_or0 = s_CSAwallace_rca24_csa2_csa_component_fa20_and0 | s_CSAwallace_rca24_csa2_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa21_xor0 = s_CSAwallace_rca24_and_15_6 ^ s_CSAwallace_rca24_and_14_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa21_and0 = s_CSAwallace_rca24_and_15_6 & s_CSAwallace_rca24_and_14_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_and_13_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa21_and1 = s_CSAwallace_rca24_csa2_csa_component_fa21_xor0 & s_CSAwallace_rca24_and_13_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa21_or0 = s_CSAwallace_rca24_csa2_csa_component_fa21_and0 | s_CSAwallace_rca24_csa2_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa22_xor0 = s_CSAwallace_rca24_and_16_6 ^ s_CSAwallace_rca24_and_15_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa22_and0 = s_CSAwallace_rca24_and_16_6 & s_CSAwallace_rca24_and_15_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_and_14_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa22_and1 = s_CSAwallace_rca24_csa2_csa_component_fa22_xor0 & s_CSAwallace_rca24_and_14_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa22_or0 = s_CSAwallace_rca24_csa2_csa_component_fa22_and0 | s_CSAwallace_rca24_csa2_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa23_xor0 = s_CSAwallace_rca24_and_17_6 ^ s_CSAwallace_rca24_and_16_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa23_and0 = s_CSAwallace_rca24_and_17_6 & s_CSAwallace_rca24_and_16_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_and_15_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa23_and1 = s_CSAwallace_rca24_csa2_csa_component_fa23_xor0 & s_CSAwallace_rca24_and_15_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa23_or0 = s_CSAwallace_rca24_csa2_csa_component_fa23_and0 | s_CSAwallace_rca24_csa2_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa24_xor0 = s_CSAwallace_rca24_and_18_6 ^ s_CSAwallace_rca24_and_17_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa24_and0 = s_CSAwallace_rca24_and_18_6 & s_CSAwallace_rca24_and_17_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_and_16_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa24_and1 = s_CSAwallace_rca24_csa2_csa_component_fa24_xor0 & s_CSAwallace_rca24_and_16_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa24_or0 = s_CSAwallace_rca24_csa2_csa_component_fa24_and0 | s_CSAwallace_rca24_csa2_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa25_xor0 = s_CSAwallace_rca24_and_19_6 ^ s_CSAwallace_rca24_and_18_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa25_and0 = s_CSAwallace_rca24_and_19_6 & s_CSAwallace_rca24_and_18_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_and_17_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa25_and1 = s_CSAwallace_rca24_csa2_csa_component_fa25_xor0 & s_CSAwallace_rca24_and_17_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa25_or0 = s_CSAwallace_rca24_csa2_csa_component_fa25_and0 | s_CSAwallace_rca24_csa2_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa26_xor0 = s_CSAwallace_rca24_and_20_6 ^ s_CSAwallace_rca24_and_19_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa26_and0 = s_CSAwallace_rca24_and_20_6 & s_CSAwallace_rca24_and_19_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_and_18_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa26_and1 = s_CSAwallace_rca24_csa2_csa_component_fa26_xor0 & s_CSAwallace_rca24_and_18_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa26_or0 = s_CSAwallace_rca24_csa2_csa_component_fa26_and0 | s_CSAwallace_rca24_csa2_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa27_xor0 = s_CSAwallace_rca24_and_21_6 ^ s_CSAwallace_rca24_and_20_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa27_and0 = s_CSAwallace_rca24_and_21_6 & s_CSAwallace_rca24_and_20_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_and_19_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa27_and1 = s_CSAwallace_rca24_csa2_csa_component_fa27_xor0 & s_CSAwallace_rca24_and_19_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa27_or0 = s_CSAwallace_rca24_csa2_csa_component_fa27_and0 | s_CSAwallace_rca24_csa2_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa28_xor0 = s_CSAwallace_rca24_and_22_6 ^ s_CSAwallace_rca24_and_21_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa28_and0 = s_CSAwallace_rca24_and_22_6 & s_CSAwallace_rca24_and_21_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_and_20_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa28_and1 = s_CSAwallace_rca24_csa2_csa_component_fa28_xor0 & s_CSAwallace_rca24_and_20_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa28_or0 = s_CSAwallace_rca24_csa2_csa_component_fa28_and0 | s_CSAwallace_rca24_csa2_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa29_xor0 = s_CSAwallace_rca24_nand_23_6 ^ s_CSAwallace_rca24_and_22_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa29_and0 = s_CSAwallace_rca24_nand_23_6 & s_CSAwallace_rca24_and_22_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_and_21_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa29_and1 = s_CSAwallace_rca24_csa2_csa_component_fa29_xor0 & s_CSAwallace_rca24_and_21_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa29_or0 = s_CSAwallace_rca24_csa2_csa_component_fa29_and0 | s_CSAwallace_rca24_csa2_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa2_csa_component_fa30_xor0 = ~s_CSAwallace_rca24_nand_23_7;
  assign s_CSAwallace_rca24_csa2_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa2_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_and_22_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa30_and1 = s_CSAwallace_rca24_csa2_csa_component_fa30_xor0 & s_CSAwallace_rca24_and_22_8;
  assign s_CSAwallace_rca24_csa2_csa_component_fa30_or0 = s_CSAwallace_rca24_nand_23_7 | s_CSAwallace_rca24_csa2_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa10_xor0 = s_CSAwallace_rca24_and_1_9 ^ s_CSAwallace_rca24_and_0_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa10_and0 = s_CSAwallace_rca24_and_1_9 & s_CSAwallace_rca24_and_0_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa11_xor0 = s_CSAwallace_rca24_and_2_9 ^ s_CSAwallace_rca24_and_1_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa11_and0 = s_CSAwallace_rca24_and_2_9 & s_CSAwallace_rca24_and_1_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa11_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_and_0_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa11_and1 = s_CSAwallace_rca24_csa3_csa_component_fa11_xor0 & s_CSAwallace_rca24_and_0_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa11_or0 = s_CSAwallace_rca24_csa3_csa_component_fa11_and0 | s_CSAwallace_rca24_csa3_csa_component_fa11_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa12_xor0 = s_CSAwallace_rca24_and_3_9 ^ s_CSAwallace_rca24_and_2_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa12_and0 = s_CSAwallace_rca24_and_3_9 & s_CSAwallace_rca24_and_2_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_and_1_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa12_and1 = s_CSAwallace_rca24_csa3_csa_component_fa12_xor0 & s_CSAwallace_rca24_and_1_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa12_or0 = s_CSAwallace_rca24_csa3_csa_component_fa12_and0 | s_CSAwallace_rca24_csa3_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa13_xor0 = s_CSAwallace_rca24_and_4_9 ^ s_CSAwallace_rca24_and_3_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa13_and0 = s_CSAwallace_rca24_and_4_9 & s_CSAwallace_rca24_and_3_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_and_2_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa13_and1 = s_CSAwallace_rca24_csa3_csa_component_fa13_xor0 & s_CSAwallace_rca24_and_2_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa13_or0 = s_CSAwallace_rca24_csa3_csa_component_fa13_and0 | s_CSAwallace_rca24_csa3_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa14_xor0 = s_CSAwallace_rca24_and_5_9 ^ s_CSAwallace_rca24_and_4_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa14_and0 = s_CSAwallace_rca24_and_5_9 & s_CSAwallace_rca24_and_4_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_and_3_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa14_and1 = s_CSAwallace_rca24_csa3_csa_component_fa14_xor0 & s_CSAwallace_rca24_and_3_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa14_or0 = s_CSAwallace_rca24_csa3_csa_component_fa14_and0 | s_CSAwallace_rca24_csa3_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa15_xor0 = s_CSAwallace_rca24_and_6_9 ^ s_CSAwallace_rca24_and_5_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa15_and0 = s_CSAwallace_rca24_and_6_9 & s_CSAwallace_rca24_and_5_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_and_4_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa15_and1 = s_CSAwallace_rca24_csa3_csa_component_fa15_xor0 & s_CSAwallace_rca24_and_4_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa15_or0 = s_CSAwallace_rca24_csa3_csa_component_fa15_and0 | s_CSAwallace_rca24_csa3_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa16_xor0 = s_CSAwallace_rca24_and_7_9 ^ s_CSAwallace_rca24_and_6_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa16_and0 = s_CSAwallace_rca24_and_7_9 & s_CSAwallace_rca24_and_6_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_and_5_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa16_and1 = s_CSAwallace_rca24_csa3_csa_component_fa16_xor0 & s_CSAwallace_rca24_and_5_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa16_or0 = s_CSAwallace_rca24_csa3_csa_component_fa16_and0 | s_CSAwallace_rca24_csa3_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa17_xor0 = s_CSAwallace_rca24_and_8_9 ^ s_CSAwallace_rca24_and_7_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa17_and0 = s_CSAwallace_rca24_and_8_9 & s_CSAwallace_rca24_and_7_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_and_6_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa17_and1 = s_CSAwallace_rca24_csa3_csa_component_fa17_xor0 & s_CSAwallace_rca24_and_6_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa17_or0 = s_CSAwallace_rca24_csa3_csa_component_fa17_and0 | s_CSAwallace_rca24_csa3_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa18_xor0 = s_CSAwallace_rca24_and_9_9 ^ s_CSAwallace_rca24_and_8_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa18_and0 = s_CSAwallace_rca24_and_9_9 & s_CSAwallace_rca24_and_8_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_and_7_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa18_and1 = s_CSAwallace_rca24_csa3_csa_component_fa18_xor0 & s_CSAwallace_rca24_and_7_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa18_or0 = s_CSAwallace_rca24_csa3_csa_component_fa18_and0 | s_CSAwallace_rca24_csa3_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa19_xor0 = s_CSAwallace_rca24_and_10_9 ^ s_CSAwallace_rca24_and_9_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa19_and0 = s_CSAwallace_rca24_and_10_9 & s_CSAwallace_rca24_and_9_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_and_8_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa19_and1 = s_CSAwallace_rca24_csa3_csa_component_fa19_xor0 & s_CSAwallace_rca24_and_8_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa19_or0 = s_CSAwallace_rca24_csa3_csa_component_fa19_and0 | s_CSAwallace_rca24_csa3_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa20_xor0 = s_CSAwallace_rca24_and_11_9 ^ s_CSAwallace_rca24_and_10_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa20_and0 = s_CSAwallace_rca24_and_11_9 & s_CSAwallace_rca24_and_10_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_and_9_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa20_and1 = s_CSAwallace_rca24_csa3_csa_component_fa20_xor0 & s_CSAwallace_rca24_and_9_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa20_or0 = s_CSAwallace_rca24_csa3_csa_component_fa20_and0 | s_CSAwallace_rca24_csa3_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa21_xor0 = s_CSAwallace_rca24_and_12_9 ^ s_CSAwallace_rca24_and_11_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa21_and0 = s_CSAwallace_rca24_and_12_9 & s_CSAwallace_rca24_and_11_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_and_10_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa21_and1 = s_CSAwallace_rca24_csa3_csa_component_fa21_xor0 & s_CSAwallace_rca24_and_10_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa21_or0 = s_CSAwallace_rca24_csa3_csa_component_fa21_and0 | s_CSAwallace_rca24_csa3_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa22_xor0 = s_CSAwallace_rca24_and_13_9 ^ s_CSAwallace_rca24_and_12_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa22_and0 = s_CSAwallace_rca24_and_13_9 & s_CSAwallace_rca24_and_12_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_and_11_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa22_and1 = s_CSAwallace_rca24_csa3_csa_component_fa22_xor0 & s_CSAwallace_rca24_and_11_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa22_or0 = s_CSAwallace_rca24_csa3_csa_component_fa22_and0 | s_CSAwallace_rca24_csa3_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa23_xor0 = s_CSAwallace_rca24_and_14_9 ^ s_CSAwallace_rca24_and_13_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa23_and0 = s_CSAwallace_rca24_and_14_9 & s_CSAwallace_rca24_and_13_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_and_12_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa23_and1 = s_CSAwallace_rca24_csa3_csa_component_fa23_xor0 & s_CSAwallace_rca24_and_12_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa23_or0 = s_CSAwallace_rca24_csa3_csa_component_fa23_and0 | s_CSAwallace_rca24_csa3_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa24_xor0 = s_CSAwallace_rca24_and_15_9 ^ s_CSAwallace_rca24_and_14_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa24_and0 = s_CSAwallace_rca24_and_15_9 & s_CSAwallace_rca24_and_14_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_and_13_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa24_and1 = s_CSAwallace_rca24_csa3_csa_component_fa24_xor0 & s_CSAwallace_rca24_and_13_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa24_or0 = s_CSAwallace_rca24_csa3_csa_component_fa24_and0 | s_CSAwallace_rca24_csa3_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa25_xor0 = s_CSAwallace_rca24_and_16_9 ^ s_CSAwallace_rca24_and_15_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa25_and0 = s_CSAwallace_rca24_and_16_9 & s_CSAwallace_rca24_and_15_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_and_14_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa25_and1 = s_CSAwallace_rca24_csa3_csa_component_fa25_xor0 & s_CSAwallace_rca24_and_14_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa25_or0 = s_CSAwallace_rca24_csa3_csa_component_fa25_and0 | s_CSAwallace_rca24_csa3_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa26_xor0 = s_CSAwallace_rca24_and_17_9 ^ s_CSAwallace_rca24_and_16_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa26_and0 = s_CSAwallace_rca24_and_17_9 & s_CSAwallace_rca24_and_16_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_and_15_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa26_and1 = s_CSAwallace_rca24_csa3_csa_component_fa26_xor0 & s_CSAwallace_rca24_and_15_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa26_or0 = s_CSAwallace_rca24_csa3_csa_component_fa26_and0 | s_CSAwallace_rca24_csa3_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa27_xor0 = s_CSAwallace_rca24_and_18_9 ^ s_CSAwallace_rca24_and_17_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa27_and0 = s_CSAwallace_rca24_and_18_9 & s_CSAwallace_rca24_and_17_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_and_16_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa27_and1 = s_CSAwallace_rca24_csa3_csa_component_fa27_xor0 & s_CSAwallace_rca24_and_16_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa27_or0 = s_CSAwallace_rca24_csa3_csa_component_fa27_and0 | s_CSAwallace_rca24_csa3_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa28_xor0 = s_CSAwallace_rca24_and_19_9 ^ s_CSAwallace_rca24_and_18_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa28_and0 = s_CSAwallace_rca24_and_19_9 & s_CSAwallace_rca24_and_18_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_and_17_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa28_and1 = s_CSAwallace_rca24_csa3_csa_component_fa28_xor0 & s_CSAwallace_rca24_and_17_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa28_or0 = s_CSAwallace_rca24_csa3_csa_component_fa28_and0 | s_CSAwallace_rca24_csa3_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa29_xor0 = s_CSAwallace_rca24_and_20_9 ^ s_CSAwallace_rca24_and_19_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa29_and0 = s_CSAwallace_rca24_and_20_9 & s_CSAwallace_rca24_and_19_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_and_18_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa29_and1 = s_CSAwallace_rca24_csa3_csa_component_fa29_xor0 & s_CSAwallace_rca24_and_18_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa29_or0 = s_CSAwallace_rca24_csa3_csa_component_fa29_and0 | s_CSAwallace_rca24_csa3_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa30_xor0 = s_CSAwallace_rca24_and_21_9 ^ s_CSAwallace_rca24_and_20_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa30_and0 = s_CSAwallace_rca24_and_21_9 & s_CSAwallace_rca24_and_20_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_and_19_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa30_and1 = s_CSAwallace_rca24_csa3_csa_component_fa30_xor0 & s_CSAwallace_rca24_and_19_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa30_or0 = s_CSAwallace_rca24_csa3_csa_component_fa30_and0 | s_CSAwallace_rca24_csa3_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa31_xor0 = s_CSAwallace_rca24_and_22_9 ^ s_CSAwallace_rca24_and_21_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa31_and0 = s_CSAwallace_rca24_and_22_9 & s_CSAwallace_rca24_and_21_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_and_20_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa31_and1 = s_CSAwallace_rca24_csa3_csa_component_fa31_xor0 & s_CSAwallace_rca24_and_20_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa31_or0 = s_CSAwallace_rca24_csa3_csa_component_fa31_and0 | s_CSAwallace_rca24_csa3_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa32_xor0 = s_CSAwallace_rca24_nand_23_9 ^ s_CSAwallace_rca24_and_22_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa32_and0 = s_CSAwallace_rca24_nand_23_9 & s_CSAwallace_rca24_and_22_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_and_21_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa32_and1 = s_CSAwallace_rca24_csa3_csa_component_fa32_xor0 & s_CSAwallace_rca24_and_21_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa32_or0 = s_CSAwallace_rca24_csa3_csa_component_fa32_and0 | s_CSAwallace_rca24_csa3_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa3_csa_component_fa33_xor0 = ~s_CSAwallace_rca24_nand_23_10;
  assign s_CSAwallace_rca24_csa3_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa3_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_and_22_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa33_and1 = s_CSAwallace_rca24_csa3_csa_component_fa33_xor0 & s_CSAwallace_rca24_and_22_11;
  assign s_CSAwallace_rca24_csa3_csa_component_fa33_or0 = s_CSAwallace_rca24_nand_23_10 | s_CSAwallace_rca24_csa3_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa13_xor0 = s_CSAwallace_rca24_and_1_12 ^ s_CSAwallace_rca24_and_0_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa13_and0 = s_CSAwallace_rca24_and_1_12 & s_CSAwallace_rca24_and_0_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa14_xor0 = s_CSAwallace_rca24_and_2_12 ^ s_CSAwallace_rca24_and_1_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa14_and0 = s_CSAwallace_rca24_and_2_12 & s_CSAwallace_rca24_and_1_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_and_0_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa14_and1 = s_CSAwallace_rca24_csa4_csa_component_fa14_xor0 & s_CSAwallace_rca24_and_0_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa14_or0 = s_CSAwallace_rca24_csa4_csa_component_fa14_and0 | s_CSAwallace_rca24_csa4_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa15_xor0 = s_CSAwallace_rca24_and_3_12 ^ s_CSAwallace_rca24_and_2_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa15_and0 = s_CSAwallace_rca24_and_3_12 & s_CSAwallace_rca24_and_2_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_and_1_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa15_and1 = s_CSAwallace_rca24_csa4_csa_component_fa15_xor0 & s_CSAwallace_rca24_and_1_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa15_or0 = s_CSAwallace_rca24_csa4_csa_component_fa15_and0 | s_CSAwallace_rca24_csa4_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa16_xor0 = s_CSAwallace_rca24_and_4_12 ^ s_CSAwallace_rca24_and_3_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa16_and0 = s_CSAwallace_rca24_and_4_12 & s_CSAwallace_rca24_and_3_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_and_2_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa16_and1 = s_CSAwallace_rca24_csa4_csa_component_fa16_xor0 & s_CSAwallace_rca24_and_2_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa16_or0 = s_CSAwallace_rca24_csa4_csa_component_fa16_and0 | s_CSAwallace_rca24_csa4_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa17_xor0 = s_CSAwallace_rca24_and_5_12 ^ s_CSAwallace_rca24_and_4_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa17_and0 = s_CSAwallace_rca24_and_5_12 & s_CSAwallace_rca24_and_4_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_and_3_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa17_and1 = s_CSAwallace_rca24_csa4_csa_component_fa17_xor0 & s_CSAwallace_rca24_and_3_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa17_or0 = s_CSAwallace_rca24_csa4_csa_component_fa17_and0 | s_CSAwallace_rca24_csa4_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa18_xor0 = s_CSAwallace_rca24_and_6_12 ^ s_CSAwallace_rca24_and_5_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa18_and0 = s_CSAwallace_rca24_and_6_12 & s_CSAwallace_rca24_and_5_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_and_4_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa18_and1 = s_CSAwallace_rca24_csa4_csa_component_fa18_xor0 & s_CSAwallace_rca24_and_4_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa18_or0 = s_CSAwallace_rca24_csa4_csa_component_fa18_and0 | s_CSAwallace_rca24_csa4_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa19_xor0 = s_CSAwallace_rca24_and_7_12 ^ s_CSAwallace_rca24_and_6_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa19_and0 = s_CSAwallace_rca24_and_7_12 & s_CSAwallace_rca24_and_6_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_and_5_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa19_and1 = s_CSAwallace_rca24_csa4_csa_component_fa19_xor0 & s_CSAwallace_rca24_and_5_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa19_or0 = s_CSAwallace_rca24_csa4_csa_component_fa19_and0 | s_CSAwallace_rca24_csa4_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa20_xor0 = s_CSAwallace_rca24_and_8_12 ^ s_CSAwallace_rca24_and_7_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa20_and0 = s_CSAwallace_rca24_and_8_12 & s_CSAwallace_rca24_and_7_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_and_6_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa20_and1 = s_CSAwallace_rca24_csa4_csa_component_fa20_xor0 & s_CSAwallace_rca24_and_6_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa20_or0 = s_CSAwallace_rca24_csa4_csa_component_fa20_and0 | s_CSAwallace_rca24_csa4_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa21_xor0 = s_CSAwallace_rca24_and_9_12 ^ s_CSAwallace_rca24_and_8_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa21_and0 = s_CSAwallace_rca24_and_9_12 & s_CSAwallace_rca24_and_8_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_and_7_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa21_and1 = s_CSAwallace_rca24_csa4_csa_component_fa21_xor0 & s_CSAwallace_rca24_and_7_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa21_or0 = s_CSAwallace_rca24_csa4_csa_component_fa21_and0 | s_CSAwallace_rca24_csa4_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa22_xor0 = s_CSAwallace_rca24_and_10_12 ^ s_CSAwallace_rca24_and_9_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa22_and0 = s_CSAwallace_rca24_and_10_12 & s_CSAwallace_rca24_and_9_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_and_8_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa22_and1 = s_CSAwallace_rca24_csa4_csa_component_fa22_xor0 & s_CSAwallace_rca24_and_8_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa22_or0 = s_CSAwallace_rca24_csa4_csa_component_fa22_and0 | s_CSAwallace_rca24_csa4_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa23_xor0 = s_CSAwallace_rca24_and_11_12 ^ s_CSAwallace_rca24_and_10_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa23_and0 = s_CSAwallace_rca24_and_11_12 & s_CSAwallace_rca24_and_10_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_and_9_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa23_and1 = s_CSAwallace_rca24_csa4_csa_component_fa23_xor0 & s_CSAwallace_rca24_and_9_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa23_or0 = s_CSAwallace_rca24_csa4_csa_component_fa23_and0 | s_CSAwallace_rca24_csa4_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa24_xor0 = s_CSAwallace_rca24_and_12_12 ^ s_CSAwallace_rca24_and_11_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa24_and0 = s_CSAwallace_rca24_and_12_12 & s_CSAwallace_rca24_and_11_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_and_10_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa24_and1 = s_CSAwallace_rca24_csa4_csa_component_fa24_xor0 & s_CSAwallace_rca24_and_10_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa24_or0 = s_CSAwallace_rca24_csa4_csa_component_fa24_and0 | s_CSAwallace_rca24_csa4_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa25_xor0 = s_CSAwallace_rca24_and_13_12 ^ s_CSAwallace_rca24_and_12_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa25_and0 = s_CSAwallace_rca24_and_13_12 & s_CSAwallace_rca24_and_12_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_and_11_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa25_and1 = s_CSAwallace_rca24_csa4_csa_component_fa25_xor0 & s_CSAwallace_rca24_and_11_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa25_or0 = s_CSAwallace_rca24_csa4_csa_component_fa25_and0 | s_CSAwallace_rca24_csa4_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa26_xor0 = s_CSAwallace_rca24_and_14_12 ^ s_CSAwallace_rca24_and_13_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa26_and0 = s_CSAwallace_rca24_and_14_12 & s_CSAwallace_rca24_and_13_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_and_12_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa26_and1 = s_CSAwallace_rca24_csa4_csa_component_fa26_xor0 & s_CSAwallace_rca24_and_12_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa26_or0 = s_CSAwallace_rca24_csa4_csa_component_fa26_and0 | s_CSAwallace_rca24_csa4_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa27_xor0 = s_CSAwallace_rca24_and_15_12 ^ s_CSAwallace_rca24_and_14_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa27_and0 = s_CSAwallace_rca24_and_15_12 & s_CSAwallace_rca24_and_14_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_and_13_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa27_and1 = s_CSAwallace_rca24_csa4_csa_component_fa27_xor0 & s_CSAwallace_rca24_and_13_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa27_or0 = s_CSAwallace_rca24_csa4_csa_component_fa27_and0 | s_CSAwallace_rca24_csa4_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa28_xor0 = s_CSAwallace_rca24_and_16_12 ^ s_CSAwallace_rca24_and_15_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa28_and0 = s_CSAwallace_rca24_and_16_12 & s_CSAwallace_rca24_and_15_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_and_14_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa28_and1 = s_CSAwallace_rca24_csa4_csa_component_fa28_xor0 & s_CSAwallace_rca24_and_14_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa28_or0 = s_CSAwallace_rca24_csa4_csa_component_fa28_and0 | s_CSAwallace_rca24_csa4_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa29_xor0 = s_CSAwallace_rca24_and_17_12 ^ s_CSAwallace_rca24_and_16_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa29_and0 = s_CSAwallace_rca24_and_17_12 & s_CSAwallace_rca24_and_16_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_and_15_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa29_and1 = s_CSAwallace_rca24_csa4_csa_component_fa29_xor0 & s_CSAwallace_rca24_and_15_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa29_or0 = s_CSAwallace_rca24_csa4_csa_component_fa29_and0 | s_CSAwallace_rca24_csa4_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa30_xor0 = s_CSAwallace_rca24_and_18_12 ^ s_CSAwallace_rca24_and_17_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa30_and0 = s_CSAwallace_rca24_and_18_12 & s_CSAwallace_rca24_and_17_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_and_16_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa30_and1 = s_CSAwallace_rca24_csa4_csa_component_fa30_xor0 & s_CSAwallace_rca24_and_16_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa30_or0 = s_CSAwallace_rca24_csa4_csa_component_fa30_and0 | s_CSAwallace_rca24_csa4_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa31_xor0 = s_CSAwallace_rca24_and_19_12 ^ s_CSAwallace_rca24_and_18_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa31_and0 = s_CSAwallace_rca24_and_19_12 & s_CSAwallace_rca24_and_18_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_and_17_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa31_and1 = s_CSAwallace_rca24_csa4_csa_component_fa31_xor0 & s_CSAwallace_rca24_and_17_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa31_or0 = s_CSAwallace_rca24_csa4_csa_component_fa31_and0 | s_CSAwallace_rca24_csa4_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa32_xor0 = s_CSAwallace_rca24_and_20_12 ^ s_CSAwallace_rca24_and_19_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa32_and0 = s_CSAwallace_rca24_and_20_12 & s_CSAwallace_rca24_and_19_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_and_18_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa32_and1 = s_CSAwallace_rca24_csa4_csa_component_fa32_xor0 & s_CSAwallace_rca24_and_18_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa32_or0 = s_CSAwallace_rca24_csa4_csa_component_fa32_and0 | s_CSAwallace_rca24_csa4_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa33_xor0 = s_CSAwallace_rca24_and_21_12 ^ s_CSAwallace_rca24_and_20_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa33_and0 = s_CSAwallace_rca24_and_21_12 & s_CSAwallace_rca24_and_20_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_and_19_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa33_and1 = s_CSAwallace_rca24_csa4_csa_component_fa33_xor0 & s_CSAwallace_rca24_and_19_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa33_or0 = s_CSAwallace_rca24_csa4_csa_component_fa33_and0 | s_CSAwallace_rca24_csa4_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa34_xor0 = s_CSAwallace_rca24_and_22_12 ^ s_CSAwallace_rca24_and_21_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa34_and0 = s_CSAwallace_rca24_and_22_12 & s_CSAwallace_rca24_and_21_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_and_20_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa34_and1 = s_CSAwallace_rca24_csa4_csa_component_fa34_xor0 & s_CSAwallace_rca24_and_20_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa34_or0 = s_CSAwallace_rca24_csa4_csa_component_fa34_and0 | s_CSAwallace_rca24_csa4_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa35_xor0 = s_CSAwallace_rca24_nand_23_12 ^ s_CSAwallace_rca24_and_22_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa35_and0 = s_CSAwallace_rca24_nand_23_12 & s_CSAwallace_rca24_and_22_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_and_21_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa35_and1 = s_CSAwallace_rca24_csa4_csa_component_fa35_xor0 & s_CSAwallace_rca24_and_21_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa35_or0 = s_CSAwallace_rca24_csa4_csa_component_fa35_and0 | s_CSAwallace_rca24_csa4_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa4_csa_component_fa36_xor0 = ~s_CSAwallace_rca24_nand_23_13;
  assign s_CSAwallace_rca24_csa4_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa4_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_and_22_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa36_and1 = s_CSAwallace_rca24_csa4_csa_component_fa36_xor0 & s_CSAwallace_rca24_and_22_14;
  assign s_CSAwallace_rca24_csa4_csa_component_fa36_or0 = s_CSAwallace_rca24_nand_23_13 | s_CSAwallace_rca24_csa4_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa16_xor0 = s_CSAwallace_rca24_and_1_15 ^ s_CSAwallace_rca24_and_0_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa16_and0 = s_CSAwallace_rca24_and_1_15 & s_CSAwallace_rca24_and_0_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa17_xor0 = s_CSAwallace_rca24_and_2_15 ^ s_CSAwallace_rca24_and_1_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa17_and0 = s_CSAwallace_rca24_and_2_15 & s_CSAwallace_rca24_and_1_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_and_0_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa17_and1 = s_CSAwallace_rca24_csa5_csa_component_fa17_xor0 & s_CSAwallace_rca24_and_0_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa17_or0 = s_CSAwallace_rca24_csa5_csa_component_fa17_and0 | s_CSAwallace_rca24_csa5_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa18_xor0 = s_CSAwallace_rca24_and_3_15 ^ s_CSAwallace_rca24_and_2_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa18_and0 = s_CSAwallace_rca24_and_3_15 & s_CSAwallace_rca24_and_2_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_and_1_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa18_and1 = s_CSAwallace_rca24_csa5_csa_component_fa18_xor0 & s_CSAwallace_rca24_and_1_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa18_or0 = s_CSAwallace_rca24_csa5_csa_component_fa18_and0 | s_CSAwallace_rca24_csa5_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa19_xor0 = s_CSAwallace_rca24_and_4_15 ^ s_CSAwallace_rca24_and_3_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa19_and0 = s_CSAwallace_rca24_and_4_15 & s_CSAwallace_rca24_and_3_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_and_2_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa19_and1 = s_CSAwallace_rca24_csa5_csa_component_fa19_xor0 & s_CSAwallace_rca24_and_2_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa19_or0 = s_CSAwallace_rca24_csa5_csa_component_fa19_and0 | s_CSAwallace_rca24_csa5_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa20_xor0 = s_CSAwallace_rca24_and_5_15 ^ s_CSAwallace_rca24_and_4_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa20_and0 = s_CSAwallace_rca24_and_5_15 & s_CSAwallace_rca24_and_4_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_and_3_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa20_and1 = s_CSAwallace_rca24_csa5_csa_component_fa20_xor0 & s_CSAwallace_rca24_and_3_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa20_or0 = s_CSAwallace_rca24_csa5_csa_component_fa20_and0 | s_CSAwallace_rca24_csa5_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa21_xor0 = s_CSAwallace_rca24_and_6_15 ^ s_CSAwallace_rca24_and_5_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa21_and0 = s_CSAwallace_rca24_and_6_15 & s_CSAwallace_rca24_and_5_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_and_4_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa21_and1 = s_CSAwallace_rca24_csa5_csa_component_fa21_xor0 & s_CSAwallace_rca24_and_4_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa21_or0 = s_CSAwallace_rca24_csa5_csa_component_fa21_and0 | s_CSAwallace_rca24_csa5_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa22_xor0 = s_CSAwallace_rca24_and_7_15 ^ s_CSAwallace_rca24_and_6_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa22_and0 = s_CSAwallace_rca24_and_7_15 & s_CSAwallace_rca24_and_6_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_and_5_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa22_and1 = s_CSAwallace_rca24_csa5_csa_component_fa22_xor0 & s_CSAwallace_rca24_and_5_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa22_or0 = s_CSAwallace_rca24_csa5_csa_component_fa22_and0 | s_CSAwallace_rca24_csa5_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa23_xor0 = s_CSAwallace_rca24_and_8_15 ^ s_CSAwallace_rca24_and_7_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa23_and0 = s_CSAwallace_rca24_and_8_15 & s_CSAwallace_rca24_and_7_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_and_6_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa23_and1 = s_CSAwallace_rca24_csa5_csa_component_fa23_xor0 & s_CSAwallace_rca24_and_6_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa23_or0 = s_CSAwallace_rca24_csa5_csa_component_fa23_and0 | s_CSAwallace_rca24_csa5_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa24_xor0 = s_CSAwallace_rca24_and_9_15 ^ s_CSAwallace_rca24_and_8_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa24_and0 = s_CSAwallace_rca24_and_9_15 & s_CSAwallace_rca24_and_8_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_and_7_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa24_and1 = s_CSAwallace_rca24_csa5_csa_component_fa24_xor0 & s_CSAwallace_rca24_and_7_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa24_or0 = s_CSAwallace_rca24_csa5_csa_component_fa24_and0 | s_CSAwallace_rca24_csa5_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa25_xor0 = s_CSAwallace_rca24_and_10_15 ^ s_CSAwallace_rca24_and_9_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa25_and0 = s_CSAwallace_rca24_and_10_15 & s_CSAwallace_rca24_and_9_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_and_8_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa25_and1 = s_CSAwallace_rca24_csa5_csa_component_fa25_xor0 & s_CSAwallace_rca24_and_8_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa25_or0 = s_CSAwallace_rca24_csa5_csa_component_fa25_and0 | s_CSAwallace_rca24_csa5_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa26_xor0 = s_CSAwallace_rca24_and_11_15 ^ s_CSAwallace_rca24_and_10_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa26_and0 = s_CSAwallace_rca24_and_11_15 & s_CSAwallace_rca24_and_10_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_and_9_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa26_and1 = s_CSAwallace_rca24_csa5_csa_component_fa26_xor0 & s_CSAwallace_rca24_and_9_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa26_or0 = s_CSAwallace_rca24_csa5_csa_component_fa26_and0 | s_CSAwallace_rca24_csa5_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa27_xor0 = s_CSAwallace_rca24_and_12_15 ^ s_CSAwallace_rca24_and_11_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa27_and0 = s_CSAwallace_rca24_and_12_15 & s_CSAwallace_rca24_and_11_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_and_10_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa27_and1 = s_CSAwallace_rca24_csa5_csa_component_fa27_xor0 & s_CSAwallace_rca24_and_10_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa27_or0 = s_CSAwallace_rca24_csa5_csa_component_fa27_and0 | s_CSAwallace_rca24_csa5_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa28_xor0 = s_CSAwallace_rca24_and_13_15 ^ s_CSAwallace_rca24_and_12_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa28_and0 = s_CSAwallace_rca24_and_13_15 & s_CSAwallace_rca24_and_12_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_and_11_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa28_and1 = s_CSAwallace_rca24_csa5_csa_component_fa28_xor0 & s_CSAwallace_rca24_and_11_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa28_or0 = s_CSAwallace_rca24_csa5_csa_component_fa28_and0 | s_CSAwallace_rca24_csa5_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa29_xor0 = s_CSAwallace_rca24_and_14_15 ^ s_CSAwallace_rca24_and_13_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa29_and0 = s_CSAwallace_rca24_and_14_15 & s_CSAwallace_rca24_and_13_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_and_12_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa29_and1 = s_CSAwallace_rca24_csa5_csa_component_fa29_xor0 & s_CSAwallace_rca24_and_12_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa29_or0 = s_CSAwallace_rca24_csa5_csa_component_fa29_and0 | s_CSAwallace_rca24_csa5_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa30_xor0 = s_CSAwallace_rca24_and_15_15 ^ s_CSAwallace_rca24_and_14_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa30_and0 = s_CSAwallace_rca24_and_15_15 & s_CSAwallace_rca24_and_14_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_and_13_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa30_and1 = s_CSAwallace_rca24_csa5_csa_component_fa30_xor0 & s_CSAwallace_rca24_and_13_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa30_or0 = s_CSAwallace_rca24_csa5_csa_component_fa30_and0 | s_CSAwallace_rca24_csa5_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa31_xor0 = s_CSAwallace_rca24_and_16_15 ^ s_CSAwallace_rca24_and_15_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa31_and0 = s_CSAwallace_rca24_and_16_15 & s_CSAwallace_rca24_and_15_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_and_14_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa31_and1 = s_CSAwallace_rca24_csa5_csa_component_fa31_xor0 & s_CSAwallace_rca24_and_14_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa31_or0 = s_CSAwallace_rca24_csa5_csa_component_fa31_and0 | s_CSAwallace_rca24_csa5_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa32_xor0 = s_CSAwallace_rca24_and_17_15 ^ s_CSAwallace_rca24_and_16_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa32_and0 = s_CSAwallace_rca24_and_17_15 & s_CSAwallace_rca24_and_16_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_and_15_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa32_and1 = s_CSAwallace_rca24_csa5_csa_component_fa32_xor0 & s_CSAwallace_rca24_and_15_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa32_or0 = s_CSAwallace_rca24_csa5_csa_component_fa32_and0 | s_CSAwallace_rca24_csa5_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa33_xor0 = s_CSAwallace_rca24_and_18_15 ^ s_CSAwallace_rca24_and_17_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa33_and0 = s_CSAwallace_rca24_and_18_15 & s_CSAwallace_rca24_and_17_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_and_16_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa33_and1 = s_CSAwallace_rca24_csa5_csa_component_fa33_xor0 & s_CSAwallace_rca24_and_16_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa33_or0 = s_CSAwallace_rca24_csa5_csa_component_fa33_and0 | s_CSAwallace_rca24_csa5_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa34_xor0 = s_CSAwallace_rca24_and_19_15 ^ s_CSAwallace_rca24_and_18_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa34_and0 = s_CSAwallace_rca24_and_19_15 & s_CSAwallace_rca24_and_18_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_and_17_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa34_and1 = s_CSAwallace_rca24_csa5_csa_component_fa34_xor0 & s_CSAwallace_rca24_and_17_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa34_or0 = s_CSAwallace_rca24_csa5_csa_component_fa34_and0 | s_CSAwallace_rca24_csa5_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa35_xor0 = s_CSAwallace_rca24_and_20_15 ^ s_CSAwallace_rca24_and_19_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa35_and0 = s_CSAwallace_rca24_and_20_15 & s_CSAwallace_rca24_and_19_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_and_18_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa35_and1 = s_CSAwallace_rca24_csa5_csa_component_fa35_xor0 & s_CSAwallace_rca24_and_18_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa35_or0 = s_CSAwallace_rca24_csa5_csa_component_fa35_and0 | s_CSAwallace_rca24_csa5_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa36_xor0 = s_CSAwallace_rca24_and_21_15 ^ s_CSAwallace_rca24_and_20_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa36_and0 = s_CSAwallace_rca24_and_21_15 & s_CSAwallace_rca24_and_20_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_and_19_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa36_and1 = s_CSAwallace_rca24_csa5_csa_component_fa36_xor0 & s_CSAwallace_rca24_and_19_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa36_or0 = s_CSAwallace_rca24_csa5_csa_component_fa36_and0 | s_CSAwallace_rca24_csa5_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa37_xor0 = s_CSAwallace_rca24_and_22_15 ^ s_CSAwallace_rca24_and_21_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa37_and0 = s_CSAwallace_rca24_and_22_15 & s_CSAwallace_rca24_and_21_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_and_20_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa37_and1 = s_CSAwallace_rca24_csa5_csa_component_fa37_xor0 & s_CSAwallace_rca24_and_20_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa37_or0 = s_CSAwallace_rca24_csa5_csa_component_fa37_and0 | s_CSAwallace_rca24_csa5_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa38_xor0 = s_CSAwallace_rca24_nand_23_15 ^ s_CSAwallace_rca24_and_22_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa38_and0 = s_CSAwallace_rca24_nand_23_15 & s_CSAwallace_rca24_and_22_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_and_21_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa38_and1 = s_CSAwallace_rca24_csa5_csa_component_fa38_xor0 & s_CSAwallace_rca24_and_21_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa38_or0 = s_CSAwallace_rca24_csa5_csa_component_fa38_and0 | s_CSAwallace_rca24_csa5_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa5_csa_component_fa39_xor0 = ~s_CSAwallace_rca24_nand_23_16;
  assign s_CSAwallace_rca24_csa5_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa5_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_and_22_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa39_and1 = s_CSAwallace_rca24_csa5_csa_component_fa39_xor0 & s_CSAwallace_rca24_and_22_17;
  assign s_CSAwallace_rca24_csa5_csa_component_fa39_or0 = s_CSAwallace_rca24_nand_23_16 | s_CSAwallace_rca24_csa5_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa19_xor0 = s_CSAwallace_rca24_and_1_18 ^ s_CSAwallace_rca24_and_0_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa19_and0 = s_CSAwallace_rca24_and_1_18 & s_CSAwallace_rca24_and_0_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa20_xor0 = s_CSAwallace_rca24_and_2_18 ^ s_CSAwallace_rca24_and_1_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa20_and0 = s_CSAwallace_rca24_and_2_18 & s_CSAwallace_rca24_and_1_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_and_0_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa20_and1 = s_CSAwallace_rca24_csa6_csa_component_fa20_xor0 & s_CSAwallace_rca24_and_0_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa20_or0 = s_CSAwallace_rca24_csa6_csa_component_fa20_and0 | s_CSAwallace_rca24_csa6_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa21_xor0 = s_CSAwallace_rca24_and_3_18 ^ s_CSAwallace_rca24_and_2_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa21_and0 = s_CSAwallace_rca24_and_3_18 & s_CSAwallace_rca24_and_2_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_and_1_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa21_and1 = s_CSAwallace_rca24_csa6_csa_component_fa21_xor0 & s_CSAwallace_rca24_and_1_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa21_or0 = s_CSAwallace_rca24_csa6_csa_component_fa21_and0 | s_CSAwallace_rca24_csa6_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa22_xor0 = s_CSAwallace_rca24_and_4_18 ^ s_CSAwallace_rca24_and_3_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa22_and0 = s_CSAwallace_rca24_and_4_18 & s_CSAwallace_rca24_and_3_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_and_2_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa22_and1 = s_CSAwallace_rca24_csa6_csa_component_fa22_xor0 & s_CSAwallace_rca24_and_2_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa22_or0 = s_CSAwallace_rca24_csa6_csa_component_fa22_and0 | s_CSAwallace_rca24_csa6_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa23_xor0 = s_CSAwallace_rca24_and_5_18 ^ s_CSAwallace_rca24_and_4_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa23_and0 = s_CSAwallace_rca24_and_5_18 & s_CSAwallace_rca24_and_4_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_and_3_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa23_and1 = s_CSAwallace_rca24_csa6_csa_component_fa23_xor0 & s_CSAwallace_rca24_and_3_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa23_or0 = s_CSAwallace_rca24_csa6_csa_component_fa23_and0 | s_CSAwallace_rca24_csa6_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa24_xor0 = s_CSAwallace_rca24_and_6_18 ^ s_CSAwallace_rca24_and_5_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa24_and0 = s_CSAwallace_rca24_and_6_18 & s_CSAwallace_rca24_and_5_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_and_4_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa24_and1 = s_CSAwallace_rca24_csa6_csa_component_fa24_xor0 & s_CSAwallace_rca24_and_4_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa24_or0 = s_CSAwallace_rca24_csa6_csa_component_fa24_and0 | s_CSAwallace_rca24_csa6_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa25_xor0 = s_CSAwallace_rca24_and_7_18 ^ s_CSAwallace_rca24_and_6_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa25_and0 = s_CSAwallace_rca24_and_7_18 & s_CSAwallace_rca24_and_6_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_and_5_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa25_and1 = s_CSAwallace_rca24_csa6_csa_component_fa25_xor0 & s_CSAwallace_rca24_and_5_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa25_or0 = s_CSAwallace_rca24_csa6_csa_component_fa25_and0 | s_CSAwallace_rca24_csa6_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa26_xor0 = s_CSAwallace_rca24_and_8_18 ^ s_CSAwallace_rca24_and_7_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa26_and0 = s_CSAwallace_rca24_and_8_18 & s_CSAwallace_rca24_and_7_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_and_6_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa26_and1 = s_CSAwallace_rca24_csa6_csa_component_fa26_xor0 & s_CSAwallace_rca24_and_6_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa26_or0 = s_CSAwallace_rca24_csa6_csa_component_fa26_and0 | s_CSAwallace_rca24_csa6_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa27_xor0 = s_CSAwallace_rca24_and_9_18 ^ s_CSAwallace_rca24_and_8_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa27_and0 = s_CSAwallace_rca24_and_9_18 & s_CSAwallace_rca24_and_8_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_and_7_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa27_and1 = s_CSAwallace_rca24_csa6_csa_component_fa27_xor0 & s_CSAwallace_rca24_and_7_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa27_or0 = s_CSAwallace_rca24_csa6_csa_component_fa27_and0 | s_CSAwallace_rca24_csa6_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa28_xor0 = s_CSAwallace_rca24_and_10_18 ^ s_CSAwallace_rca24_and_9_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa28_and0 = s_CSAwallace_rca24_and_10_18 & s_CSAwallace_rca24_and_9_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_and_8_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa28_and1 = s_CSAwallace_rca24_csa6_csa_component_fa28_xor0 & s_CSAwallace_rca24_and_8_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa28_or0 = s_CSAwallace_rca24_csa6_csa_component_fa28_and0 | s_CSAwallace_rca24_csa6_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa29_xor0 = s_CSAwallace_rca24_and_11_18 ^ s_CSAwallace_rca24_and_10_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa29_and0 = s_CSAwallace_rca24_and_11_18 & s_CSAwallace_rca24_and_10_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_and_9_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa29_and1 = s_CSAwallace_rca24_csa6_csa_component_fa29_xor0 & s_CSAwallace_rca24_and_9_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa29_or0 = s_CSAwallace_rca24_csa6_csa_component_fa29_and0 | s_CSAwallace_rca24_csa6_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa30_xor0 = s_CSAwallace_rca24_and_12_18 ^ s_CSAwallace_rca24_and_11_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa30_and0 = s_CSAwallace_rca24_and_12_18 & s_CSAwallace_rca24_and_11_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_and_10_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa30_and1 = s_CSAwallace_rca24_csa6_csa_component_fa30_xor0 & s_CSAwallace_rca24_and_10_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa30_or0 = s_CSAwallace_rca24_csa6_csa_component_fa30_and0 | s_CSAwallace_rca24_csa6_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa31_xor0 = s_CSAwallace_rca24_and_13_18 ^ s_CSAwallace_rca24_and_12_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa31_and0 = s_CSAwallace_rca24_and_13_18 & s_CSAwallace_rca24_and_12_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_and_11_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa31_and1 = s_CSAwallace_rca24_csa6_csa_component_fa31_xor0 & s_CSAwallace_rca24_and_11_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa31_or0 = s_CSAwallace_rca24_csa6_csa_component_fa31_and0 | s_CSAwallace_rca24_csa6_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa32_xor0 = s_CSAwallace_rca24_and_14_18 ^ s_CSAwallace_rca24_and_13_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa32_and0 = s_CSAwallace_rca24_and_14_18 & s_CSAwallace_rca24_and_13_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_and_12_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa32_and1 = s_CSAwallace_rca24_csa6_csa_component_fa32_xor0 & s_CSAwallace_rca24_and_12_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa32_or0 = s_CSAwallace_rca24_csa6_csa_component_fa32_and0 | s_CSAwallace_rca24_csa6_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa33_xor0 = s_CSAwallace_rca24_and_15_18 ^ s_CSAwallace_rca24_and_14_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa33_and0 = s_CSAwallace_rca24_and_15_18 & s_CSAwallace_rca24_and_14_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_and_13_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa33_and1 = s_CSAwallace_rca24_csa6_csa_component_fa33_xor0 & s_CSAwallace_rca24_and_13_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa33_or0 = s_CSAwallace_rca24_csa6_csa_component_fa33_and0 | s_CSAwallace_rca24_csa6_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa34_xor0 = s_CSAwallace_rca24_and_16_18 ^ s_CSAwallace_rca24_and_15_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa34_and0 = s_CSAwallace_rca24_and_16_18 & s_CSAwallace_rca24_and_15_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_and_14_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa34_and1 = s_CSAwallace_rca24_csa6_csa_component_fa34_xor0 & s_CSAwallace_rca24_and_14_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa34_or0 = s_CSAwallace_rca24_csa6_csa_component_fa34_and0 | s_CSAwallace_rca24_csa6_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa35_xor0 = s_CSAwallace_rca24_and_17_18 ^ s_CSAwallace_rca24_and_16_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa35_and0 = s_CSAwallace_rca24_and_17_18 & s_CSAwallace_rca24_and_16_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_and_15_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa35_and1 = s_CSAwallace_rca24_csa6_csa_component_fa35_xor0 & s_CSAwallace_rca24_and_15_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa35_or0 = s_CSAwallace_rca24_csa6_csa_component_fa35_and0 | s_CSAwallace_rca24_csa6_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa36_xor0 = s_CSAwallace_rca24_and_18_18 ^ s_CSAwallace_rca24_and_17_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa36_and0 = s_CSAwallace_rca24_and_18_18 & s_CSAwallace_rca24_and_17_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_and_16_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa36_and1 = s_CSAwallace_rca24_csa6_csa_component_fa36_xor0 & s_CSAwallace_rca24_and_16_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa36_or0 = s_CSAwallace_rca24_csa6_csa_component_fa36_and0 | s_CSAwallace_rca24_csa6_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa37_xor0 = s_CSAwallace_rca24_and_19_18 ^ s_CSAwallace_rca24_and_18_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa37_and0 = s_CSAwallace_rca24_and_19_18 & s_CSAwallace_rca24_and_18_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_and_17_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa37_and1 = s_CSAwallace_rca24_csa6_csa_component_fa37_xor0 & s_CSAwallace_rca24_and_17_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa37_or0 = s_CSAwallace_rca24_csa6_csa_component_fa37_and0 | s_CSAwallace_rca24_csa6_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa38_xor0 = s_CSAwallace_rca24_and_20_18 ^ s_CSAwallace_rca24_and_19_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa38_and0 = s_CSAwallace_rca24_and_20_18 & s_CSAwallace_rca24_and_19_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_and_18_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa38_and1 = s_CSAwallace_rca24_csa6_csa_component_fa38_xor0 & s_CSAwallace_rca24_and_18_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa38_or0 = s_CSAwallace_rca24_csa6_csa_component_fa38_and0 | s_CSAwallace_rca24_csa6_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa39_xor0 = s_CSAwallace_rca24_and_21_18 ^ s_CSAwallace_rca24_and_20_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa39_and0 = s_CSAwallace_rca24_and_21_18 & s_CSAwallace_rca24_and_20_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_and_19_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa39_and1 = s_CSAwallace_rca24_csa6_csa_component_fa39_xor0 & s_CSAwallace_rca24_and_19_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa39_or0 = s_CSAwallace_rca24_csa6_csa_component_fa39_and0 | s_CSAwallace_rca24_csa6_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa40_xor0 = s_CSAwallace_rca24_and_22_18 ^ s_CSAwallace_rca24_and_21_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa40_and0 = s_CSAwallace_rca24_and_22_18 & s_CSAwallace_rca24_and_21_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa40_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa40_xor0 ^ s_CSAwallace_rca24_and_20_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa40_and1 = s_CSAwallace_rca24_csa6_csa_component_fa40_xor0 & s_CSAwallace_rca24_and_20_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa40_or0 = s_CSAwallace_rca24_csa6_csa_component_fa40_and0 | s_CSAwallace_rca24_csa6_csa_component_fa40_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa41_xor0 = s_CSAwallace_rca24_nand_23_18 ^ s_CSAwallace_rca24_and_22_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa41_and0 = s_CSAwallace_rca24_nand_23_18 & s_CSAwallace_rca24_and_22_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa41_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa41_xor0 ^ s_CSAwallace_rca24_and_21_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa41_and1 = s_CSAwallace_rca24_csa6_csa_component_fa41_xor0 & s_CSAwallace_rca24_and_21_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa41_or0 = s_CSAwallace_rca24_csa6_csa_component_fa41_and0 | s_CSAwallace_rca24_csa6_csa_component_fa41_and1;
  assign s_CSAwallace_rca24_csa6_csa_component_fa42_xor0 = ~s_CSAwallace_rca24_nand_23_19;
  assign s_CSAwallace_rca24_csa6_csa_component_fa42_xor1 = s_CSAwallace_rca24_csa6_csa_component_fa42_xor0 ^ s_CSAwallace_rca24_and_22_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa42_and1 = s_CSAwallace_rca24_csa6_csa_component_fa42_xor0 & s_CSAwallace_rca24_and_22_20;
  assign s_CSAwallace_rca24_csa6_csa_component_fa42_or0 = s_CSAwallace_rca24_nand_23_19 | s_CSAwallace_rca24_csa6_csa_component_fa42_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa22_xor0 = s_CSAwallace_rca24_and_1_21 ^ s_CSAwallace_rca24_and_0_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa22_and0 = s_CSAwallace_rca24_and_1_21 & s_CSAwallace_rca24_and_0_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa23_xor0 = s_CSAwallace_rca24_and_2_21 ^ s_CSAwallace_rca24_and_1_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa23_and0 = s_CSAwallace_rca24_and_2_21 & s_CSAwallace_rca24_and_1_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_nand_0_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa23_and1 = s_CSAwallace_rca24_csa7_csa_component_fa23_xor0 & s_CSAwallace_rca24_nand_0_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa23_or0 = s_CSAwallace_rca24_csa7_csa_component_fa23_and0 | s_CSAwallace_rca24_csa7_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa24_xor0 = s_CSAwallace_rca24_and_3_21 ^ s_CSAwallace_rca24_and_2_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa24_and0 = s_CSAwallace_rca24_and_3_21 & s_CSAwallace_rca24_and_2_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_nand_1_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa24_and1 = s_CSAwallace_rca24_csa7_csa_component_fa24_xor0 & s_CSAwallace_rca24_nand_1_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa24_or0 = s_CSAwallace_rca24_csa7_csa_component_fa24_and0 | s_CSAwallace_rca24_csa7_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa25_xor0 = s_CSAwallace_rca24_and_4_21 ^ s_CSAwallace_rca24_and_3_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa25_and0 = s_CSAwallace_rca24_and_4_21 & s_CSAwallace_rca24_and_3_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_nand_2_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa25_and1 = s_CSAwallace_rca24_csa7_csa_component_fa25_xor0 & s_CSAwallace_rca24_nand_2_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa25_or0 = s_CSAwallace_rca24_csa7_csa_component_fa25_and0 | s_CSAwallace_rca24_csa7_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa26_xor0 = s_CSAwallace_rca24_and_5_21 ^ s_CSAwallace_rca24_and_4_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa26_and0 = s_CSAwallace_rca24_and_5_21 & s_CSAwallace_rca24_and_4_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_nand_3_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa26_and1 = s_CSAwallace_rca24_csa7_csa_component_fa26_xor0 & s_CSAwallace_rca24_nand_3_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa26_or0 = s_CSAwallace_rca24_csa7_csa_component_fa26_and0 | s_CSAwallace_rca24_csa7_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa27_xor0 = s_CSAwallace_rca24_and_6_21 ^ s_CSAwallace_rca24_and_5_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa27_and0 = s_CSAwallace_rca24_and_6_21 & s_CSAwallace_rca24_and_5_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_nand_4_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa27_and1 = s_CSAwallace_rca24_csa7_csa_component_fa27_xor0 & s_CSAwallace_rca24_nand_4_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa27_or0 = s_CSAwallace_rca24_csa7_csa_component_fa27_and0 | s_CSAwallace_rca24_csa7_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa28_xor0 = s_CSAwallace_rca24_and_7_21 ^ s_CSAwallace_rca24_and_6_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa28_and0 = s_CSAwallace_rca24_and_7_21 & s_CSAwallace_rca24_and_6_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_nand_5_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa28_and1 = s_CSAwallace_rca24_csa7_csa_component_fa28_xor0 & s_CSAwallace_rca24_nand_5_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa28_or0 = s_CSAwallace_rca24_csa7_csa_component_fa28_and0 | s_CSAwallace_rca24_csa7_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa29_xor0 = s_CSAwallace_rca24_and_8_21 ^ s_CSAwallace_rca24_and_7_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa29_and0 = s_CSAwallace_rca24_and_8_21 & s_CSAwallace_rca24_and_7_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_nand_6_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa29_and1 = s_CSAwallace_rca24_csa7_csa_component_fa29_xor0 & s_CSAwallace_rca24_nand_6_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa29_or0 = s_CSAwallace_rca24_csa7_csa_component_fa29_and0 | s_CSAwallace_rca24_csa7_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa30_xor0 = s_CSAwallace_rca24_and_9_21 ^ s_CSAwallace_rca24_and_8_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa30_and0 = s_CSAwallace_rca24_and_9_21 & s_CSAwallace_rca24_and_8_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_nand_7_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa30_and1 = s_CSAwallace_rca24_csa7_csa_component_fa30_xor0 & s_CSAwallace_rca24_nand_7_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa30_or0 = s_CSAwallace_rca24_csa7_csa_component_fa30_and0 | s_CSAwallace_rca24_csa7_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa31_xor0 = s_CSAwallace_rca24_and_10_21 ^ s_CSAwallace_rca24_and_9_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa31_and0 = s_CSAwallace_rca24_and_10_21 & s_CSAwallace_rca24_and_9_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_nand_8_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa31_and1 = s_CSAwallace_rca24_csa7_csa_component_fa31_xor0 & s_CSAwallace_rca24_nand_8_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa31_or0 = s_CSAwallace_rca24_csa7_csa_component_fa31_and0 | s_CSAwallace_rca24_csa7_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa32_xor0 = s_CSAwallace_rca24_and_11_21 ^ s_CSAwallace_rca24_and_10_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa32_and0 = s_CSAwallace_rca24_and_11_21 & s_CSAwallace_rca24_and_10_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_nand_9_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa32_and1 = s_CSAwallace_rca24_csa7_csa_component_fa32_xor0 & s_CSAwallace_rca24_nand_9_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa32_or0 = s_CSAwallace_rca24_csa7_csa_component_fa32_and0 | s_CSAwallace_rca24_csa7_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa33_xor0 = s_CSAwallace_rca24_and_12_21 ^ s_CSAwallace_rca24_and_11_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa33_and0 = s_CSAwallace_rca24_and_12_21 & s_CSAwallace_rca24_and_11_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_nand_10_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa33_and1 = s_CSAwallace_rca24_csa7_csa_component_fa33_xor0 & s_CSAwallace_rca24_nand_10_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa33_or0 = s_CSAwallace_rca24_csa7_csa_component_fa33_and0 | s_CSAwallace_rca24_csa7_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa34_xor0 = s_CSAwallace_rca24_and_13_21 ^ s_CSAwallace_rca24_and_12_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa34_and0 = s_CSAwallace_rca24_and_13_21 & s_CSAwallace_rca24_and_12_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_nand_11_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa34_and1 = s_CSAwallace_rca24_csa7_csa_component_fa34_xor0 & s_CSAwallace_rca24_nand_11_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa34_or0 = s_CSAwallace_rca24_csa7_csa_component_fa34_and0 | s_CSAwallace_rca24_csa7_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa35_xor0 = s_CSAwallace_rca24_and_14_21 ^ s_CSAwallace_rca24_and_13_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa35_and0 = s_CSAwallace_rca24_and_14_21 & s_CSAwallace_rca24_and_13_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_nand_12_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa35_and1 = s_CSAwallace_rca24_csa7_csa_component_fa35_xor0 & s_CSAwallace_rca24_nand_12_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa35_or0 = s_CSAwallace_rca24_csa7_csa_component_fa35_and0 | s_CSAwallace_rca24_csa7_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa36_xor0 = s_CSAwallace_rca24_and_15_21 ^ s_CSAwallace_rca24_and_14_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa36_and0 = s_CSAwallace_rca24_and_15_21 & s_CSAwallace_rca24_and_14_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_nand_13_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa36_and1 = s_CSAwallace_rca24_csa7_csa_component_fa36_xor0 & s_CSAwallace_rca24_nand_13_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa36_or0 = s_CSAwallace_rca24_csa7_csa_component_fa36_and0 | s_CSAwallace_rca24_csa7_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa37_xor0 = s_CSAwallace_rca24_and_16_21 ^ s_CSAwallace_rca24_and_15_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa37_and0 = s_CSAwallace_rca24_and_16_21 & s_CSAwallace_rca24_and_15_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_nand_14_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa37_and1 = s_CSAwallace_rca24_csa7_csa_component_fa37_xor0 & s_CSAwallace_rca24_nand_14_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa37_or0 = s_CSAwallace_rca24_csa7_csa_component_fa37_and0 | s_CSAwallace_rca24_csa7_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa38_xor0 = s_CSAwallace_rca24_and_17_21 ^ s_CSAwallace_rca24_and_16_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa38_and0 = s_CSAwallace_rca24_and_17_21 & s_CSAwallace_rca24_and_16_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_nand_15_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa38_and1 = s_CSAwallace_rca24_csa7_csa_component_fa38_xor0 & s_CSAwallace_rca24_nand_15_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa38_or0 = s_CSAwallace_rca24_csa7_csa_component_fa38_and0 | s_CSAwallace_rca24_csa7_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa39_xor0 = s_CSAwallace_rca24_and_18_21 ^ s_CSAwallace_rca24_and_17_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa39_and0 = s_CSAwallace_rca24_and_18_21 & s_CSAwallace_rca24_and_17_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_nand_16_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa39_and1 = s_CSAwallace_rca24_csa7_csa_component_fa39_xor0 & s_CSAwallace_rca24_nand_16_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa39_or0 = s_CSAwallace_rca24_csa7_csa_component_fa39_and0 | s_CSAwallace_rca24_csa7_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa40_xor0 = s_CSAwallace_rca24_and_19_21 ^ s_CSAwallace_rca24_and_18_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa40_and0 = s_CSAwallace_rca24_and_19_21 & s_CSAwallace_rca24_and_18_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa40_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa40_xor0 ^ s_CSAwallace_rca24_nand_17_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa40_and1 = s_CSAwallace_rca24_csa7_csa_component_fa40_xor0 & s_CSAwallace_rca24_nand_17_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa40_or0 = s_CSAwallace_rca24_csa7_csa_component_fa40_and0 | s_CSAwallace_rca24_csa7_csa_component_fa40_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa41_xor0 = s_CSAwallace_rca24_and_20_21 ^ s_CSAwallace_rca24_and_19_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa41_and0 = s_CSAwallace_rca24_and_20_21 & s_CSAwallace_rca24_and_19_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa41_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa41_xor0 ^ s_CSAwallace_rca24_nand_18_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa41_and1 = s_CSAwallace_rca24_csa7_csa_component_fa41_xor0 & s_CSAwallace_rca24_nand_18_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa41_or0 = s_CSAwallace_rca24_csa7_csa_component_fa41_and0 | s_CSAwallace_rca24_csa7_csa_component_fa41_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa42_xor0 = s_CSAwallace_rca24_and_21_21 ^ s_CSAwallace_rca24_and_20_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa42_and0 = s_CSAwallace_rca24_and_21_21 & s_CSAwallace_rca24_and_20_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa42_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa42_xor0 ^ s_CSAwallace_rca24_nand_19_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa42_and1 = s_CSAwallace_rca24_csa7_csa_component_fa42_xor0 & s_CSAwallace_rca24_nand_19_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa42_or0 = s_CSAwallace_rca24_csa7_csa_component_fa42_and0 | s_CSAwallace_rca24_csa7_csa_component_fa42_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa43_xor0 = s_CSAwallace_rca24_and_22_21 ^ s_CSAwallace_rca24_and_21_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa43_and0 = s_CSAwallace_rca24_and_22_21 & s_CSAwallace_rca24_and_21_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa43_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa43_xor0 ^ s_CSAwallace_rca24_nand_20_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa43_and1 = s_CSAwallace_rca24_csa7_csa_component_fa43_xor0 & s_CSAwallace_rca24_nand_20_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa43_or0 = s_CSAwallace_rca24_csa7_csa_component_fa43_and0 | s_CSAwallace_rca24_csa7_csa_component_fa43_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa44_xor0 = s_CSAwallace_rca24_nand_23_21 ^ s_CSAwallace_rca24_and_22_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa44_and0 = s_CSAwallace_rca24_nand_23_21 & s_CSAwallace_rca24_and_22_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa44_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa44_xor0 ^ s_CSAwallace_rca24_nand_21_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa44_and1 = s_CSAwallace_rca24_csa7_csa_component_fa44_xor0 & s_CSAwallace_rca24_nand_21_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa44_or0 = s_CSAwallace_rca24_csa7_csa_component_fa44_and0 | s_CSAwallace_rca24_csa7_csa_component_fa44_and1;
  assign s_CSAwallace_rca24_csa7_csa_component_fa45_xor0 = ~s_CSAwallace_rca24_nand_23_22;
  assign s_CSAwallace_rca24_csa7_csa_component_fa45_xor1 = s_CSAwallace_rca24_csa7_csa_component_fa45_xor0 ^ s_CSAwallace_rca24_nand_22_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa45_and1 = s_CSAwallace_rca24_csa7_csa_component_fa45_xor0 & s_CSAwallace_rca24_nand_22_23;
  assign s_CSAwallace_rca24_csa7_csa_component_fa45_or0 = s_CSAwallace_rca24_nand_23_22 | s_CSAwallace_rca24_csa7_csa_component_fa45_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa2_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa2_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa1_and0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa2_and0 = s_CSAwallace_rca24_csa0_csa_component_fa2_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa1_and0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa3_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa3_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa2_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa3_and0 = s_CSAwallace_rca24_csa0_csa_component_fa3_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa2_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa3_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa3_xor0 ^ s_CSAwallace_rca24_and_0_3;
  assign s_CSAwallace_rca24_csa8_csa_component_fa3_and1 = s_CSAwallace_rca24_csa8_csa_component_fa3_xor0 & s_CSAwallace_rca24_and_0_3;
  assign s_CSAwallace_rca24_csa8_csa_component_fa3_or0 = s_CSAwallace_rca24_csa8_csa_component_fa3_and0 | s_CSAwallace_rca24_csa8_csa_component_fa3_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa4_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa4_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa3_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa4_and0 = s_CSAwallace_rca24_csa0_csa_component_fa4_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa3_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa4_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa4_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa4_xor0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa4_and1 = s_CSAwallace_rca24_csa8_csa_component_fa4_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa4_xor0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa4_or0 = s_CSAwallace_rca24_csa8_csa_component_fa4_and0 | s_CSAwallace_rca24_csa8_csa_component_fa4_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa5_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa5_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa4_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa5_and0 = s_CSAwallace_rca24_csa0_csa_component_fa5_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa4_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa5_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa5_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa5_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa5_and1 = s_CSAwallace_rca24_csa8_csa_component_fa5_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa5_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa5_or0 = s_CSAwallace_rca24_csa8_csa_component_fa5_and0 | s_CSAwallace_rca24_csa8_csa_component_fa5_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa6_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa6_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa5_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa6_and0 = s_CSAwallace_rca24_csa0_csa_component_fa6_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa5_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa6_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa6_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa6_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa6_and1 = s_CSAwallace_rca24_csa8_csa_component_fa6_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa6_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa6_or0 = s_CSAwallace_rca24_csa8_csa_component_fa6_and0 | s_CSAwallace_rca24_csa8_csa_component_fa6_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa7_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa7_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa6_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa7_and0 = s_CSAwallace_rca24_csa0_csa_component_fa7_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa6_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa7_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa7_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa7_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa7_and1 = s_CSAwallace_rca24_csa8_csa_component_fa7_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa7_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa7_or0 = s_CSAwallace_rca24_csa8_csa_component_fa7_and0 | s_CSAwallace_rca24_csa8_csa_component_fa7_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa8_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa8_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa7_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa8_and0 = s_CSAwallace_rca24_csa0_csa_component_fa8_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa7_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa8_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa8_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa8_and1 = s_CSAwallace_rca24_csa8_csa_component_fa8_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa8_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa8_or0 = s_CSAwallace_rca24_csa8_csa_component_fa8_and0 | s_CSAwallace_rca24_csa8_csa_component_fa8_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa9_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa9_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa9_and0 = s_CSAwallace_rca24_csa0_csa_component_fa9_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa9_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa9_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa9_and1 = s_CSAwallace_rca24_csa8_csa_component_fa9_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa9_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa9_or0 = s_CSAwallace_rca24_csa8_csa_component_fa9_and0 | s_CSAwallace_rca24_csa8_csa_component_fa9_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa10_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa10_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa10_and0 = s_CSAwallace_rca24_csa0_csa_component_fa10_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa10_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa10_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa10_and1 = s_CSAwallace_rca24_csa8_csa_component_fa10_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa10_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa10_or0 = s_CSAwallace_rca24_csa8_csa_component_fa10_and0 | s_CSAwallace_rca24_csa8_csa_component_fa10_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa11_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa11_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa11_and0 = s_CSAwallace_rca24_csa0_csa_component_fa11_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa11_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa11_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa11_and1 = s_CSAwallace_rca24_csa8_csa_component_fa11_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa11_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa11_or0 = s_CSAwallace_rca24_csa8_csa_component_fa11_and0 | s_CSAwallace_rca24_csa8_csa_component_fa11_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa12_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa12_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa12_and0 = s_CSAwallace_rca24_csa0_csa_component_fa12_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa12_and1 = s_CSAwallace_rca24_csa8_csa_component_fa12_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa12_or0 = s_CSAwallace_rca24_csa8_csa_component_fa12_and0 | s_CSAwallace_rca24_csa8_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa13_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa13_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa13_and0 = s_CSAwallace_rca24_csa0_csa_component_fa13_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa13_and1 = s_CSAwallace_rca24_csa8_csa_component_fa13_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa13_or0 = s_CSAwallace_rca24_csa8_csa_component_fa13_and0 | s_CSAwallace_rca24_csa8_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa14_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa14_and0 = s_CSAwallace_rca24_csa0_csa_component_fa14_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa14_and1 = s_CSAwallace_rca24_csa8_csa_component_fa14_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa14_or0 = s_CSAwallace_rca24_csa8_csa_component_fa14_and0 | s_CSAwallace_rca24_csa8_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa15_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa15_and0 = s_CSAwallace_rca24_csa0_csa_component_fa15_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa15_and1 = s_CSAwallace_rca24_csa8_csa_component_fa15_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa15_or0 = s_CSAwallace_rca24_csa8_csa_component_fa15_and0 | s_CSAwallace_rca24_csa8_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa16_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa16_and0 = s_CSAwallace_rca24_csa0_csa_component_fa16_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa16_and1 = s_CSAwallace_rca24_csa8_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa16_or0 = s_CSAwallace_rca24_csa8_csa_component_fa16_and0 | s_CSAwallace_rca24_csa8_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa17_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa17_and0 = s_CSAwallace_rca24_csa0_csa_component_fa17_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa17_and1 = s_CSAwallace_rca24_csa8_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa17_or0 = s_CSAwallace_rca24_csa8_csa_component_fa17_and0 | s_CSAwallace_rca24_csa8_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa18_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa18_and0 = s_CSAwallace_rca24_csa0_csa_component_fa18_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa18_and1 = s_CSAwallace_rca24_csa8_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa18_or0 = s_CSAwallace_rca24_csa8_csa_component_fa18_and0 | s_CSAwallace_rca24_csa8_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa19_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa19_and0 = s_CSAwallace_rca24_csa0_csa_component_fa19_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa19_and1 = s_CSAwallace_rca24_csa8_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa19_or0 = s_CSAwallace_rca24_csa8_csa_component_fa19_and0 | s_CSAwallace_rca24_csa8_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa20_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa20_and0 = s_CSAwallace_rca24_csa0_csa_component_fa20_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa20_and1 = s_CSAwallace_rca24_csa8_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa20_or0 = s_CSAwallace_rca24_csa8_csa_component_fa20_and0 | s_CSAwallace_rca24_csa8_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa21_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa21_and0 = s_CSAwallace_rca24_csa0_csa_component_fa21_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa21_and1 = s_CSAwallace_rca24_csa8_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa21_or0 = s_CSAwallace_rca24_csa8_csa_component_fa21_and0 | s_CSAwallace_rca24_csa8_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa22_and0 = s_CSAwallace_rca24_csa0_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa22_and1 = s_CSAwallace_rca24_csa8_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa22_or0 = s_CSAwallace_rca24_csa8_csa_component_fa22_and0 | s_CSAwallace_rca24_csa8_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa23_and0 = s_CSAwallace_rca24_csa0_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa23_and1 = s_CSAwallace_rca24_csa8_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa23_or0 = s_CSAwallace_rca24_csa8_csa_component_fa23_and0 | s_CSAwallace_rca24_csa8_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa0_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa0_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa24_and0 = s_CSAwallace_rca24_csa0_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa0_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa24_and1 = s_CSAwallace_rca24_csa8_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa24_or0 = s_CSAwallace_rca24_csa8_csa_component_fa24_and0 | s_CSAwallace_rca24_csa8_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa25_xor0 = s_CSAwallace_rca24_nand_23_2 ^ s_CSAwallace_rca24_csa0_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa25_and0 = s_CSAwallace_rca24_nand_23_2 & s_CSAwallace_rca24_csa0_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa8_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa8_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa25_and1 = s_CSAwallace_rca24_csa8_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa8_csa_component_fa25_or0 = s_CSAwallace_rca24_csa8_csa_component_fa25_and0 | s_CSAwallace_rca24_csa8_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa6_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa5_or0 ^ s_CSAwallace_rca24_and_0_6;
  assign s_CSAwallace_rca24_csa9_csa_component_fa6_and0 = s_CSAwallace_rca24_csa1_csa_component_fa5_or0 & s_CSAwallace_rca24_and_0_6;
  assign s_CSAwallace_rca24_csa9_csa_component_fa7_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa6_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa7_xor0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa7_and0 = s_CSAwallace_rca24_csa1_csa_component_fa6_or0 & s_CSAwallace_rca24_csa2_csa_component_fa7_xor0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa8_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa7_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa8_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa8_and0 = s_CSAwallace_rca24_csa1_csa_component_fa7_or0 & s_CSAwallace_rca24_csa2_csa_component_fa8_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa8_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa8_and1 = s_CSAwallace_rca24_csa9_csa_component_fa8_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa8_or0 = s_CSAwallace_rca24_csa9_csa_component_fa8_and0 | s_CSAwallace_rca24_csa9_csa_component_fa8_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa9_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa8_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa9_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa9_and0 = s_CSAwallace_rca24_csa1_csa_component_fa8_or0 & s_CSAwallace_rca24_csa2_csa_component_fa9_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa9_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa9_and1 = s_CSAwallace_rca24_csa9_csa_component_fa9_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa9_or0 = s_CSAwallace_rca24_csa9_csa_component_fa9_and0 | s_CSAwallace_rca24_csa9_csa_component_fa9_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa10_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa9_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa10_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa10_and0 = s_CSAwallace_rca24_csa1_csa_component_fa9_or0 & s_CSAwallace_rca24_csa2_csa_component_fa10_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa10_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa10_and1 = s_CSAwallace_rca24_csa9_csa_component_fa10_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa10_or0 = s_CSAwallace_rca24_csa9_csa_component_fa10_and0 | s_CSAwallace_rca24_csa9_csa_component_fa10_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa11_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa10_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa11_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa11_and0 = s_CSAwallace_rca24_csa1_csa_component_fa10_or0 & s_CSAwallace_rca24_csa2_csa_component_fa11_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa11_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa11_and1 = s_CSAwallace_rca24_csa9_csa_component_fa11_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa11_or0 = s_CSAwallace_rca24_csa9_csa_component_fa11_and0 | s_CSAwallace_rca24_csa9_csa_component_fa11_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa12_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa11_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa12_and0 = s_CSAwallace_rca24_csa1_csa_component_fa11_or0 & s_CSAwallace_rca24_csa2_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa12_and1 = s_CSAwallace_rca24_csa9_csa_component_fa12_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa12_or0 = s_CSAwallace_rca24_csa9_csa_component_fa12_and0 | s_CSAwallace_rca24_csa9_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa13_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa12_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa13_and0 = s_CSAwallace_rca24_csa1_csa_component_fa12_or0 & s_CSAwallace_rca24_csa2_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa13_and1 = s_CSAwallace_rca24_csa9_csa_component_fa13_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa13_or0 = s_CSAwallace_rca24_csa9_csa_component_fa13_and0 | s_CSAwallace_rca24_csa9_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa13_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa14_and0 = s_CSAwallace_rca24_csa1_csa_component_fa13_or0 & s_CSAwallace_rca24_csa2_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa14_and1 = s_CSAwallace_rca24_csa9_csa_component_fa14_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa14_or0 = s_CSAwallace_rca24_csa9_csa_component_fa14_and0 | s_CSAwallace_rca24_csa9_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa14_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa15_and0 = s_CSAwallace_rca24_csa1_csa_component_fa14_or0 & s_CSAwallace_rca24_csa2_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa15_and1 = s_CSAwallace_rca24_csa9_csa_component_fa15_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa15_or0 = s_CSAwallace_rca24_csa9_csa_component_fa15_and0 | s_CSAwallace_rca24_csa9_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa15_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa16_and0 = s_CSAwallace_rca24_csa1_csa_component_fa15_or0 & s_CSAwallace_rca24_csa2_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa16_and1 = s_CSAwallace_rca24_csa9_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa16_or0 = s_CSAwallace_rca24_csa9_csa_component_fa16_and0 | s_CSAwallace_rca24_csa9_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa16_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa17_and0 = s_CSAwallace_rca24_csa1_csa_component_fa16_or0 & s_CSAwallace_rca24_csa2_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa17_and1 = s_CSAwallace_rca24_csa9_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa17_or0 = s_CSAwallace_rca24_csa9_csa_component_fa17_and0 | s_CSAwallace_rca24_csa9_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa17_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa18_and0 = s_CSAwallace_rca24_csa1_csa_component_fa17_or0 & s_CSAwallace_rca24_csa2_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa18_and1 = s_CSAwallace_rca24_csa9_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa18_or0 = s_CSAwallace_rca24_csa9_csa_component_fa18_and0 | s_CSAwallace_rca24_csa9_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa18_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa19_and0 = s_CSAwallace_rca24_csa1_csa_component_fa18_or0 & s_CSAwallace_rca24_csa2_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa19_and1 = s_CSAwallace_rca24_csa9_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa19_or0 = s_CSAwallace_rca24_csa9_csa_component_fa19_and0 | s_CSAwallace_rca24_csa9_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa19_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa20_and0 = s_CSAwallace_rca24_csa1_csa_component_fa19_or0 & s_CSAwallace_rca24_csa2_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa20_and1 = s_CSAwallace_rca24_csa9_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa20_or0 = s_CSAwallace_rca24_csa9_csa_component_fa20_and0 | s_CSAwallace_rca24_csa9_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa20_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa21_and0 = s_CSAwallace_rca24_csa1_csa_component_fa20_or0 & s_CSAwallace_rca24_csa2_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa21_and1 = s_CSAwallace_rca24_csa9_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa21_or0 = s_CSAwallace_rca24_csa9_csa_component_fa21_and0 | s_CSAwallace_rca24_csa9_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa21_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa22_and0 = s_CSAwallace_rca24_csa1_csa_component_fa21_or0 & s_CSAwallace_rca24_csa2_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa22_and1 = s_CSAwallace_rca24_csa9_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa22_or0 = s_CSAwallace_rca24_csa9_csa_component_fa22_and0 | s_CSAwallace_rca24_csa9_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa22_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa23_and0 = s_CSAwallace_rca24_csa1_csa_component_fa22_or0 & s_CSAwallace_rca24_csa2_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa23_and1 = s_CSAwallace_rca24_csa9_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa23_or0 = s_CSAwallace_rca24_csa9_csa_component_fa23_and0 | s_CSAwallace_rca24_csa9_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa23_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa24_and0 = s_CSAwallace_rca24_csa1_csa_component_fa23_or0 & s_CSAwallace_rca24_csa2_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa24_and1 = s_CSAwallace_rca24_csa9_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa24_or0 = s_CSAwallace_rca24_csa9_csa_component_fa24_and0 | s_CSAwallace_rca24_csa9_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa24_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa25_and0 = s_CSAwallace_rca24_csa1_csa_component_fa24_or0 & s_CSAwallace_rca24_csa2_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa25_and1 = s_CSAwallace_rca24_csa9_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa25_or0 = s_CSAwallace_rca24_csa9_csa_component_fa25_and0 | s_CSAwallace_rca24_csa9_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa25_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa26_and0 = s_CSAwallace_rca24_csa1_csa_component_fa25_or0 & s_CSAwallace_rca24_csa2_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa26_and1 = s_CSAwallace_rca24_csa9_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa26_or0 = s_CSAwallace_rca24_csa9_csa_component_fa26_and0 | s_CSAwallace_rca24_csa9_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa26_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa27_and0 = s_CSAwallace_rca24_csa1_csa_component_fa26_or0 & s_CSAwallace_rca24_csa2_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa27_and1 = s_CSAwallace_rca24_csa9_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa27_or0 = s_CSAwallace_rca24_csa9_csa_component_fa27_and0 | s_CSAwallace_rca24_csa9_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa27_or0 ^ s_CSAwallace_rca24_csa2_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa28_and0 = s_CSAwallace_rca24_csa1_csa_component_fa27_or0 & s_CSAwallace_rca24_csa2_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa28_and1 = s_CSAwallace_rca24_csa9_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa28_or0 = s_CSAwallace_rca24_csa9_csa_component_fa28_and0 | s_CSAwallace_rca24_csa9_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa29_xor0 = ~s_CSAwallace_rca24_csa2_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa29_and1 = s_CSAwallace_rca24_csa9_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa29_or0 = s_CSAwallace_rca24_csa2_csa_component_fa29_xor1 | s_CSAwallace_rca24_csa9_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa30_xor0 = ~s_CSAwallace_rca24_csa2_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa30_and1 = s_CSAwallace_rca24_csa9_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa30_or0 = s_CSAwallace_rca24_csa2_csa_component_fa30_xor1 | s_CSAwallace_rca24_csa9_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa9_csa_component_fa31_xor0 = ~s_CSAwallace_rca24_nand_23_8;
  assign s_CSAwallace_rca24_csa9_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa9_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa2_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa31_and1 = s_CSAwallace_rca24_csa9_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa2_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa9_csa_component_fa31_or0 = s_CSAwallace_rca24_nand_23_8 | s_CSAwallace_rca24_csa9_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa11_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa11_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa10_and0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa11_and0 = s_CSAwallace_rca24_csa3_csa_component_fa11_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa10_and0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa12_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa12_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa12_and0 = s_CSAwallace_rca24_csa3_csa_component_fa12_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_and_0_12;
  assign s_CSAwallace_rca24_csa10_csa_component_fa12_and1 = s_CSAwallace_rca24_csa10_csa_component_fa12_xor0 & s_CSAwallace_rca24_and_0_12;
  assign s_CSAwallace_rca24_csa10_csa_component_fa12_or0 = s_CSAwallace_rca24_csa10_csa_component_fa12_and0 | s_CSAwallace_rca24_csa10_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa13_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa13_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa13_and0 = s_CSAwallace_rca24_csa3_csa_component_fa13_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa13_xor0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa13_and1 = s_CSAwallace_rca24_csa10_csa_component_fa13_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa13_xor0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa13_or0 = s_CSAwallace_rca24_csa10_csa_component_fa13_and0 | s_CSAwallace_rca24_csa10_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa14_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa14_and0 = s_CSAwallace_rca24_csa3_csa_component_fa14_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa14_and1 = s_CSAwallace_rca24_csa10_csa_component_fa14_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa14_or0 = s_CSAwallace_rca24_csa10_csa_component_fa14_and0 | s_CSAwallace_rca24_csa10_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa15_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa15_and0 = s_CSAwallace_rca24_csa3_csa_component_fa15_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa15_and1 = s_CSAwallace_rca24_csa10_csa_component_fa15_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa15_or0 = s_CSAwallace_rca24_csa10_csa_component_fa15_and0 | s_CSAwallace_rca24_csa10_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa16_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa16_and0 = s_CSAwallace_rca24_csa3_csa_component_fa16_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa16_and1 = s_CSAwallace_rca24_csa10_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa16_or0 = s_CSAwallace_rca24_csa10_csa_component_fa16_and0 | s_CSAwallace_rca24_csa10_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa17_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa17_and0 = s_CSAwallace_rca24_csa3_csa_component_fa17_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa17_and1 = s_CSAwallace_rca24_csa10_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa17_or0 = s_CSAwallace_rca24_csa10_csa_component_fa17_and0 | s_CSAwallace_rca24_csa10_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa18_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa18_and0 = s_CSAwallace_rca24_csa3_csa_component_fa18_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa18_and1 = s_CSAwallace_rca24_csa10_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa18_or0 = s_CSAwallace_rca24_csa10_csa_component_fa18_and0 | s_CSAwallace_rca24_csa10_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa19_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa19_and0 = s_CSAwallace_rca24_csa3_csa_component_fa19_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa19_and1 = s_CSAwallace_rca24_csa10_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa19_or0 = s_CSAwallace_rca24_csa10_csa_component_fa19_and0 | s_CSAwallace_rca24_csa10_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa20_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa20_and0 = s_CSAwallace_rca24_csa3_csa_component_fa20_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa20_and1 = s_CSAwallace_rca24_csa10_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa20_or0 = s_CSAwallace_rca24_csa10_csa_component_fa20_and0 | s_CSAwallace_rca24_csa10_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa21_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa21_and0 = s_CSAwallace_rca24_csa3_csa_component_fa21_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa21_and1 = s_CSAwallace_rca24_csa10_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa21_or0 = s_CSAwallace_rca24_csa10_csa_component_fa21_and0 | s_CSAwallace_rca24_csa10_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa22_and0 = s_CSAwallace_rca24_csa3_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa22_and1 = s_CSAwallace_rca24_csa10_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa22_or0 = s_CSAwallace_rca24_csa10_csa_component_fa22_and0 | s_CSAwallace_rca24_csa10_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa23_and0 = s_CSAwallace_rca24_csa3_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa23_and1 = s_CSAwallace_rca24_csa10_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa23_or0 = s_CSAwallace_rca24_csa10_csa_component_fa23_and0 | s_CSAwallace_rca24_csa10_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa24_and0 = s_CSAwallace_rca24_csa3_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa24_and1 = s_CSAwallace_rca24_csa10_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa24_or0 = s_CSAwallace_rca24_csa10_csa_component_fa24_and0 | s_CSAwallace_rca24_csa10_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa25_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa25_and0 = s_CSAwallace_rca24_csa3_csa_component_fa25_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa25_and1 = s_CSAwallace_rca24_csa10_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa25_or0 = s_CSAwallace_rca24_csa10_csa_component_fa25_and0 | s_CSAwallace_rca24_csa10_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa26_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa26_and0 = s_CSAwallace_rca24_csa3_csa_component_fa26_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa26_and1 = s_CSAwallace_rca24_csa10_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa26_or0 = s_CSAwallace_rca24_csa10_csa_component_fa26_and0 | s_CSAwallace_rca24_csa10_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa27_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa27_and0 = s_CSAwallace_rca24_csa3_csa_component_fa27_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa27_and1 = s_CSAwallace_rca24_csa10_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa27_or0 = s_CSAwallace_rca24_csa10_csa_component_fa27_and0 | s_CSAwallace_rca24_csa10_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa28_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa28_and0 = s_CSAwallace_rca24_csa3_csa_component_fa28_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa28_and1 = s_CSAwallace_rca24_csa10_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa28_or0 = s_CSAwallace_rca24_csa10_csa_component_fa28_and0 | s_CSAwallace_rca24_csa10_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa29_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa29_and0 = s_CSAwallace_rca24_csa3_csa_component_fa29_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa29_and1 = s_CSAwallace_rca24_csa10_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa29_or0 = s_CSAwallace_rca24_csa10_csa_component_fa29_and0 | s_CSAwallace_rca24_csa10_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa30_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa30_and0 = s_CSAwallace_rca24_csa3_csa_component_fa30_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa30_and1 = s_CSAwallace_rca24_csa10_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa30_or0 = s_CSAwallace_rca24_csa10_csa_component_fa30_and0 | s_CSAwallace_rca24_csa10_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa31_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa31_and0 = s_CSAwallace_rca24_csa3_csa_component_fa31_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa31_and1 = s_CSAwallace_rca24_csa10_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa31_or0 = s_CSAwallace_rca24_csa10_csa_component_fa31_and0 | s_CSAwallace_rca24_csa10_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa32_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa32_and0 = s_CSAwallace_rca24_csa3_csa_component_fa32_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa32_and1 = s_CSAwallace_rca24_csa10_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa32_or0 = s_CSAwallace_rca24_csa10_csa_component_fa32_and0 | s_CSAwallace_rca24_csa10_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa33_xor0 = s_CSAwallace_rca24_csa3_csa_component_fa33_xor1 ^ s_CSAwallace_rca24_csa3_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa33_and0 = s_CSAwallace_rca24_csa3_csa_component_fa33_xor1 & s_CSAwallace_rca24_csa3_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa33_and1 = s_CSAwallace_rca24_csa10_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa33_or0 = s_CSAwallace_rca24_csa10_csa_component_fa33_and0 | s_CSAwallace_rca24_csa10_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa34_xor0 = s_CSAwallace_rca24_nand_23_11 ^ s_CSAwallace_rca24_csa3_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa34_and0 = s_CSAwallace_rca24_nand_23_11 & s_CSAwallace_rca24_csa3_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa10_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa10_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa4_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa34_and1 = s_CSAwallace_rca24_csa10_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa4_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa10_csa_component_fa34_or0 = s_CSAwallace_rca24_csa10_csa_component_fa34_and0 | s_CSAwallace_rca24_csa10_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa14_or0 ^ s_CSAwallace_rca24_and_0_15;
  assign s_CSAwallace_rca24_csa11_csa_component_fa15_and0 = s_CSAwallace_rca24_csa4_csa_component_fa14_or0 & s_CSAwallace_rca24_and_0_15;
  assign s_CSAwallace_rca24_csa11_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa15_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa16_xor0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa16_and0 = s_CSAwallace_rca24_csa4_csa_component_fa15_or0 & s_CSAwallace_rca24_csa5_csa_component_fa16_xor0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa16_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa17_and0 = s_CSAwallace_rca24_csa4_csa_component_fa16_or0 & s_CSAwallace_rca24_csa5_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa17_and1 = s_CSAwallace_rca24_csa11_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa17_or0 = s_CSAwallace_rca24_csa11_csa_component_fa17_and0 | s_CSAwallace_rca24_csa11_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa17_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa18_and0 = s_CSAwallace_rca24_csa4_csa_component_fa17_or0 & s_CSAwallace_rca24_csa5_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa18_and1 = s_CSAwallace_rca24_csa11_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa18_or0 = s_CSAwallace_rca24_csa11_csa_component_fa18_and0 | s_CSAwallace_rca24_csa11_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa18_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa19_and0 = s_CSAwallace_rca24_csa4_csa_component_fa18_or0 & s_CSAwallace_rca24_csa5_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa19_and1 = s_CSAwallace_rca24_csa11_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa19_or0 = s_CSAwallace_rca24_csa11_csa_component_fa19_and0 | s_CSAwallace_rca24_csa11_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa19_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa20_and0 = s_CSAwallace_rca24_csa4_csa_component_fa19_or0 & s_CSAwallace_rca24_csa5_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa20_and1 = s_CSAwallace_rca24_csa11_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa20_or0 = s_CSAwallace_rca24_csa11_csa_component_fa20_and0 | s_CSAwallace_rca24_csa11_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa20_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa21_and0 = s_CSAwallace_rca24_csa4_csa_component_fa20_or0 & s_CSAwallace_rca24_csa5_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa21_and1 = s_CSAwallace_rca24_csa11_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa21_or0 = s_CSAwallace_rca24_csa11_csa_component_fa21_and0 | s_CSAwallace_rca24_csa11_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa21_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa22_and0 = s_CSAwallace_rca24_csa4_csa_component_fa21_or0 & s_CSAwallace_rca24_csa5_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa22_and1 = s_CSAwallace_rca24_csa11_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa22_or0 = s_CSAwallace_rca24_csa11_csa_component_fa22_and0 | s_CSAwallace_rca24_csa11_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa22_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa23_and0 = s_CSAwallace_rca24_csa4_csa_component_fa22_or0 & s_CSAwallace_rca24_csa5_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa23_and1 = s_CSAwallace_rca24_csa11_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa23_or0 = s_CSAwallace_rca24_csa11_csa_component_fa23_and0 | s_CSAwallace_rca24_csa11_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa23_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa24_and0 = s_CSAwallace_rca24_csa4_csa_component_fa23_or0 & s_CSAwallace_rca24_csa5_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa24_and1 = s_CSAwallace_rca24_csa11_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa24_or0 = s_CSAwallace_rca24_csa11_csa_component_fa24_and0 | s_CSAwallace_rca24_csa11_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa24_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa25_and0 = s_CSAwallace_rca24_csa4_csa_component_fa24_or0 & s_CSAwallace_rca24_csa5_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa25_and1 = s_CSAwallace_rca24_csa11_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa25_or0 = s_CSAwallace_rca24_csa11_csa_component_fa25_and0 | s_CSAwallace_rca24_csa11_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa25_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa26_and0 = s_CSAwallace_rca24_csa4_csa_component_fa25_or0 & s_CSAwallace_rca24_csa5_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa26_and1 = s_CSAwallace_rca24_csa11_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa26_or0 = s_CSAwallace_rca24_csa11_csa_component_fa26_and0 | s_CSAwallace_rca24_csa11_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa26_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa27_and0 = s_CSAwallace_rca24_csa4_csa_component_fa26_or0 & s_CSAwallace_rca24_csa5_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa27_and1 = s_CSAwallace_rca24_csa11_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa27_or0 = s_CSAwallace_rca24_csa11_csa_component_fa27_and0 | s_CSAwallace_rca24_csa11_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa27_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa28_and0 = s_CSAwallace_rca24_csa4_csa_component_fa27_or0 & s_CSAwallace_rca24_csa5_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa28_and1 = s_CSAwallace_rca24_csa11_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa28_or0 = s_CSAwallace_rca24_csa11_csa_component_fa28_and0 | s_CSAwallace_rca24_csa11_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa28_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa29_and0 = s_CSAwallace_rca24_csa4_csa_component_fa28_or0 & s_CSAwallace_rca24_csa5_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa29_and1 = s_CSAwallace_rca24_csa11_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa29_or0 = s_CSAwallace_rca24_csa11_csa_component_fa29_and0 | s_CSAwallace_rca24_csa11_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa29_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa30_and0 = s_CSAwallace_rca24_csa4_csa_component_fa29_or0 & s_CSAwallace_rca24_csa5_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa30_and1 = s_CSAwallace_rca24_csa11_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa30_or0 = s_CSAwallace_rca24_csa11_csa_component_fa30_and0 | s_CSAwallace_rca24_csa11_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa30_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa31_and0 = s_CSAwallace_rca24_csa4_csa_component_fa30_or0 & s_CSAwallace_rca24_csa5_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa31_and1 = s_CSAwallace_rca24_csa11_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa31_or0 = s_CSAwallace_rca24_csa11_csa_component_fa31_and0 | s_CSAwallace_rca24_csa11_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa31_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa32_and0 = s_CSAwallace_rca24_csa4_csa_component_fa31_or0 & s_CSAwallace_rca24_csa5_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa32_and1 = s_CSAwallace_rca24_csa11_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa32_or0 = s_CSAwallace_rca24_csa11_csa_component_fa32_and0 | s_CSAwallace_rca24_csa11_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa33_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa32_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa33_and0 = s_CSAwallace_rca24_csa4_csa_component_fa32_or0 & s_CSAwallace_rca24_csa5_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa33_and1 = s_CSAwallace_rca24_csa11_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa33_or0 = s_CSAwallace_rca24_csa11_csa_component_fa33_and0 | s_CSAwallace_rca24_csa11_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa34_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa33_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa34_and0 = s_CSAwallace_rca24_csa4_csa_component_fa33_or0 & s_CSAwallace_rca24_csa5_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa34_and1 = s_CSAwallace_rca24_csa11_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa34_or0 = s_CSAwallace_rca24_csa11_csa_component_fa34_and0 | s_CSAwallace_rca24_csa11_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa35_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa34_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa35_and0 = s_CSAwallace_rca24_csa4_csa_component_fa34_or0 & s_CSAwallace_rca24_csa5_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa35_and1 = s_CSAwallace_rca24_csa11_csa_component_fa35_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa35_or0 = s_CSAwallace_rca24_csa11_csa_component_fa35_and0 | s_CSAwallace_rca24_csa11_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa36_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa35_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa36_and0 = s_CSAwallace_rca24_csa4_csa_component_fa35_or0 & s_CSAwallace_rca24_csa5_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa36_and1 = s_CSAwallace_rca24_csa11_csa_component_fa36_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa36_or0 = s_CSAwallace_rca24_csa11_csa_component_fa36_and0 | s_CSAwallace_rca24_csa11_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa37_xor0 = s_CSAwallace_rca24_csa4_csa_component_fa36_or0 ^ s_CSAwallace_rca24_csa5_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa37_and0 = s_CSAwallace_rca24_csa4_csa_component_fa36_or0 & s_CSAwallace_rca24_csa5_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa37_and1 = s_CSAwallace_rca24_csa11_csa_component_fa37_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa37_or0 = s_CSAwallace_rca24_csa11_csa_component_fa37_and0 | s_CSAwallace_rca24_csa11_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa38_xor0 = ~s_CSAwallace_rca24_csa5_csa_component_fa38_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa38_and1 = s_CSAwallace_rca24_csa11_csa_component_fa38_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa38_or0 = s_CSAwallace_rca24_csa5_csa_component_fa38_xor1 | s_CSAwallace_rca24_csa11_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa39_xor0 = ~s_CSAwallace_rca24_csa5_csa_component_fa39_xor1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa39_and1 = s_CSAwallace_rca24_csa11_csa_component_fa39_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa39_or0 = s_CSAwallace_rca24_csa5_csa_component_fa39_xor1 | s_CSAwallace_rca24_csa11_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa11_csa_component_fa40_xor0 = ~s_CSAwallace_rca24_nand_23_17;
  assign s_CSAwallace_rca24_csa11_csa_component_fa40_xor1 = s_CSAwallace_rca24_csa11_csa_component_fa40_xor0 ^ s_CSAwallace_rca24_csa5_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa40_and1 = s_CSAwallace_rca24_csa11_csa_component_fa40_xor0 & s_CSAwallace_rca24_csa5_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa11_csa_component_fa40_or0 = s_CSAwallace_rca24_nand_23_17 | s_CSAwallace_rca24_csa11_csa_component_fa40_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa20_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa19_and0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa20_and0 = s_CSAwallace_rca24_csa6_csa_component_fa20_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa19_and0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa21_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa21_and0 = s_CSAwallace_rca24_csa6_csa_component_fa21_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_and_0_21;
  assign s_CSAwallace_rca24_csa12_csa_component_fa21_and1 = s_CSAwallace_rca24_csa12_csa_component_fa21_xor0 & s_CSAwallace_rca24_and_0_21;
  assign s_CSAwallace_rca24_csa12_csa_component_fa21_or0 = s_CSAwallace_rca24_csa12_csa_component_fa21_and0 | s_CSAwallace_rca24_csa12_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa22_and0 = s_CSAwallace_rca24_csa6_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa22_xor0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa22_and1 = s_CSAwallace_rca24_csa12_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa22_xor0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa22_or0 = s_CSAwallace_rca24_csa12_csa_component_fa22_and0 | s_CSAwallace_rca24_csa12_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa23_and0 = s_CSAwallace_rca24_csa6_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa23_and1 = s_CSAwallace_rca24_csa12_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa23_or0 = s_CSAwallace_rca24_csa12_csa_component_fa23_and0 | s_CSAwallace_rca24_csa12_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa24_and0 = s_CSAwallace_rca24_csa6_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa24_and1 = s_CSAwallace_rca24_csa12_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa24_or0 = s_CSAwallace_rca24_csa12_csa_component_fa24_and0 | s_CSAwallace_rca24_csa12_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa25_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa25_and0 = s_CSAwallace_rca24_csa6_csa_component_fa25_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa25_and1 = s_CSAwallace_rca24_csa12_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa25_or0 = s_CSAwallace_rca24_csa12_csa_component_fa25_and0 | s_CSAwallace_rca24_csa12_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa26_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa26_and0 = s_CSAwallace_rca24_csa6_csa_component_fa26_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa26_and1 = s_CSAwallace_rca24_csa12_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa26_or0 = s_CSAwallace_rca24_csa12_csa_component_fa26_and0 | s_CSAwallace_rca24_csa12_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa27_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa27_and0 = s_CSAwallace_rca24_csa6_csa_component_fa27_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa27_and1 = s_CSAwallace_rca24_csa12_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa27_or0 = s_CSAwallace_rca24_csa12_csa_component_fa27_and0 | s_CSAwallace_rca24_csa12_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa28_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa28_and0 = s_CSAwallace_rca24_csa6_csa_component_fa28_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa28_and1 = s_CSAwallace_rca24_csa12_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa28_or0 = s_CSAwallace_rca24_csa12_csa_component_fa28_and0 | s_CSAwallace_rca24_csa12_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa29_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa29_and0 = s_CSAwallace_rca24_csa6_csa_component_fa29_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa29_and1 = s_CSAwallace_rca24_csa12_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa29_or0 = s_CSAwallace_rca24_csa12_csa_component_fa29_and0 | s_CSAwallace_rca24_csa12_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa30_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa30_and0 = s_CSAwallace_rca24_csa6_csa_component_fa30_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa30_and1 = s_CSAwallace_rca24_csa12_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa30_or0 = s_CSAwallace_rca24_csa12_csa_component_fa30_and0 | s_CSAwallace_rca24_csa12_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa31_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa31_and0 = s_CSAwallace_rca24_csa6_csa_component_fa31_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa31_and1 = s_CSAwallace_rca24_csa12_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa31_or0 = s_CSAwallace_rca24_csa12_csa_component_fa31_and0 | s_CSAwallace_rca24_csa12_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa32_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa32_and0 = s_CSAwallace_rca24_csa6_csa_component_fa32_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa32_and1 = s_CSAwallace_rca24_csa12_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa32_or0 = s_CSAwallace_rca24_csa12_csa_component_fa32_and0 | s_CSAwallace_rca24_csa12_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa33_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa33_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa33_and0 = s_CSAwallace_rca24_csa6_csa_component_fa33_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa33_and1 = s_CSAwallace_rca24_csa12_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa33_or0 = s_CSAwallace_rca24_csa12_csa_component_fa33_and0 | s_CSAwallace_rca24_csa12_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa34_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa34_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa34_and0 = s_CSAwallace_rca24_csa6_csa_component_fa34_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa34_and1 = s_CSAwallace_rca24_csa12_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa34_or0 = s_CSAwallace_rca24_csa12_csa_component_fa34_and0 | s_CSAwallace_rca24_csa12_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa35_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa35_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa35_and0 = s_CSAwallace_rca24_csa6_csa_component_fa35_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa35_and1 = s_CSAwallace_rca24_csa12_csa_component_fa35_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa35_or0 = s_CSAwallace_rca24_csa12_csa_component_fa35_and0 | s_CSAwallace_rca24_csa12_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa36_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa36_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa36_and0 = s_CSAwallace_rca24_csa6_csa_component_fa36_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa36_and1 = s_CSAwallace_rca24_csa12_csa_component_fa36_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa36_or0 = s_CSAwallace_rca24_csa12_csa_component_fa36_and0 | s_CSAwallace_rca24_csa12_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa37_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa37_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa37_and0 = s_CSAwallace_rca24_csa6_csa_component_fa37_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa37_and1 = s_CSAwallace_rca24_csa12_csa_component_fa37_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa37_or0 = s_CSAwallace_rca24_csa12_csa_component_fa37_and0 | s_CSAwallace_rca24_csa12_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa38_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa38_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa38_and0 = s_CSAwallace_rca24_csa6_csa_component_fa38_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa38_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa38_and1 = s_CSAwallace_rca24_csa12_csa_component_fa38_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa38_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa38_or0 = s_CSAwallace_rca24_csa12_csa_component_fa38_and0 | s_CSAwallace_rca24_csa12_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa39_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa39_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa39_and0 = s_CSAwallace_rca24_csa6_csa_component_fa39_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa39_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa39_and1 = s_CSAwallace_rca24_csa12_csa_component_fa39_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa39_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa39_or0 = s_CSAwallace_rca24_csa12_csa_component_fa39_and0 | s_CSAwallace_rca24_csa12_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa40_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa40_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa40_and0 = s_CSAwallace_rca24_csa6_csa_component_fa40_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa40_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa40_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa40_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa40_and1 = s_CSAwallace_rca24_csa12_csa_component_fa40_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa40_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa40_or0 = s_CSAwallace_rca24_csa12_csa_component_fa40_and0 | s_CSAwallace_rca24_csa12_csa_component_fa40_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa41_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa41_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa41_and0 = s_CSAwallace_rca24_csa6_csa_component_fa41_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa41_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa41_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa41_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa41_and1 = s_CSAwallace_rca24_csa12_csa_component_fa41_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa41_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa41_or0 = s_CSAwallace_rca24_csa12_csa_component_fa41_and0 | s_CSAwallace_rca24_csa12_csa_component_fa41_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa42_xor0 = s_CSAwallace_rca24_csa6_csa_component_fa42_xor1 ^ s_CSAwallace_rca24_csa6_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa42_and0 = s_CSAwallace_rca24_csa6_csa_component_fa42_xor1 & s_CSAwallace_rca24_csa6_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa42_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa42_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa42_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa42_and1 = s_CSAwallace_rca24_csa12_csa_component_fa42_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa42_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa42_or0 = s_CSAwallace_rca24_csa12_csa_component_fa42_and0 | s_CSAwallace_rca24_csa12_csa_component_fa42_and1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa43_xor0 = s_CSAwallace_rca24_nand_23_20 ^ s_CSAwallace_rca24_csa6_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa43_and0 = s_CSAwallace_rca24_nand_23_20 & s_CSAwallace_rca24_csa6_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa12_csa_component_fa43_xor1 = s_CSAwallace_rca24_csa12_csa_component_fa43_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa43_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa43_and1 = s_CSAwallace_rca24_csa12_csa_component_fa43_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa43_xor1;
  assign s_CSAwallace_rca24_csa12_csa_component_fa43_or0 = s_CSAwallace_rca24_csa12_csa_component_fa43_and0 | s_CSAwallace_rca24_csa12_csa_component_fa43_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa3_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa3_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa2_and0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa3_and0 = s_CSAwallace_rca24_csa8_csa_component_fa3_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa2_and0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa4_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa4_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa3_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa4_and0 = s_CSAwallace_rca24_csa8_csa_component_fa4_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa3_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa5_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa5_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa4_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa5_and0 = s_CSAwallace_rca24_csa8_csa_component_fa5_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa4_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa5_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa5_xor0 ^ s_CSAwallace_rca24_csa1_csa_component_fa4_and0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa5_and1 = s_CSAwallace_rca24_csa13_csa_component_fa5_xor0 & s_CSAwallace_rca24_csa1_csa_component_fa4_and0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa5_or0 = s_CSAwallace_rca24_csa13_csa_component_fa5_and0 | s_CSAwallace_rca24_csa13_csa_component_fa5_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa6_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa6_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa5_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa6_and0 = s_CSAwallace_rca24_csa8_csa_component_fa6_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa5_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa6_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa6_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa6_xor0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa6_and1 = s_CSAwallace_rca24_csa13_csa_component_fa6_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa6_xor0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa6_or0 = s_CSAwallace_rca24_csa13_csa_component_fa6_and0 | s_CSAwallace_rca24_csa13_csa_component_fa6_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa7_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa7_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa6_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa7_and0 = s_CSAwallace_rca24_csa8_csa_component_fa7_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa6_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa7_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa7_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa7_xor0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa7_and1 = s_CSAwallace_rca24_csa13_csa_component_fa7_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa7_xor0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa7_or0 = s_CSAwallace_rca24_csa13_csa_component_fa7_and0 | s_CSAwallace_rca24_csa13_csa_component_fa7_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa8_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa8_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa7_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa8_and0 = s_CSAwallace_rca24_csa8_csa_component_fa8_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa7_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa8_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa8_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa8_and1 = s_CSAwallace_rca24_csa13_csa_component_fa8_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa8_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa8_or0 = s_CSAwallace_rca24_csa13_csa_component_fa8_and0 | s_CSAwallace_rca24_csa13_csa_component_fa8_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa9_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa9_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa9_and0 = s_CSAwallace_rca24_csa8_csa_component_fa9_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa9_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa9_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa9_and1 = s_CSAwallace_rca24_csa13_csa_component_fa9_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa9_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa9_or0 = s_CSAwallace_rca24_csa13_csa_component_fa9_and0 | s_CSAwallace_rca24_csa13_csa_component_fa9_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa10_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa10_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa10_and0 = s_CSAwallace_rca24_csa8_csa_component_fa10_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa10_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa10_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa10_and1 = s_CSAwallace_rca24_csa13_csa_component_fa10_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa10_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa10_or0 = s_CSAwallace_rca24_csa13_csa_component_fa10_and0 | s_CSAwallace_rca24_csa13_csa_component_fa10_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa11_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa11_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa11_and0 = s_CSAwallace_rca24_csa8_csa_component_fa11_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa11_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa11_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa11_and1 = s_CSAwallace_rca24_csa13_csa_component_fa11_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa11_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa11_or0 = s_CSAwallace_rca24_csa13_csa_component_fa11_and0 | s_CSAwallace_rca24_csa13_csa_component_fa11_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa12_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa12_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa12_and0 = s_CSAwallace_rca24_csa8_csa_component_fa12_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa12_and1 = s_CSAwallace_rca24_csa13_csa_component_fa12_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa12_or0 = s_CSAwallace_rca24_csa13_csa_component_fa12_and0 | s_CSAwallace_rca24_csa13_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa13_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa13_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa13_and0 = s_CSAwallace_rca24_csa8_csa_component_fa13_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa13_and1 = s_CSAwallace_rca24_csa13_csa_component_fa13_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa13_or0 = s_CSAwallace_rca24_csa13_csa_component_fa13_and0 | s_CSAwallace_rca24_csa13_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa14_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa14_and0 = s_CSAwallace_rca24_csa8_csa_component_fa14_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa14_and1 = s_CSAwallace_rca24_csa13_csa_component_fa14_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa14_or0 = s_CSAwallace_rca24_csa13_csa_component_fa14_and0 | s_CSAwallace_rca24_csa13_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa15_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa15_and0 = s_CSAwallace_rca24_csa8_csa_component_fa15_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa15_and1 = s_CSAwallace_rca24_csa13_csa_component_fa15_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa15_or0 = s_CSAwallace_rca24_csa13_csa_component_fa15_and0 | s_CSAwallace_rca24_csa13_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa16_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa16_and0 = s_CSAwallace_rca24_csa8_csa_component_fa16_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa16_and1 = s_CSAwallace_rca24_csa13_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa16_or0 = s_CSAwallace_rca24_csa13_csa_component_fa16_and0 | s_CSAwallace_rca24_csa13_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa17_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa17_and0 = s_CSAwallace_rca24_csa8_csa_component_fa17_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa17_and1 = s_CSAwallace_rca24_csa13_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa17_or0 = s_CSAwallace_rca24_csa13_csa_component_fa17_and0 | s_CSAwallace_rca24_csa13_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa18_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa18_and0 = s_CSAwallace_rca24_csa8_csa_component_fa18_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa18_and1 = s_CSAwallace_rca24_csa13_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa18_or0 = s_CSAwallace_rca24_csa13_csa_component_fa18_and0 | s_CSAwallace_rca24_csa13_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa19_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa19_and0 = s_CSAwallace_rca24_csa8_csa_component_fa19_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa19_and1 = s_CSAwallace_rca24_csa13_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa19_or0 = s_CSAwallace_rca24_csa13_csa_component_fa19_and0 | s_CSAwallace_rca24_csa13_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa20_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa20_and0 = s_CSAwallace_rca24_csa8_csa_component_fa20_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa20_and1 = s_CSAwallace_rca24_csa13_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa20_or0 = s_CSAwallace_rca24_csa13_csa_component_fa20_and0 | s_CSAwallace_rca24_csa13_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa21_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa21_and0 = s_CSAwallace_rca24_csa8_csa_component_fa21_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa21_and1 = s_CSAwallace_rca24_csa13_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa21_or0 = s_CSAwallace_rca24_csa13_csa_component_fa21_and0 | s_CSAwallace_rca24_csa13_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa22_and0 = s_CSAwallace_rca24_csa8_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa22_and1 = s_CSAwallace_rca24_csa13_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa22_or0 = s_CSAwallace_rca24_csa13_csa_component_fa22_and0 | s_CSAwallace_rca24_csa13_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa23_and0 = s_CSAwallace_rca24_csa8_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa23_and1 = s_CSAwallace_rca24_csa13_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa23_or0 = s_CSAwallace_rca24_csa13_csa_component_fa23_and0 | s_CSAwallace_rca24_csa13_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa24_and0 = s_CSAwallace_rca24_csa8_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa24_and1 = s_CSAwallace_rca24_csa13_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa24_or0 = s_CSAwallace_rca24_csa13_csa_component_fa24_and0 | s_CSAwallace_rca24_csa13_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa8_csa_component_fa25_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa25_and0 = s_CSAwallace_rca24_csa8_csa_component_fa25_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa25_and1 = s_CSAwallace_rca24_csa13_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa25_or0 = s_CSAwallace_rca24_csa13_csa_component_fa25_and0 | s_CSAwallace_rca24_csa13_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa1_csa_component_fa26_xor1 ^ s_CSAwallace_rca24_csa8_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa26_and0 = s_CSAwallace_rca24_csa1_csa_component_fa26_xor1 & s_CSAwallace_rca24_csa8_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa13_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa26_and1 = s_CSAwallace_rca24_csa13_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa26_or0 = s_CSAwallace_rca24_csa13_csa_component_fa26_and0 | s_CSAwallace_rca24_csa13_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa27_xor0 = ~s_CSAwallace_rca24_csa1_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa27_and1 = s_CSAwallace_rca24_csa13_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa27_or0 = s_CSAwallace_rca24_csa1_csa_component_fa27_xor1 | s_CSAwallace_rca24_csa13_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa28_xor0 = ~s_CSAwallace_rca24_nand_23_5;
  assign s_CSAwallace_rca24_csa13_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa13_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa28_and1 = s_CSAwallace_rca24_csa13_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa13_csa_component_fa28_or0 = s_CSAwallace_rca24_nand_23_5 | s_CSAwallace_rca24_csa13_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa9_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa8_or0 ^ s_CSAwallace_rca24_and_0_9;
  assign s_CSAwallace_rca24_csa14_csa_component_fa9_and0 = s_CSAwallace_rca24_csa9_csa_component_fa8_or0 & s_CSAwallace_rca24_and_0_9;
  assign s_CSAwallace_rca24_csa14_csa_component_fa10_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa9_or0 ^ s_CSAwallace_rca24_csa3_csa_component_fa10_xor0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa10_and0 = s_CSAwallace_rca24_csa9_csa_component_fa9_or0 & s_CSAwallace_rca24_csa3_csa_component_fa10_xor0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa11_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa10_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa11_xor0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa11_and0 = s_CSAwallace_rca24_csa9_csa_component_fa10_or0 & s_CSAwallace_rca24_csa10_csa_component_fa11_xor0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa12_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa11_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa12_and0 = s_CSAwallace_rca24_csa9_csa_component_fa11_or0 & s_CSAwallace_rca24_csa10_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa11_and0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa12_and1 = s_CSAwallace_rca24_csa14_csa_component_fa12_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa11_and0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa12_or0 = s_CSAwallace_rca24_csa14_csa_component_fa12_and0 | s_CSAwallace_rca24_csa14_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa13_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa12_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa13_and0 = s_CSAwallace_rca24_csa9_csa_component_fa12_or0 & s_CSAwallace_rca24_csa10_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa13_and1 = s_CSAwallace_rca24_csa14_csa_component_fa13_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa13_or0 = s_CSAwallace_rca24_csa14_csa_component_fa13_and0 | s_CSAwallace_rca24_csa14_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa13_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa14_and0 = s_CSAwallace_rca24_csa9_csa_component_fa13_or0 & s_CSAwallace_rca24_csa10_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa14_and1 = s_CSAwallace_rca24_csa14_csa_component_fa14_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa14_or0 = s_CSAwallace_rca24_csa14_csa_component_fa14_and0 | s_CSAwallace_rca24_csa14_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa14_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa15_and0 = s_CSAwallace_rca24_csa9_csa_component_fa14_or0 & s_CSAwallace_rca24_csa10_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa15_and1 = s_CSAwallace_rca24_csa14_csa_component_fa15_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa15_or0 = s_CSAwallace_rca24_csa14_csa_component_fa15_and0 | s_CSAwallace_rca24_csa14_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa15_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa16_and0 = s_CSAwallace_rca24_csa9_csa_component_fa15_or0 & s_CSAwallace_rca24_csa10_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa16_and1 = s_CSAwallace_rca24_csa14_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa16_or0 = s_CSAwallace_rca24_csa14_csa_component_fa16_and0 | s_CSAwallace_rca24_csa14_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa16_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa17_and0 = s_CSAwallace_rca24_csa9_csa_component_fa16_or0 & s_CSAwallace_rca24_csa10_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa17_and1 = s_CSAwallace_rca24_csa14_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa17_or0 = s_CSAwallace_rca24_csa14_csa_component_fa17_and0 | s_CSAwallace_rca24_csa14_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa17_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa18_and0 = s_CSAwallace_rca24_csa9_csa_component_fa17_or0 & s_CSAwallace_rca24_csa10_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa18_and1 = s_CSAwallace_rca24_csa14_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa18_or0 = s_CSAwallace_rca24_csa14_csa_component_fa18_and0 | s_CSAwallace_rca24_csa14_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa18_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa19_and0 = s_CSAwallace_rca24_csa9_csa_component_fa18_or0 & s_CSAwallace_rca24_csa10_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa19_and1 = s_CSAwallace_rca24_csa14_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa19_or0 = s_CSAwallace_rca24_csa14_csa_component_fa19_and0 | s_CSAwallace_rca24_csa14_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa19_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa20_and0 = s_CSAwallace_rca24_csa9_csa_component_fa19_or0 & s_CSAwallace_rca24_csa10_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa20_and1 = s_CSAwallace_rca24_csa14_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa20_or0 = s_CSAwallace_rca24_csa14_csa_component_fa20_and0 | s_CSAwallace_rca24_csa14_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa20_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa21_and0 = s_CSAwallace_rca24_csa9_csa_component_fa20_or0 & s_CSAwallace_rca24_csa10_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa21_and1 = s_CSAwallace_rca24_csa14_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa21_or0 = s_CSAwallace_rca24_csa14_csa_component_fa21_and0 | s_CSAwallace_rca24_csa14_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa21_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa22_and0 = s_CSAwallace_rca24_csa9_csa_component_fa21_or0 & s_CSAwallace_rca24_csa10_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa22_and1 = s_CSAwallace_rca24_csa14_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa22_or0 = s_CSAwallace_rca24_csa14_csa_component_fa22_and0 | s_CSAwallace_rca24_csa14_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa22_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa23_and0 = s_CSAwallace_rca24_csa9_csa_component_fa22_or0 & s_CSAwallace_rca24_csa10_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa23_and1 = s_CSAwallace_rca24_csa14_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa23_or0 = s_CSAwallace_rca24_csa14_csa_component_fa23_and0 | s_CSAwallace_rca24_csa14_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa23_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa24_and0 = s_CSAwallace_rca24_csa9_csa_component_fa23_or0 & s_CSAwallace_rca24_csa10_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa24_and1 = s_CSAwallace_rca24_csa14_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa24_or0 = s_CSAwallace_rca24_csa14_csa_component_fa24_and0 | s_CSAwallace_rca24_csa14_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa24_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa25_and0 = s_CSAwallace_rca24_csa9_csa_component_fa24_or0 & s_CSAwallace_rca24_csa10_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa25_and1 = s_CSAwallace_rca24_csa14_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa25_or0 = s_CSAwallace_rca24_csa14_csa_component_fa25_and0 | s_CSAwallace_rca24_csa14_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa25_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa26_and0 = s_CSAwallace_rca24_csa9_csa_component_fa25_or0 & s_CSAwallace_rca24_csa10_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa26_and1 = s_CSAwallace_rca24_csa14_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa26_or0 = s_CSAwallace_rca24_csa14_csa_component_fa26_and0 | s_CSAwallace_rca24_csa14_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa26_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa27_and0 = s_CSAwallace_rca24_csa9_csa_component_fa26_or0 & s_CSAwallace_rca24_csa10_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa27_and1 = s_CSAwallace_rca24_csa14_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa27_or0 = s_CSAwallace_rca24_csa14_csa_component_fa27_and0 | s_CSAwallace_rca24_csa14_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa27_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa28_and0 = s_CSAwallace_rca24_csa9_csa_component_fa27_or0 & s_CSAwallace_rca24_csa10_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa28_and1 = s_CSAwallace_rca24_csa14_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa28_or0 = s_CSAwallace_rca24_csa14_csa_component_fa28_and0 | s_CSAwallace_rca24_csa14_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa28_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa29_and0 = s_CSAwallace_rca24_csa9_csa_component_fa28_or0 & s_CSAwallace_rca24_csa10_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa29_and1 = s_CSAwallace_rca24_csa14_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa29_or0 = s_CSAwallace_rca24_csa14_csa_component_fa29_and0 | s_CSAwallace_rca24_csa14_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa29_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa30_and0 = s_CSAwallace_rca24_csa9_csa_component_fa29_or0 & s_CSAwallace_rca24_csa10_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa30_and1 = s_CSAwallace_rca24_csa14_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa30_or0 = s_CSAwallace_rca24_csa14_csa_component_fa30_and0 | s_CSAwallace_rca24_csa14_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa30_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa31_and0 = s_CSAwallace_rca24_csa9_csa_component_fa30_or0 & s_CSAwallace_rca24_csa10_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa31_and1 = s_CSAwallace_rca24_csa14_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa31_or0 = s_CSAwallace_rca24_csa14_csa_component_fa31_and0 | s_CSAwallace_rca24_csa14_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa31_or0 ^ s_CSAwallace_rca24_csa10_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa32_and0 = s_CSAwallace_rca24_csa9_csa_component_fa31_or0 & s_CSAwallace_rca24_csa10_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa32_and1 = s_CSAwallace_rca24_csa14_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa32_or0 = s_CSAwallace_rca24_csa14_csa_component_fa32_and0 | s_CSAwallace_rca24_csa14_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa33_xor0 = ~s_CSAwallace_rca24_csa10_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa33_and1 = s_CSAwallace_rca24_csa14_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa33_or0 = s_CSAwallace_rca24_csa10_csa_component_fa33_xor1 | s_CSAwallace_rca24_csa14_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa34_xor0 = ~s_CSAwallace_rca24_csa10_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa34_and1 = s_CSAwallace_rca24_csa14_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa34_or0 = s_CSAwallace_rca24_csa10_csa_component_fa34_xor1 | s_CSAwallace_rca24_csa14_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa35_xor0 = ~s_CSAwallace_rca24_csa4_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa14_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_csa10_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa35_and1 = s_CSAwallace_rca24_csa14_csa_component_fa35_xor0 & s_CSAwallace_rca24_csa10_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa35_or0 = s_CSAwallace_rca24_csa4_csa_component_fa35_xor1 | s_CSAwallace_rca24_csa14_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa36_xor0 = ~s_CSAwallace_rca24_csa4_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa14_csa_component_fa36_xor1 = ~s_CSAwallace_rca24_csa14_csa_component_fa36_xor0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa36_or0 = s_CSAwallace_rca24_csa4_csa_component_fa36_xor1 | s_CSAwallace_rca24_csa14_csa_component_fa36_xor0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa37_xor0 = ~s_CSAwallace_rca24_nand_23_14;
  assign s_CSAwallace_rca24_csa14_csa_component_fa37_xor1 = ~s_CSAwallace_rca24_csa14_csa_component_fa37_xor0;
  assign s_CSAwallace_rca24_csa14_csa_component_fa37_or0 = s_CSAwallace_rca24_nand_23_14 | s_CSAwallace_rca24_csa14_csa_component_fa37_xor0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa11_csa_component_fa15_and0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa16_and0 = s_CSAwallace_rca24_csa11_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa11_csa_component_fa15_and0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa17_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa17_and0 = s_CSAwallace_rca24_csa11_csa_component_fa17_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa18_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa18_and0 = s_CSAwallace_rca24_csa11_csa_component_fa18_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_and_0_18;
  assign s_CSAwallace_rca24_csa15_csa_component_fa18_and1 = s_CSAwallace_rca24_csa15_csa_component_fa18_xor0 & s_CSAwallace_rca24_and_0_18;
  assign s_CSAwallace_rca24_csa15_csa_component_fa18_or0 = s_CSAwallace_rca24_csa15_csa_component_fa18_and0 | s_CSAwallace_rca24_csa15_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa19_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa19_and0 = s_CSAwallace_rca24_csa11_csa_component_fa19_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa6_csa_component_fa19_xor0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa19_and1 = s_CSAwallace_rca24_csa15_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa6_csa_component_fa19_xor0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa19_or0 = s_CSAwallace_rca24_csa15_csa_component_fa19_and0 | s_CSAwallace_rca24_csa15_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa20_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa20_and0 = s_CSAwallace_rca24_csa11_csa_component_fa20_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa20_xor0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa20_and1 = s_CSAwallace_rca24_csa15_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa20_xor0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa20_or0 = s_CSAwallace_rca24_csa15_csa_component_fa20_and0 | s_CSAwallace_rca24_csa15_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa21_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa21_and0 = s_CSAwallace_rca24_csa11_csa_component_fa21_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa21_and1 = s_CSAwallace_rca24_csa15_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa21_or0 = s_CSAwallace_rca24_csa15_csa_component_fa21_and0 | s_CSAwallace_rca24_csa15_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa22_and0 = s_CSAwallace_rca24_csa11_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa22_and1 = s_CSAwallace_rca24_csa15_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa22_or0 = s_CSAwallace_rca24_csa15_csa_component_fa22_and0 | s_CSAwallace_rca24_csa15_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa23_and0 = s_CSAwallace_rca24_csa11_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa23_and1 = s_CSAwallace_rca24_csa15_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa23_or0 = s_CSAwallace_rca24_csa15_csa_component_fa23_and0 | s_CSAwallace_rca24_csa15_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa24_and0 = s_CSAwallace_rca24_csa11_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa24_and1 = s_CSAwallace_rca24_csa15_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa24_or0 = s_CSAwallace_rca24_csa15_csa_component_fa24_and0 | s_CSAwallace_rca24_csa15_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa25_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa25_and0 = s_CSAwallace_rca24_csa11_csa_component_fa25_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa25_and1 = s_CSAwallace_rca24_csa15_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa25_or0 = s_CSAwallace_rca24_csa15_csa_component_fa25_and0 | s_CSAwallace_rca24_csa15_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa26_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa26_and0 = s_CSAwallace_rca24_csa11_csa_component_fa26_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa26_and1 = s_CSAwallace_rca24_csa15_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa26_or0 = s_CSAwallace_rca24_csa15_csa_component_fa26_and0 | s_CSAwallace_rca24_csa15_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa27_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa27_and0 = s_CSAwallace_rca24_csa11_csa_component_fa27_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa27_and1 = s_CSAwallace_rca24_csa15_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa27_or0 = s_CSAwallace_rca24_csa15_csa_component_fa27_and0 | s_CSAwallace_rca24_csa15_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa28_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa28_and0 = s_CSAwallace_rca24_csa11_csa_component_fa28_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa28_and1 = s_CSAwallace_rca24_csa15_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa28_or0 = s_CSAwallace_rca24_csa15_csa_component_fa28_and0 | s_CSAwallace_rca24_csa15_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa29_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa29_and0 = s_CSAwallace_rca24_csa11_csa_component_fa29_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa29_and1 = s_CSAwallace_rca24_csa15_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa29_or0 = s_CSAwallace_rca24_csa15_csa_component_fa29_and0 | s_CSAwallace_rca24_csa15_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa30_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa30_and0 = s_CSAwallace_rca24_csa11_csa_component_fa30_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa30_and1 = s_CSAwallace_rca24_csa15_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa30_or0 = s_CSAwallace_rca24_csa15_csa_component_fa30_and0 | s_CSAwallace_rca24_csa15_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa31_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa31_and0 = s_CSAwallace_rca24_csa11_csa_component_fa31_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa31_and1 = s_CSAwallace_rca24_csa15_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa31_or0 = s_CSAwallace_rca24_csa15_csa_component_fa31_and0 | s_CSAwallace_rca24_csa15_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa32_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa32_and0 = s_CSAwallace_rca24_csa11_csa_component_fa32_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa32_and1 = s_CSAwallace_rca24_csa15_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa32_or0 = s_CSAwallace_rca24_csa15_csa_component_fa32_and0 | s_CSAwallace_rca24_csa15_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa33_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa33_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa33_and0 = s_CSAwallace_rca24_csa11_csa_component_fa33_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa33_and1 = s_CSAwallace_rca24_csa15_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa33_or0 = s_CSAwallace_rca24_csa15_csa_component_fa33_and0 | s_CSAwallace_rca24_csa15_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa34_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa34_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa34_and0 = s_CSAwallace_rca24_csa11_csa_component_fa34_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa34_and1 = s_CSAwallace_rca24_csa15_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa34_or0 = s_CSAwallace_rca24_csa15_csa_component_fa34_and0 | s_CSAwallace_rca24_csa15_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa35_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa35_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa35_and0 = s_CSAwallace_rca24_csa11_csa_component_fa35_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa35_and1 = s_CSAwallace_rca24_csa15_csa_component_fa35_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa35_or0 = s_CSAwallace_rca24_csa15_csa_component_fa35_and0 | s_CSAwallace_rca24_csa15_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa36_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa36_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa36_and0 = s_CSAwallace_rca24_csa11_csa_component_fa36_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa36_and1 = s_CSAwallace_rca24_csa15_csa_component_fa36_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa36_or0 = s_CSAwallace_rca24_csa15_csa_component_fa36_and0 | s_CSAwallace_rca24_csa15_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa37_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa37_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa37_and0 = s_CSAwallace_rca24_csa11_csa_component_fa37_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa37_and1 = s_CSAwallace_rca24_csa15_csa_component_fa37_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa37_or0 = s_CSAwallace_rca24_csa15_csa_component_fa37_and0 | s_CSAwallace_rca24_csa15_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa38_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa38_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa38_and0 = s_CSAwallace_rca24_csa11_csa_component_fa38_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa38_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa38_and1 = s_CSAwallace_rca24_csa15_csa_component_fa38_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa38_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa38_or0 = s_CSAwallace_rca24_csa15_csa_component_fa38_and0 | s_CSAwallace_rca24_csa15_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa39_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa39_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa39_and0 = s_CSAwallace_rca24_csa11_csa_component_fa39_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa39_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa39_and1 = s_CSAwallace_rca24_csa15_csa_component_fa39_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa39_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa39_or0 = s_CSAwallace_rca24_csa15_csa_component_fa39_and0 | s_CSAwallace_rca24_csa15_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa40_xor0 = s_CSAwallace_rca24_csa11_csa_component_fa40_xor1 ^ s_CSAwallace_rca24_csa11_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa40_and0 = s_CSAwallace_rca24_csa11_csa_component_fa40_xor1 & s_CSAwallace_rca24_csa11_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa40_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa40_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa40_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa40_and1 = s_CSAwallace_rca24_csa15_csa_component_fa40_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa40_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa40_or0 = s_CSAwallace_rca24_csa15_csa_component_fa40_and0 | s_CSAwallace_rca24_csa15_csa_component_fa40_and1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa41_xor0 = ~s_CSAwallace_rca24_csa11_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa15_csa_component_fa41_xor1 = s_CSAwallace_rca24_csa15_csa_component_fa41_xor0 ^ s_CSAwallace_rca24_csa12_csa_component_fa41_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa41_and1 = s_CSAwallace_rca24_csa15_csa_component_fa41_xor0 & s_CSAwallace_rca24_csa12_csa_component_fa41_xor1;
  assign s_CSAwallace_rca24_csa15_csa_component_fa41_or0 = s_CSAwallace_rca24_csa11_csa_component_fa40_or0 | s_CSAwallace_rca24_csa15_csa_component_fa41_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa4_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa4_xor0 ^ s_CSAwallace_rca24_csa13_csa_component_fa3_and0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa4_and0 = s_CSAwallace_rca24_csa13_csa_component_fa4_xor0 & s_CSAwallace_rca24_csa13_csa_component_fa3_and0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa5_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa5_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa4_and0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa5_and0 = s_CSAwallace_rca24_csa13_csa_component_fa5_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa4_and0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa6_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa6_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa5_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa6_and0 = s_CSAwallace_rca24_csa13_csa_component_fa6_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa5_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa7_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa7_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa6_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa7_and0 = s_CSAwallace_rca24_csa13_csa_component_fa7_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa6_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa7_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa7_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa6_and0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa7_and1 = s_CSAwallace_rca24_csa16_csa_component_fa7_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa6_and0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa7_or0 = s_CSAwallace_rca24_csa16_csa_component_fa7_and0 | s_CSAwallace_rca24_csa16_csa_component_fa7_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa8_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa8_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa7_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa8_and0 = s_CSAwallace_rca24_csa13_csa_component_fa8_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa7_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa8_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_csa9_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa8_and1 = s_CSAwallace_rca24_csa16_csa_component_fa8_xor0 & s_CSAwallace_rca24_csa9_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa8_or0 = s_CSAwallace_rca24_csa16_csa_component_fa8_and0 | s_CSAwallace_rca24_csa16_csa_component_fa8_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa9_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa9_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa9_and0 = s_CSAwallace_rca24_csa13_csa_component_fa9_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa9_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa9_xor0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa9_and1 = s_CSAwallace_rca24_csa16_csa_component_fa9_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa9_xor0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa9_or0 = s_CSAwallace_rca24_csa16_csa_component_fa9_and0 | s_CSAwallace_rca24_csa16_csa_component_fa9_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa10_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa10_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa10_and0 = s_CSAwallace_rca24_csa13_csa_component_fa10_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa10_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa10_xor0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa10_and1 = s_CSAwallace_rca24_csa16_csa_component_fa10_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa10_xor0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa10_or0 = s_CSAwallace_rca24_csa16_csa_component_fa10_and0 | s_CSAwallace_rca24_csa16_csa_component_fa10_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa11_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa11_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa11_and0 = s_CSAwallace_rca24_csa13_csa_component_fa11_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa11_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa11_xor0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa11_and1 = s_CSAwallace_rca24_csa16_csa_component_fa11_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa11_xor0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa11_or0 = s_CSAwallace_rca24_csa16_csa_component_fa11_and0 | s_CSAwallace_rca24_csa16_csa_component_fa11_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa12_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa12_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa12_and0 = s_CSAwallace_rca24_csa13_csa_component_fa12_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa12_and1 = s_CSAwallace_rca24_csa16_csa_component_fa12_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa12_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa12_or0 = s_CSAwallace_rca24_csa16_csa_component_fa12_and0 | s_CSAwallace_rca24_csa16_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa13_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa13_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa13_and0 = s_CSAwallace_rca24_csa13_csa_component_fa13_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa13_and1 = s_CSAwallace_rca24_csa16_csa_component_fa13_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa13_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa13_or0 = s_CSAwallace_rca24_csa16_csa_component_fa13_and0 | s_CSAwallace_rca24_csa16_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa14_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa14_and0 = s_CSAwallace_rca24_csa13_csa_component_fa14_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa14_and1 = s_CSAwallace_rca24_csa16_csa_component_fa14_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa14_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa14_or0 = s_CSAwallace_rca24_csa16_csa_component_fa14_and0 | s_CSAwallace_rca24_csa16_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa15_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa15_and0 = s_CSAwallace_rca24_csa13_csa_component_fa15_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa15_and1 = s_CSAwallace_rca24_csa16_csa_component_fa15_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa15_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa15_or0 = s_CSAwallace_rca24_csa16_csa_component_fa15_and0 | s_CSAwallace_rca24_csa16_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa16_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa16_and0 = s_CSAwallace_rca24_csa13_csa_component_fa16_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa16_and1 = s_CSAwallace_rca24_csa16_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa16_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa16_or0 = s_CSAwallace_rca24_csa16_csa_component_fa16_and0 | s_CSAwallace_rca24_csa16_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa17_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa17_and0 = s_CSAwallace_rca24_csa13_csa_component_fa17_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa17_and1 = s_CSAwallace_rca24_csa16_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa17_or0 = s_CSAwallace_rca24_csa16_csa_component_fa17_and0 | s_CSAwallace_rca24_csa16_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa18_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa18_and0 = s_CSAwallace_rca24_csa13_csa_component_fa18_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa18_and1 = s_CSAwallace_rca24_csa16_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa18_or0 = s_CSAwallace_rca24_csa16_csa_component_fa18_and0 | s_CSAwallace_rca24_csa16_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa19_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa19_and0 = s_CSAwallace_rca24_csa13_csa_component_fa19_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa19_and1 = s_CSAwallace_rca24_csa16_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa19_or0 = s_CSAwallace_rca24_csa16_csa_component_fa19_and0 | s_CSAwallace_rca24_csa16_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa20_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa20_and0 = s_CSAwallace_rca24_csa13_csa_component_fa20_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa20_and1 = s_CSAwallace_rca24_csa16_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa20_or0 = s_CSAwallace_rca24_csa16_csa_component_fa20_and0 | s_CSAwallace_rca24_csa16_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa21_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa21_and0 = s_CSAwallace_rca24_csa13_csa_component_fa21_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa21_and1 = s_CSAwallace_rca24_csa16_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa21_or0 = s_CSAwallace_rca24_csa16_csa_component_fa21_and0 | s_CSAwallace_rca24_csa16_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa22_and0 = s_CSAwallace_rca24_csa13_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa22_and1 = s_CSAwallace_rca24_csa16_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa22_or0 = s_CSAwallace_rca24_csa16_csa_component_fa22_and0 | s_CSAwallace_rca24_csa16_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa23_and0 = s_CSAwallace_rca24_csa13_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa23_and1 = s_CSAwallace_rca24_csa16_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa23_or0 = s_CSAwallace_rca24_csa16_csa_component_fa23_and0 | s_CSAwallace_rca24_csa16_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa24_and0 = s_CSAwallace_rca24_csa13_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa24_and1 = s_CSAwallace_rca24_csa16_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa24_or0 = s_CSAwallace_rca24_csa16_csa_component_fa24_and0 | s_CSAwallace_rca24_csa16_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa25_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa25_and0 = s_CSAwallace_rca24_csa13_csa_component_fa25_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa25_and1 = s_CSAwallace_rca24_csa16_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa25_or0 = s_CSAwallace_rca24_csa16_csa_component_fa25_and0 | s_CSAwallace_rca24_csa16_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa26_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa26_and0 = s_CSAwallace_rca24_csa13_csa_component_fa26_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa26_and1 = s_CSAwallace_rca24_csa16_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa26_or0 = s_CSAwallace_rca24_csa16_csa_component_fa26_and0 | s_CSAwallace_rca24_csa16_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa27_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa27_and0 = s_CSAwallace_rca24_csa13_csa_component_fa27_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa27_and1 = s_CSAwallace_rca24_csa16_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa27_or0 = s_CSAwallace_rca24_csa16_csa_component_fa27_and0 | s_CSAwallace_rca24_csa16_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa13_csa_component_fa28_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa28_and0 = s_CSAwallace_rca24_csa13_csa_component_fa28_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa28_and1 = s_CSAwallace_rca24_csa16_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa28_or0 = s_CSAwallace_rca24_csa16_csa_component_fa28_and0 | s_CSAwallace_rca24_csa16_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa9_csa_component_fa29_xor1 ^ s_CSAwallace_rca24_csa13_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa29_and0 = s_CSAwallace_rca24_csa9_csa_component_fa29_xor1 & s_CSAwallace_rca24_csa13_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa16_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa29_and1 = s_CSAwallace_rca24_csa16_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa29_or0 = s_CSAwallace_rca24_csa16_csa_component_fa29_and0 | s_CSAwallace_rca24_csa16_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa30_xor0 = ~s_CSAwallace_rca24_csa9_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa30_and1 = s_CSAwallace_rca24_csa16_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa30_or0 = s_CSAwallace_rca24_csa9_csa_component_fa30_xor1 | s_CSAwallace_rca24_csa16_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa31_xor0 = ~s_CSAwallace_rca24_csa9_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa16_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa31_and1 = s_CSAwallace_rca24_csa16_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa16_csa_component_fa31_or0 = s_CSAwallace_rca24_csa9_csa_component_fa31_xor1 | s_CSAwallace_rca24_csa16_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa13_or0 ^ s_CSAwallace_rca24_csa4_csa_component_fa13_and0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa14_and0 = s_CSAwallace_rca24_csa14_csa_component_fa13_or0 & s_CSAwallace_rca24_csa4_csa_component_fa13_and0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa14_or0 ^ s_CSAwallace_rca24_csa11_csa_component_fa15_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa15_and0 = s_CSAwallace_rca24_csa14_csa_component_fa14_or0 & s_CSAwallace_rca24_csa11_csa_component_fa15_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa15_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa16_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa16_and0 = s_CSAwallace_rca24_csa14_csa_component_fa15_or0 & s_CSAwallace_rca24_csa15_csa_component_fa16_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa16_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa17_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa17_and0 = s_CSAwallace_rca24_csa14_csa_component_fa16_or0 & s_CSAwallace_rca24_csa15_csa_component_fa17_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa17_and1 = s_CSAwallace_rca24_csa17_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa17_or0 = s_CSAwallace_rca24_csa17_csa_component_fa17_and0 | s_CSAwallace_rca24_csa17_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa17_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa18_and0 = s_CSAwallace_rca24_csa14_csa_component_fa17_or0 & s_CSAwallace_rca24_csa15_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa17_and0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa18_and1 = s_CSAwallace_rca24_csa17_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa17_and0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa18_or0 = s_CSAwallace_rca24_csa17_csa_component_fa18_and0 | s_CSAwallace_rca24_csa17_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa18_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa19_and0 = s_CSAwallace_rca24_csa14_csa_component_fa18_or0 & s_CSAwallace_rca24_csa15_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa19_and1 = s_CSAwallace_rca24_csa17_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa19_or0 = s_CSAwallace_rca24_csa17_csa_component_fa19_and0 | s_CSAwallace_rca24_csa17_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa19_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa20_and0 = s_CSAwallace_rca24_csa14_csa_component_fa19_or0 & s_CSAwallace_rca24_csa15_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa20_and1 = s_CSAwallace_rca24_csa17_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa20_or0 = s_CSAwallace_rca24_csa17_csa_component_fa20_and0 | s_CSAwallace_rca24_csa17_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa20_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa21_and0 = s_CSAwallace_rca24_csa14_csa_component_fa20_or0 & s_CSAwallace_rca24_csa15_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa21_and1 = s_CSAwallace_rca24_csa17_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa21_or0 = s_CSAwallace_rca24_csa17_csa_component_fa21_and0 | s_CSAwallace_rca24_csa17_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa21_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa22_and0 = s_CSAwallace_rca24_csa14_csa_component_fa21_or0 & s_CSAwallace_rca24_csa15_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa22_and1 = s_CSAwallace_rca24_csa17_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa22_or0 = s_CSAwallace_rca24_csa17_csa_component_fa22_and0 | s_CSAwallace_rca24_csa17_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa22_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa23_and0 = s_CSAwallace_rca24_csa14_csa_component_fa22_or0 & s_CSAwallace_rca24_csa15_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa23_and1 = s_CSAwallace_rca24_csa17_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa23_or0 = s_CSAwallace_rca24_csa17_csa_component_fa23_and0 | s_CSAwallace_rca24_csa17_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa23_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa24_and0 = s_CSAwallace_rca24_csa14_csa_component_fa23_or0 & s_CSAwallace_rca24_csa15_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa24_and1 = s_CSAwallace_rca24_csa17_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa24_or0 = s_CSAwallace_rca24_csa17_csa_component_fa24_and0 | s_CSAwallace_rca24_csa17_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa24_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa25_and0 = s_CSAwallace_rca24_csa14_csa_component_fa24_or0 & s_CSAwallace_rca24_csa15_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa25_and1 = s_CSAwallace_rca24_csa17_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa25_or0 = s_CSAwallace_rca24_csa17_csa_component_fa25_and0 | s_CSAwallace_rca24_csa17_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa25_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa26_and0 = s_CSAwallace_rca24_csa14_csa_component_fa25_or0 & s_CSAwallace_rca24_csa15_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa26_and1 = s_CSAwallace_rca24_csa17_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa26_or0 = s_CSAwallace_rca24_csa17_csa_component_fa26_and0 | s_CSAwallace_rca24_csa17_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa26_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa27_and0 = s_CSAwallace_rca24_csa14_csa_component_fa26_or0 & s_CSAwallace_rca24_csa15_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa27_and1 = s_CSAwallace_rca24_csa17_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa27_or0 = s_CSAwallace_rca24_csa17_csa_component_fa27_and0 | s_CSAwallace_rca24_csa17_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa27_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa28_and0 = s_CSAwallace_rca24_csa14_csa_component_fa27_or0 & s_CSAwallace_rca24_csa15_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa28_and1 = s_CSAwallace_rca24_csa17_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa28_or0 = s_CSAwallace_rca24_csa17_csa_component_fa28_and0 | s_CSAwallace_rca24_csa17_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa28_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa29_and0 = s_CSAwallace_rca24_csa14_csa_component_fa28_or0 & s_CSAwallace_rca24_csa15_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa29_and1 = s_CSAwallace_rca24_csa17_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa29_or0 = s_CSAwallace_rca24_csa17_csa_component_fa29_and0 | s_CSAwallace_rca24_csa17_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa29_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa30_and0 = s_CSAwallace_rca24_csa14_csa_component_fa29_or0 & s_CSAwallace_rca24_csa15_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa30_and1 = s_CSAwallace_rca24_csa17_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa30_or0 = s_CSAwallace_rca24_csa17_csa_component_fa30_and0 | s_CSAwallace_rca24_csa17_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa30_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa31_and0 = s_CSAwallace_rca24_csa14_csa_component_fa30_or0 & s_CSAwallace_rca24_csa15_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa31_and1 = s_CSAwallace_rca24_csa17_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa31_or0 = s_CSAwallace_rca24_csa17_csa_component_fa31_and0 | s_CSAwallace_rca24_csa17_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa31_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa32_and0 = s_CSAwallace_rca24_csa14_csa_component_fa31_or0 & s_CSAwallace_rca24_csa15_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa32_and1 = s_CSAwallace_rca24_csa17_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa32_or0 = s_CSAwallace_rca24_csa17_csa_component_fa32_and0 | s_CSAwallace_rca24_csa17_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa33_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa32_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa33_and0 = s_CSAwallace_rca24_csa14_csa_component_fa32_or0 & s_CSAwallace_rca24_csa15_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa33_and1 = s_CSAwallace_rca24_csa17_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa33_or0 = s_CSAwallace_rca24_csa17_csa_component_fa33_and0 | s_CSAwallace_rca24_csa17_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa34_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa33_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa34_and0 = s_CSAwallace_rca24_csa14_csa_component_fa33_or0 & s_CSAwallace_rca24_csa15_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa34_and1 = s_CSAwallace_rca24_csa17_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa34_or0 = s_CSAwallace_rca24_csa17_csa_component_fa34_and0 | s_CSAwallace_rca24_csa17_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa35_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa34_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa35_and0 = s_CSAwallace_rca24_csa14_csa_component_fa34_or0 & s_CSAwallace_rca24_csa15_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa35_and1 = s_CSAwallace_rca24_csa17_csa_component_fa35_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa35_or0 = s_CSAwallace_rca24_csa17_csa_component_fa35_and0 | s_CSAwallace_rca24_csa17_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa36_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa35_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa36_and0 = s_CSAwallace_rca24_csa14_csa_component_fa35_or0 & s_CSAwallace_rca24_csa15_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa36_and1 = s_CSAwallace_rca24_csa17_csa_component_fa36_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa36_or0 = s_CSAwallace_rca24_csa17_csa_component_fa36_and0 | s_CSAwallace_rca24_csa17_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa37_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa36_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa37_and0 = s_CSAwallace_rca24_csa14_csa_component_fa36_or0 & s_CSAwallace_rca24_csa15_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa37_and1 = s_CSAwallace_rca24_csa17_csa_component_fa37_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa37_or0 = s_CSAwallace_rca24_csa17_csa_component_fa37_and0 | s_CSAwallace_rca24_csa17_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa38_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa37_or0 ^ s_CSAwallace_rca24_csa15_csa_component_fa38_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa38_and0 = s_CSAwallace_rca24_csa14_csa_component_fa37_or0 & s_CSAwallace_rca24_csa15_csa_component_fa38_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa38_and1 = s_CSAwallace_rca24_csa17_csa_component_fa38_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa38_or0 = s_CSAwallace_rca24_csa17_csa_component_fa38_and0 | s_CSAwallace_rca24_csa17_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa39_xor0 = ~s_CSAwallace_rca24_csa15_csa_component_fa39_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa39_and1 = s_CSAwallace_rca24_csa17_csa_component_fa39_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa39_or0 = s_CSAwallace_rca24_csa15_csa_component_fa39_xor1 | s_CSAwallace_rca24_csa17_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa40_xor0 = ~s_CSAwallace_rca24_csa15_csa_component_fa40_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa40_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa40_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa40_and1 = s_CSAwallace_rca24_csa17_csa_component_fa40_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa40_or0 = s_CSAwallace_rca24_csa15_csa_component_fa40_xor1 | s_CSAwallace_rca24_csa17_csa_component_fa40_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa41_xor0 = ~s_CSAwallace_rca24_csa15_csa_component_fa41_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa41_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa41_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa41_and1 = s_CSAwallace_rca24_csa17_csa_component_fa41_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa41_or0 = s_CSAwallace_rca24_csa15_csa_component_fa41_xor1 | s_CSAwallace_rca24_csa17_csa_component_fa41_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa42_xor0 = ~s_CSAwallace_rca24_csa12_csa_component_fa42_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa42_xor1 = s_CSAwallace_rca24_csa17_csa_component_fa42_xor0 ^ s_CSAwallace_rca24_csa15_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa42_and1 = s_CSAwallace_rca24_csa17_csa_component_fa42_xor0 & s_CSAwallace_rca24_csa15_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa42_or0 = s_CSAwallace_rca24_csa12_csa_component_fa42_xor1 | s_CSAwallace_rca24_csa17_csa_component_fa42_and1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa43_xor0 = ~s_CSAwallace_rca24_csa12_csa_component_fa43_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa43_xor1 = ~s_CSAwallace_rca24_csa17_csa_component_fa43_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa43_or0 = s_CSAwallace_rca24_csa12_csa_component_fa43_xor1 | s_CSAwallace_rca24_csa17_csa_component_fa43_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa44_xor0 = ~s_CSAwallace_rca24_csa7_csa_component_fa44_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa44_xor1 = ~s_CSAwallace_rca24_csa17_csa_component_fa44_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa44_or0 = s_CSAwallace_rca24_csa7_csa_component_fa44_xor1 | s_CSAwallace_rca24_csa17_csa_component_fa44_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa45_xor0 = ~s_CSAwallace_rca24_csa7_csa_component_fa45_xor1;
  assign s_CSAwallace_rca24_csa17_csa_component_fa45_xor1 = ~s_CSAwallace_rca24_csa17_csa_component_fa45_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa45_or0 = s_CSAwallace_rca24_csa7_csa_component_fa45_xor1 | s_CSAwallace_rca24_csa17_csa_component_fa45_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa46_xor0 = ~s_CSAwallace_rca24_and_23_23;
  assign s_CSAwallace_rca24_csa17_csa_component_fa46_xor1 = ~s_CSAwallace_rca24_csa17_csa_component_fa46_xor0;
  assign s_CSAwallace_rca24_csa17_csa_component_fa46_or0 = s_CSAwallace_rca24_and_23_23 | s_CSAwallace_rca24_csa17_csa_component_fa46_xor0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa5_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa5_xor0 ^ s_CSAwallace_rca24_csa16_csa_component_fa4_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa5_and0 = s_CSAwallace_rca24_csa16_csa_component_fa5_xor0 & s_CSAwallace_rca24_csa16_csa_component_fa4_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa6_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa6_xor0 ^ s_CSAwallace_rca24_csa16_csa_component_fa5_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa6_and0 = s_CSAwallace_rca24_csa16_csa_component_fa6_xor0 & s_CSAwallace_rca24_csa16_csa_component_fa5_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa7_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa7_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa6_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa7_and0 = s_CSAwallace_rca24_csa16_csa_component_fa7_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa6_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa8_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa8_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa7_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa8_and0 = s_CSAwallace_rca24_csa16_csa_component_fa8_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa7_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa9_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa9_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa9_and0 = s_CSAwallace_rca24_csa16_csa_component_fa9_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa8_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa10_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa10_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa10_and0 = s_CSAwallace_rca24_csa16_csa_component_fa10_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa9_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa10_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa9_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa10_and1 = s_CSAwallace_rca24_csa18_csa_component_fa10_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa9_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa10_or0 = s_CSAwallace_rca24_csa18_csa_component_fa10_and0 | s_CSAwallace_rca24_csa18_csa_component_fa10_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa11_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa11_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa11_and0 = s_CSAwallace_rca24_csa16_csa_component_fa11_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa11_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa10_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa11_and1 = s_CSAwallace_rca24_csa18_csa_component_fa11_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa10_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa11_or0 = s_CSAwallace_rca24_csa18_csa_component_fa11_and0 | s_CSAwallace_rca24_csa18_csa_component_fa11_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa12_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa12_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa12_and0 = s_CSAwallace_rca24_csa16_csa_component_fa12_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa12_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa11_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa12_and1 = s_CSAwallace_rca24_csa18_csa_component_fa12_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa11_and0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa12_or0 = s_CSAwallace_rca24_csa18_csa_component_fa12_and0 | s_CSAwallace_rca24_csa18_csa_component_fa12_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa13_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa13_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa13_and0 = s_CSAwallace_rca24_csa16_csa_component_fa13_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa13_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_csa14_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa13_and1 = s_CSAwallace_rca24_csa18_csa_component_fa13_xor0 & s_CSAwallace_rca24_csa14_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa13_or0 = s_CSAwallace_rca24_csa18_csa_component_fa13_and0 | s_CSAwallace_rca24_csa18_csa_component_fa13_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa14_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa14_and0 = s_CSAwallace_rca24_csa16_csa_component_fa14_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa14_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa14_xor0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa14_and1 = s_CSAwallace_rca24_csa18_csa_component_fa14_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa14_xor0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa14_or0 = s_CSAwallace_rca24_csa18_csa_component_fa14_and0 | s_CSAwallace_rca24_csa18_csa_component_fa14_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa15_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa15_and0 = s_CSAwallace_rca24_csa16_csa_component_fa15_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa15_xor0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa15_and1 = s_CSAwallace_rca24_csa18_csa_component_fa15_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa15_xor0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa15_or0 = s_CSAwallace_rca24_csa18_csa_component_fa15_and0 | s_CSAwallace_rca24_csa18_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa16_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa16_and0 = s_CSAwallace_rca24_csa16_csa_component_fa16_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa16_xor0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa16_and1 = s_CSAwallace_rca24_csa18_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa16_xor0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa16_or0 = s_CSAwallace_rca24_csa18_csa_component_fa16_and0 | s_CSAwallace_rca24_csa18_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa17_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa17_and0 = s_CSAwallace_rca24_csa16_csa_component_fa17_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa17_and1 = s_CSAwallace_rca24_csa18_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa17_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa17_or0 = s_CSAwallace_rca24_csa18_csa_component_fa17_and0 | s_CSAwallace_rca24_csa18_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa18_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa18_and0 = s_CSAwallace_rca24_csa16_csa_component_fa18_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa18_and1 = s_CSAwallace_rca24_csa18_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa18_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa18_or0 = s_CSAwallace_rca24_csa18_csa_component_fa18_and0 | s_CSAwallace_rca24_csa18_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa19_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa19_and0 = s_CSAwallace_rca24_csa16_csa_component_fa19_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa19_and1 = s_CSAwallace_rca24_csa18_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa19_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa19_or0 = s_CSAwallace_rca24_csa18_csa_component_fa19_and0 | s_CSAwallace_rca24_csa18_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa20_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa20_and0 = s_CSAwallace_rca24_csa16_csa_component_fa20_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa20_and1 = s_CSAwallace_rca24_csa18_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa20_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa20_or0 = s_CSAwallace_rca24_csa18_csa_component_fa20_and0 | s_CSAwallace_rca24_csa18_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa21_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa21_and0 = s_CSAwallace_rca24_csa16_csa_component_fa21_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa21_and1 = s_CSAwallace_rca24_csa18_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa21_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa21_or0 = s_CSAwallace_rca24_csa18_csa_component_fa21_and0 | s_CSAwallace_rca24_csa18_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa22_and0 = s_CSAwallace_rca24_csa16_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa22_and1 = s_CSAwallace_rca24_csa18_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa22_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa22_or0 = s_CSAwallace_rca24_csa18_csa_component_fa22_and0 | s_CSAwallace_rca24_csa18_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa23_and0 = s_CSAwallace_rca24_csa16_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa23_and1 = s_CSAwallace_rca24_csa18_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa23_or0 = s_CSAwallace_rca24_csa18_csa_component_fa23_and0 | s_CSAwallace_rca24_csa18_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa24_and0 = s_CSAwallace_rca24_csa16_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa24_and1 = s_CSAwallace_rca24_csa18_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa24_or0 = s_CSAwallace_rca24_csa18_csa_component_fa24_and0 | s_CSAwallace_rca24_csa18_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa25_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa25_and0 = s_CSAwallace_rca24_csa16_csa_component_fa25_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa25_and1 = s_CSAwallace_rca24_csa18_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa25_or0 = s_CSAwallace_rca24_csa18_csa_component_fa25_and0 | s_CSAwallace_rca24_csa18_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa26_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa26_and0 = s_CSAwallace_rca24_csa16_csa_component_fa26_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa26_and1 = s_CSAwallace_rca24_csa18_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa26_or0 = s_CSAwallace_rca24_csa18_csa_component_fa26_and0 | s_CSAwallace_rca24_csa18_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa27_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa27_and0 = s_CSAwallace_rca24_csa16_csa_component_fa27_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa27_and1 = s_CSAwallace_rca24_csa18_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa27_or0 = s_CSAwallace_rca24_csa18_csa_component_fa27_and0 | s_CSAwallace_rca24_csa18_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa28_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa28_and0 = s_CSAwallace_rca24_csa16_csa_component_fa28_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa28_and1 = s_CSAwallace_rca24_csa18_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa28_or0 = s_CSAwallace_rca24_csa18_csa_component_fa28_and0 | s_CSAwallace_rca24_csa18_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa29_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa29_and0 = s_CSAwallace_rca24_csa16_csa_component_fa29_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa29_and1 = s_CSAwallace_rca24_csa18_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa29_or0 = s_CSAwallace_rca24_csa18_csa_component_fa29_and0 | s_CSAwallace_rca24_csa18_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa30_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa30_and0 = s_CSAwallace_rca24_csa16_csa_component_fa30_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa30_and1 = s_CSAwallace_rca24_csa18_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa30_or0 = s_CSAwallace_rca24_csa18_csa_component_fa30_and0 | s_CSAwallace_rca24_csa18_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa16_csa_component_fa31_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa31_and0 = s_CSAwallace_rca24_csa16_csa_component_fa31_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa31_and1 = s_CSAwallace_rca24_csa18_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa31_or0 = s_CSAwallace_rca24_csa18_csa_component_fa31_and0 | s_CSAwallace_rca24_csa18_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa14_csa_component_fa32_xor1 ^ s_CSAwallace_rca24_csa16_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa32_and0 = s_CSAwallace_rca24_csa14_csa_component_fa32_xor1 & s_CSAwallace_rca24_csa16_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa18_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa32_and1 = s_CSAwallace_rca24_csa18_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa32_or0 = s_CSAwallace_rca24_csa18_csa_component_fa32_and0 | s_CSAwallace_rca24_csa18_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa33_xor0 = ~s_CSAwallace_rca24_csa14_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa33_and1 = s_CSAwallace_rca24_csa18_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa33_or0 = s_CSAwallace_rca24_csa14_csa_component_fa33_xor1 | s_CSAwallace_rca24_csa18_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa34_xor0 = ~s_CSAwallace_rca24_csa14_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa34_and1 = s_CSAwallace_rca24_csa18_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa34_or0 = s_CSAwallace_rca24_csa14_csa_component_fa34_xor1 | s_CSAwallace_rca24_csa18_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa35_xor0 = ~s_CSAwallace_rca24_csa14_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa35_and1 = s_CSAwallace_rca24_csa18_csa_component_fa35_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa35_or0 = s_CSAwallace_rca24_csa14_csa_component_fa35_xor1 | s_CSAwallace_rca24_csa18_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa36_xor0 = ~s_CSAwallace_rca24_csa14_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa36_and1 = s_CSAwallace_rca24_csa18_csa_component_fa36_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa36_or0 = s_CSAwallace_rca24_csa14_csa_component_fa36_xor1 | s_CSAwallace_rca24_csa18_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa37_xor0 = ~s_CSAwallace_rca24_csa14_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa18_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa37_and1 = s_CSAwallace_rca24_csa18_csa_component_fa37_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa18_csa_component_fa37_or0 = s_CSAwallace_rca24_csa14_csa_component_fa37_xor1 | s_CSAwallace_rca24_csa18_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa20_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa20_and0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa21_and0 = s_CSAwallace_rca24_csa17_csa_component_fa20_or0 & s_CSAwallace_rca24_csa12_csa_component_fa20_and0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa21_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa22_and0 = s_CSAwallace_rca24_csa17_csa_component_fa21_or0 & s_CSAwallace_rca24_csa12_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa22_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa23_and0 = s_CSAwallace_rca24_csa17_csa_component_fa22_or0 & s_CSAwallace_rca24_csa12_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa22_and0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa23_and1 = s_CSAwallace_rca24_csa19_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa22_and0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa23_or0 = s_CSAwallace_rca24_csa19_csa_component_fa23_and0 | s_CSAwallace_rca24_csa19_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa23_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa24_and0 = s_CSAwallace_rca24_csa17_csa_component_fa23_or0 & s_CSAwallace_rca24_csa12_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa24_and1 = s_CSAwallace_rca24_csa19_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa24_or0 = s_CSAwallace_rca24_csa19_csa_component_fa24_and0 | s_CSAwallace_rca24_csa19_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa24_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa25_and0 = s_CSAwallace_rca24_csa17_csa_component_fa24_or0 & s_CSAwallace_rca24_csa12_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa25_and1 = s_CSAwallace_rca24_csa19_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa25_or0 = s_CSAwallace_rca24_csa19_csa_component_fa25_and0 | s_CSAwallace_rca24_csa19_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa25_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa26_and0 = s_CSAwallace_rca24_csa17_csa_component_fa25_or0 & s_CSAwallace_rca24_csa12_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa26_and1 = s_CSAwallace_rca24_csa19_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa26_or0 = s_CSAwallace_rca24_csa19_csa_component_fa26_and0 | s_CSAwallace_rca24_csa19_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa26_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa27_and0 = s_CSAwallace_rca24_csa17_csa_component_fa26_or0 & s_CSAwallace_rca24_csa12_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa27_and1 = s_CSAwallace_rca24_csa19_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa27_or0 = s_CSAwallace_rca24_csa19_csa_component_fa27_and0 | s_CSAwallace_rca24_csa19_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa27_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa28_and0 = s_CSAwallace_rca24_csa17_csa_component_fa27_or0 & s_CSAwallace_rca24_csa12_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa28_and1 = s_CSAwallace_rca24_csa19_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa28_or0 = s_CSAwallace_rca24_csa19_csa_component_fa28_and0 | s_CSAwallace_rca24_csa19_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa28_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa29_and0 = s_CSAwallace_rca24_csa17_csa_component_fa28_or0 & s_CSAwallace_rca24_csa12_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa29_and1 = s_CSAwallace_rca24_csa19_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa29_or0 = s_CSAwallace_rca24_csa19_csa_component_fa29_and0 | s_CSAwallace_rca24_csa19_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa29_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa30_and0 = s_CSAwallace_rca24_csa17_csa_component_fa29_or0 & s_CSAwallace_rca24_csa12_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa30_and1 = s_CSAwallace_rca24_csa19_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa30_or0 = s_CSAwallace_rca24_csa19_csa_component_fa30_and0 | s_CSAwallace_rca24_csa19_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa30_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa31_and0 = s_CSAwallace_rca24_csa17_csa_component_fa30_or0 & s_CSAwallace_rca24_csa12_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa31_and1 = s_CSAwallace_rca24_csa19_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa31_or0 = s_CSAwallace_rca24_csa19_csa_component_fa31_and0 | s_CSAwallace_rca24_csa19_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa31_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa32_and0 = s_CSAwallace_rca24_csa17_csa_component_fa31_or0 & s_CSAwallace_rca24_csa12_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa32_and1 = s_CSAwallace_rca24_csa19_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa32_or0 = s_CSAwallace_rca24_csa19_csa_component_fa32_and0 | s_CSAwallace_rca24_csa19_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa33_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa32_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa33_and0 = s_CSAwallace_rca24_csa17_csa_component_fa32_or0 & s_CSAwallace_rca24_csa12_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa33_and1 = s_CSAwallace_rca24_csa19_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa33_or0 = s_CSAwallace_rca24_csa19_csa_component_fa33_and0 | s_CSAwallace_rca24_csa19_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa34_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa33_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa34_and0 = s_CSAwallace_rca24_csa17_csa_component_fa33_or0 & s_CSAwallace_rca24_csa12_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa34_and1 = s_CSAwallace_rca24_csa19_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa34_or0 = s_CSAwallace_rca24_csa19_csa_component_fa34_and0 | s_CSAwallace_rca24_csa19_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa35_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa34_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa35_and0 = s_CSAwallace_rca24_csa17_csa_component_fa34_or0 & s_CSAwallace_rca24_csa12_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa35_and1 = s_CSAwallace_rca24_csa19_csa_component_fa35_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa35_or0 = s_CSAwallace_rca24_csa19_csa_component_fa35_and0 | s_CSAwallace_rca24_csa19_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa36_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa35_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa36_and0 = s_CSAwallace_rca24_csa17_csa_component_fa35_or0 & s_CSAwallace_rca24_csa12_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa36_and1 = s_CSAwallace_rca24_csa19_csa_component_fa36_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa36_or0 = s_CSAwallace_rca24_csa19_csa_component_fa36_and0 | s_CSAwallace_rca24_csa19_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa37_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa36_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa37_and0 = s_CSAwallace_rca24_csa17_csa_component_fa36_or0 & s_CSAwallace_rca24_csa12_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa37_and1 = s_CSAwallace_rca24_csa19_csa_component_fa37_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa37_or0 = s_CSAwallace_rca24_csa19_csa_component_fa37_and0 | s_CSAwallace_rca24_csa19_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa38_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa37_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa38_and0 = s_CSAwallace_rca24_csa17_csa_component_fa37_or0 & s_CSAwallace_rca24_csa12_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa38_and1 = s_CSAwallace_rca24_csa19_csa_component_fa38_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa38_or0 = s_CSAwallace_rca24_csa19_csa_component_fa38_and0 | s_CSAwallace_rca24_csa19_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa39_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa38_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa39_and0 = s_CSAwallace_rca24_csa17_csa_component_fa38_or0 & s_CSAwallace_rca24_csa12_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa39_and1 = s_CSAwallace_rca24_csa19_csa_component_fa39_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa39_or0 = s_CSAwallace_rca24_csa19_csa_component_fa39_and0 | s_CSAwallace_rca24_csa19_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa40_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa39_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa40_and0 = s_CSAwallace_rca24_csa17_csa_component_fa39_or0 & s_CSAwallace_rca24_csa12_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa40_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa40_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa40_and1 = s_CSAwallace_rca24_csa19_csa_component_fa40_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa40_or0 = s_CSAwallace_rca24_csa19_csa_component_fa40_and0 | s_CSAwallace_rca24_csa19_csa_component_fa40_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa41_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa40_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa41_and0 = s_CSAwallace_rca24_csa17_csa_component_fa40_or0 & s_CSAwallace_rca24_csa12_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa41_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa41_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa41_and1 = s_CSAwallace_rca24_csa19_csa_component_fa41_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa41_or0 = s_CSAwallace_rca24_csa19_csa_component_fa41_and0 | s_CSAwallace_rca24_csa19_csa_component_fa41_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa42_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa41_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa42_and0 = s_CSAwallace_rca24_csa17_csa_component_fa41_or0 & s_CSAwallace_rca24_csa12_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa42_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa42_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa42_and1 = s_CSAwallace_rca24_csa19_csa_component_fa42_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa42_or0 = s_CSAwallace_rca24_csa19_csa_component_fa42_and0 | s_CSAwallace_rca24_csa19_csa_component_fa42_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa43_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa42_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa43_and0 = s_CSAwallace_rca24_csa17_csa_component_fa42_or0 & s_CSAwallace_rca24_csa12_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa43_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa43_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa43_and1 = s_CSAwallace_rca24_csa19_csa_component_fa43_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa43_or0 = s_CSAwallace_rca24_csa19_csa_component_fa43_and0 | s_CSAwallace_rca24_csa19_csa_component_fa43_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa44_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa43_or0 ^ s_CSAwallace_rca24_csa12_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa44_and0 = s_CSAwallace_rca24_csa17_csa_component_fa43_or0 & s_CSAwallace_rca24_csa12_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa44_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa44_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa44_and1 = s_CSAwallace_rca24_csa19_csa_component_fa44_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa44_or0 = s_CSAwallace_rca24_csa19_csa_component_fa44_and0 | s_CSAwallace_rca24_csa19_csa_component_fa44_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa45_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa44_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa45_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa45_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa44_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa45_and1 = s_CSAwallace_rca24_csa19_csa_component_fa45_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa44_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa45_or0 = s_CSAwallace_rca24_csa17_csa_component_fa44_or0 | s_CSAwallace_rca24_csa19_csa_component_fa45_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa46_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa45_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa46_xor1 = s_CSAwallace_rca24_csa19_csa_component_fa46_xor0 ^ s_CSAwallace_rca24_csa7_csa_component_fa45_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa46_and1 = s_CSAwallace_rca24_csa19_csa_component_fa46_xor0 & s_CSAwallace_rca24_csa7_csa_component_fa45_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa46_or0 = s_CSAwallace_rca24_csa17_csa_component_fa45_or0 | s_CSAwallace_rca24_csa19_csa_component_fa46_and1;
  assign s_CSAwallace_rca24_csa19_csa_component_fa47_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa46_or0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa47_xor1 = ~s_CSAwallace_rca24_csa19_csa_component_fa47_xor0;
  assign s_CSAwallace_rca24_csa19_csa_component_fa47_or0 = s_CSAwallace_rca24_csa17_csa_component_fa46_or0 | s_CSAwallace_rca24_csa19_csa_component_fa47_xor0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa6_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa6_xor0 ^ s_CSAwallace_rca24_csa18_csa_component_fa5_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa6_and0 = s_CSAwallace_rca24_csa18_csa_component_fa6_xor0 & s_CSAwallace_rca24_csa18_csa_component_fa5_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa7_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa7_xor0 ^ s_CSAwallace_rca24_csa18_csa_component_fa6_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa7_and0 = s_CSAwallace_rca24_csa18_csa_component_fa7_xor0 & s_CSAwallace_rca24_csa18_csa_component_fa6_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa8_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_csa18_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa8_and0 = s_CSAwallace_rca24_csa18_csa_component_fa8_xor0 & s_CSAwallace_rca24_csa18_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa9_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_csa18_csa_component_fa8_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa9_and0 = s_CSAwallace_rca24_csa18_csa_component_fa9_xor0 & s_CSAwallace_rca24_csa18_csa_component_fa8_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa10_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa10_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa9_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa10_and0 = s_CSAwallace_rca24_csa18_csa_component_fa10_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa9_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa11_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa11_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa11_and0 = s_CSAwallace_rca24_csa18_csa_component_fa11_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa10_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa12_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa12_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa12_and0 = s_CSAwallace_rca24_csa18_csa_component_fa12_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa11_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa13_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa13_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa13_and0 = s_CSAwallace_rca24_csa18_csa_component_fa13_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa12_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa14_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa14_and0 = s_CSAwallace_rca24_csa18_csa_component_fa14_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa13_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa15_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa15_and0 = s_CSAwallace_rca24_csa18_csa_component_fa15_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa14_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa15_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa14_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa15_and1 = s_CSAwallace_rca24_csa20_csa_component_fa15_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa14_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa15_or0 = s_CSAwallace_rca24_csa20_csa_component_fa15_and0 | s_CSAwallace_rca24_csa20_csa_component_fa15_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa16_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa16_and0 = s_CSAwallace_rca24_csa18_csa_component_fa16_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa16_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa15_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa16_and1 = s_CSAwallace_rca24_csa20_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa15_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa16_or0 = s_CSAwallace_rca24_csa20_csa_component_fa16_and0 | s_CSAwallace_rca24_csa20_csa_component_fa16_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa17_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa17_and0 = s_CSAwallace_rca24_csa18_csa_component_fa17_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa17_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa17_and1 = s_CSAwallace_rca24_csa20_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa17_or0 = s_CSAwallace_rca24_csa20_csa_component_fa17_and0 | s_CSAwallace_rca24_csa20_csa_component_fa17_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa18_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa18_and0 = s_CSAwallace_rca24_csa18_csa_component_fa18_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa18_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa18_and1 = s_CSAwallace_rca24_csa20_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa18_or0 = s_CSAwallace_rca24_csa20_csa_component_fa18_and0 | s_CSAwallace_rca24_csa20_csa_component_fa18_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa19_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa19_and0 = s_CSAwallace_rca24_csa18_csa_component_fa19_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa19_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa19_and1 = s_CSAwallace_rca24_csa20_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa19_or0 = s_CSAwallace_rca24_csa20_csa_component_fa19_and0 | s_CSAwallace_rca24_csa20_csa_component_fa19_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa20_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa20_and0 = s_CSAwallace_rca24_csa18_csa_component_fa20_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa20_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa17_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa20_and1 = s_CSAwallace_rca24_csa20_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa17_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa20_or0 = s_CSAwallace_rca24_csa20_csa_component_fa20_and0 | s_CSAwallace_rca24_csa20_csa_component_fa20_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa21_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa21_and0 = s_CSAwallace_rca24_csa18_csa_component_fa21_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa21_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa21_xor0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa21_and1 = s_CSAwallace_rca24_csa20_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa21_xor0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa21_or0 = s_CSAwallace_rca24_csa20_csa_component_fa21_and0 | s_CSAwallace_rca24_csa20_csa_component_fa21_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa22_and0 = s_CSAwallace_rca24_csa18_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa22_xor0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa22_and1 = s_CSAwallace_rca24_csa20_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa22_xor0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa22_or0 = s_CSAwallace_rca24_csa20_csa_component_fa22_and0 | s_CSAwallace_rca24_csa20_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa23_and0 = s_CSAwallace_rca24_csa18_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa23_and1 = s_CSAwallace_rca24_csa20_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa23_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa23_or0 = s_CSAwallace_rca24_csa20_csa_component_fa23_and0 | s_CSAwallace_rca24_csa20_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa24_and0 = s_CSAwallace_rca24_csa18_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa24_and1 = s_CSAwallace_rca24_csa20_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa24_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa24_or0 = s_CSAwallace_rca24_csa20_csa_component_fa24_and0 | s_CSAwallace_rca24_csa20_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa25_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa25_and0 = s_CSAwallace_rca24_csa18_csa_component_fa25_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa25_and1 = s_CSAwallace_rca24_csa20_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa25_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa25_or0 = s_CSAwallace_rca24_csa20_csa_component_fa25_and0 | s_CSAwallace_rca24_csa20_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa26_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa26_and0 = s_CSAwallace_rca24_csa18_csa_component_fa26_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa26_and1 = s_CSAwallace_rca24_csa20_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa26_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa26_or0 = s_CSAwallace_rca24_csa20_csa_component_fa26_and0 | s_CSAwallace_rca24_csa20_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa27_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa27_and0 = s_CSAwallace_rca24_csa18_csa_component_fa27_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa27_and1 = s_CSAwallace_rca24_csa20_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa27_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa27_or0 = s_CSAwallace_rca24_csa20_csa_component_fa27_and0 | s_CSAwallace_rca24_csa20_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa28_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa28_and0 = s_CSAwallace_rca24_csa18_csa_component_fa28_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa28_and1 = s_CSAwallace_rca24_csa20_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa28_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa28_or0 = s_CSAwallace_rca24_csa20_csa_component_fa28_and0 | s_CSAwallace_rca24_csa20_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa29_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa29_and0 = s_CSAwallace_rca24_csa18_csa_component_fa29_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa29_and1 = s_CSAwallace_rca24_csa20_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa29_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa29_or0 = s_CSAwallace_rca24_csa20_csa_component_fa29_and0 | s_CSAwallace_rca24_csa20_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa30_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa30_and0 = s_CSAwallace_rca24_csa18_csa_component_fa30_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa30_and1 = s_CSAwallace_rca24_csa20_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa30_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa30_or0 = s_CSAwallace_rca24_csa20_csa_component_fa30_and0 | s_CSAwallace_rca24_csa20_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa31_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa31_and0 = s_CSAwallace_rca24_csa18_csa_component_fa31_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa31_and1 = s_CSAwallace_rca24_csa20_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa31_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa31_or0 = s_CSAwallace_rca24_csa20_csa_component_fa31_and0 | s_CSAwallace_rca24_csa20_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa32_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa32_and0 = s_CSAwallace_rca24_csa18_csa_component_fa32_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa32_and1 = s_CSAwallace_rca24_csa20_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa32_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa32_or0 = s_CSAwallace_rca24_csa20_csa_component_fa32_and0 | s_CSAwallace_rca24_csa20_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa33_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa33_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa33_and0 = s_CSAwallace_rca24_csa18_csa_component_fa33_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa33_and1 = s_CSAwallace_rca24_csa20_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa33_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa33_or0 = s_CSAwallace_rca24_csa20_csa_component_fa33_and0 | s_CSAwallace_rca24_csa20_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa34_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa34_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa34_and0 = s_CSAwallace_rca24_csa18_csa_component_fa34_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa34_and1 = s_CSAwallace_rca24_csa20_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa34_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa34_or0 = s_CSAwallace_rca24_csa20_csa_component_fa34_and0 | s_CSAwallace_rca24_csa20_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa35_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa35_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa35_and0 = s_CSAwallace_rca24_csa18_csa_component_fa35_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa35_and1 = s_CSAwallace_rca24_csa20_csa_component_fa35_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa35_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa35_or0 = s_CSAwallace_rca24_csa20_csa_component_fa35_and0 | s_CSAwallace_rca24_csa20_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa36_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa36_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa36_and0 = s_CSAwallace_rca24_csa18_csa_component_fa36_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa36_and1 = s_CSAwallace_rca24_csa20_csa_component_fa36_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa36_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa36_or0 = s_CSAwallace_rca24_csa20_csa_component_fa36_and0 | s_CSAwallace_rca24_csa20_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa37_xor0 = s_CSAwallace_rca24_csa18_csa_component_fa37_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa37_and0 = s_CSAwallace_rca24_csa18_csa_component_fa37_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa37_and1 = s_CSAwallace_rca24_csa20_csa_component_fa37_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa37_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa37_or0 = s_CSAwallace_rca24_csa20_csa_component_fa37_and0 | s_CSAwallace_rca24_csa20_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa38_xor0 = s_CSAwallace_rca24_csa17_csa_component_fa38_xor1 ^ s_CSAwallace_rca24_csa18_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa38_and0 = s_CSAwallace_rca24_csa17_csa_component_fa38_xor1 & s_CSAwallace_rca24_csa18_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa20_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa38_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa38_and1 = s_CSAwallace_rca24_csa20_csa_component_fa38_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa38_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa38_or0 = s_CSAwallace_rca24_csa20_csa_component_fa38_and0 | s_CSAwallace_rca24_csa20_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa39_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa39_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa39_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa39_and1 = s_CSAwallace_rca24_csa20_csa_component_fa39_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa39_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa39_or0 = s_CSAwallace_rca24_csa17_csa_component_fa39_xor1 | s_CSAwallace_rca24_csa20_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa40_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa40_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa40_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa40_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa40_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa40_and1 = s_CSAwallace_rca24_csa20_csa_component_fa40_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa40_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa40_or0 = s_CSAwallace_rca24_csa17_csa_component_fa40_xor1 | s_CSAwallace_rca24_csa20_csa_component_fa40_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa41_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa41_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa41_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa41_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa41_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa41_and1 = s_CSAwallace_rca24_csa20_csa_component_fa41_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa41_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa41_or0 = s_CSAwallace_rca24_csa17_csa_component_fa41_xor1 | s_CSAwallace_rca24_csa20_csa_component_fa41_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa42_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa42_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa42_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa42_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa42_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa42_and1 = s_CSAwallace_rca24_csa20_csa_component_fa42_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa42_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa42_or0 = s_CSAwallace_rca24_csa17_csa_component_fa42_xor1 | s_CSAwallace_rca24_csa20_csa_component_fa42_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa43_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa43_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa43_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa43_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa43_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa43_and1 = s_CSAwallace_rca24_csa20_csa_component_fa43_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa43_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa43_or0 = s_CSAwallace_rca24_csa17_csa_component_fa43_xor1 | s_CSAwallace_rca24_csa20_csa_component_fa43_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa44_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa44_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa44_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa44_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa44_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa44_and1 = s_CSAwallace_rca24_csa20_csa_component_fa44_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa44_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa44_or0 = s_CSAwallace_rca24_csa17_csa_component_fa44_xor1 | s_CSAwallace_rca24_csa20_csa_component_fa44_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa45_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa45_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa45_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa45_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa45_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa45_and1 = s_CSAwallace_rca24_csa20_csa_component_fa45_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa45_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa45_or0 = s_CSAwallace_rca24_csa17_csa_component_fa45_xor1 | s_CSAwallace_rca24_csa20_csa_component_fa45_and1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa46_xor0 = ~s_CSAwallace_rca24_csa17_csa_component_fa46_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa46_xor1 = s_CSAwallace_rca24_csa20_csa_component_fa46_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa46_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa46_and1 = s_CSAwallace_rca24_csa20_csa_component_fa46_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa46_xor1;
  assign s_CSAwallace_rca24_csa20_csa_component_fa46_or0 = s_CSAwallace_rca24_csa17_csa_component_fa46_xor1 | s_CSAwallace_rca24_csa20_csa_component_fa46_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa7_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa7_xor0 ^ s_CSAwallace_rca24_csa20_csa_component_fa6_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa7_and0 = s_CSAwallace_rca24_csa20_csa_component_fa7_xor0 & s_CSAwallace_rca24_csa20_csa_component_fa6_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa8_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_csa20_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa8_and0 = s_CSAwallace_rca24_csa20_csa_component_fa8_xor0 & s_CSAwallace_rca24_csa20_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa9_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_csa20_csa_component_fa8_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa9_and0 = s_CSAwallace_rca24_csa20_csa_component_fa9_xor0 & s_CSAwallace_rca24_csa20_csa_component_fa8_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa10_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_csa20_csa_component_fa9_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa10_and0 = s_CSAwallace_rca24_csa20_csa_component_fa10_xor0 & s_CSAwallace_rca24_csa20_csa_component_fa9_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa11_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_csa20_csa_component_fa10_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa11_and0 = s_CSAwallace_rca24_csa20_csa_component_fa11_xor0 & s_CSAwallace_rca24_csa20_csa_component_fa10_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa12_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_csa20_csa_component_fa11_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa12_and0 = s_CSAwallace_rca24_csa20_csa_component_fa12_xor0 & s_CSAwallace_rca24_csa20_csa_component_fa11_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa13_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_csa20_csa_component_fa12_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa13_and0 = s_CSAwallace_rca24_csa20_csa_component_fa13_xor0 & s_CSAwallace_rca24_csa20_csa_component_fa12_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa14_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_csa20_csa_component_fa13_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa14_and0 = s_CSAwallace_rca24_csa20_csa_component_fa14_xor0 & s_CSAwallace_rca24_csa20_csa_component_fa13_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa15_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa15_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa14_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa15_and0 = s_CSAwallace_rca24_csa20_csa_component_fa15_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa14_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa16_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa16_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa16_and0 = s_CSAwallace_rca24_csa20_csa_component_fa16_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa15_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa17_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa17_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa17_and0 = s_CSAwallace_rca24_csa20_csa_component_fa17_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa16_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa18_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa18_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa18_and0 = s_CSAwallace_rca24_csa20_csa_component_fa18_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa17_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa19_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa19_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa19_and0 = s_CSAwallace_rca24_csa20_csa_component_fa19_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa18_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa20_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa20_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa20_and0 = s_CSAwallace_rca24_csa20_csa_component_fa20_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa19_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa21_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa21_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa21_and0 = s_CSAwallace_rca24_csa20_csa_component_fa21_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa20_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa22_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa22_and0 = s_CSAwallace_rca24_csa20_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa21_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa22_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa22_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa21_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa22_and1 = s_CSAwallace_rca24_csa21_csa_component_fa22_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa21_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa22_or0 = s_CSAwallace_rca24_csa21_csa_component_fa22_and0 | s_CSAwallace_rca24_csa21_csa_component_fa22_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa23_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa23_and0 = s_CSAwallace_rca24_csa20_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa23_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa23_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa22_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa23_and1 = s_CSAwallace_rca24_csa21_csa_component_fa23_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa22_and0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa23_or0 = s_CSAwallace_rca24_csa21_csa_component_fa23_and0 | s_CSAwallace_rca24_csa21_csa_component_fa23_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa24_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa24_and0 = s_CSAwallace_rca24_csa20_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa24_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa24_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa24_and1 = s_CSAwallace_rca24_csa21_csa_component_fa24_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa24_or0 = s_CSAwallace_rca24_csa21_csa_component_fa24_and0 | s_CSAwallace_rca24_csa21_csa_component_fa24_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa25_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa25_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa25_and0 = s_CSAwallace_rca24_csa20_csa_component_fa25_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa25_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa25_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa25_and1 = s_CSAwallace_rca24_csa21_csa_component_fa25_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa25_or0 = s_CSAwallace_rca24_csa21_csa_component_fa25_and0 | s_CSAwallace_rca24_csa21_csa_component_fa25_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa26_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa26_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa26_and0 = s_CSAwallace_rca24_csa20_csa_component_fa26_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa26_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa26_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa26_and1 = s_CSAwallace_rca24_csa21_csa_component_fa26_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa26_or0 = s_CSAwallace_rca24_csa21_csa_component_fa26_and0 | s_CSAwallace_rca24_csa21_csa_component_fa26_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa27_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa27_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa27_and0 = s_CSAwallace_rca24_csa20_csa_component_fa27_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa27_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa27_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa27_and1 = s_CSAwallace_rca24_csa21_csa_component_fa27_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa27_or0 = s_CSAwallace_rca24_csa21_csa_component_fa27_and0 | s_CSAwallace_rca24_csa21_csa_component_fa27_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa28_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa28_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa28_and0 = s_CSAwallace_rca24_csa20_csa_component_fa28_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa28_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa28_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa28_and1 = s_CSAwallace_rca24_csa21_csa_component_fa28_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa28_or0 = s_CSAwallace_rca24_csa21_csa_component_fa28_and0 | s_CSAwallace_rca24_csa21_csa_component_fa28_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa29_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa29_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa29_and0 = s_CSAwallace_rca24_csa20_csa_component_fa29_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa29_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa29_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa29_and1 = s_CSAwallace_rca24_csa21_csa_component_fa29_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa29_or0 = s_CSAwallace_rca24_csa21_csa_component_fa29_and0 | s_CSAwallace_rca24_csa21_csa_component_fa29_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa30_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa30_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa30_and0 = s_CSAwallace_rca24_csa20_csa_component_fa30_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa30_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa30_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa30_and1 = s_CSAwallace_rca24_csa21_csa_component_fa30_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa30_or0 = s_CSAwallace_rca24_csa21_csa_component_fa30_and0 | s_CSAwallace_rca24_csa21_csa_component_fa30_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa31_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa31_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa31_and0 = s_CSAwallace_rca24_csa20_csa_component_fa31_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa31_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa31_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa31_and1 = s_CSAwallace_rca24_csa21_csa_component_fa31_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa31_or0 = s_CSAwallace_rca24_csa21_csa_component_fa31_and0 | s_CSAwallace_rca24_csa21_csa_component_fa31_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa32_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa32_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa32_and0 = s_CSAwallace_rca24_csa20_csa_component_fa32_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa32_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa32_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa32_and1 = s_CSAwallace_rca24_csa21_csa_component_fa32_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa32_or0 = s_CSAwallace_rca24_csa21_csa_component_fa32_and0 | s_CSAwallace_rca24_csa21_csa_component_fa32_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa33_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa33_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa33_and0 = s_CSAwallace_rca24_csa20_csa_component_fa33_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa33_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa33_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa33_and1 = s_CSAwallace_rca24_csa21_csa_component_fa33_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa33_or0 = s_CSAwallace_rca24_csa21_csa_component_fa33_and0 | s_CSAwallace_rca24_csa21_csa_component_fa33_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa34_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa34_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa34_and0 = s_CSAwallace_rca24_csa20_csa_component_fa34_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa34_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa34_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa34_and1 = s_CSAwallace_rca24_csa21_csa_component_fa34_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa34_or0 = s_CSAwallace_rca24_csa21_csa_component_fa34_and0 | s_CSAwallace_rca24_csa21_csa_component_fa34_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa35_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa35_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa35_and0 = s_CSAwallace_rca24_csa20_csa_component_fa35_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa35_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa35_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa35_and1 = s_CSAwallace_rca24_csa21_csa_component_fa35_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa35_or0 = s_CSAwallace_rca24_csa21_csa_component_fa35_and0 | s_CSAwallace_rca24_csa21_csa_component_fa35_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa36_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa36_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa36_and0 = s_CSAwallace_rca24_csa20_csa_component_fa36_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa36_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa36_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa36_and1 = s_CSAwallace_rca24_csa21_csa_component_fa36_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa36_or0 = s_CSAwallace_rca24_csa21_csa_component_fa36_and0 | s_CSAwallace_rca24_csa21_csa_component_fa36_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa37_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa37_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa37_and0 = s_CSAwallace_rca24_csa20_csa_component_fa37_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa37_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa37_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa37_and1 = s_CSAwallace_rca24_csa21_csa_component_fa37_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa37_or0 = s_CSAwallace_rca24_csa21_csa_component_fa37_and0 | s_CSAwallace_rca24_csa21_csa_component_fa37_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa38_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa38_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa38_and0 = s_CSAwallace_rca24_csa20_csa_component_fa38_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa38_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa38_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa38_and1 = s_CSAwallace_rca24_csa21_csa_component_fa38_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa38_or0 = s_CSAwallace_rca24_csa21_csa_component_fa38_and0 | s_CSAwallace_rca24_csa21_csa_component_fa38_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa39_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa39_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa39_and0 = s_CSAwallace_rca24_csa20_csa_component_fa39_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa39_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa39_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa39_and1 = s_CSAwallace_rca24_csa21_csa_component_fa39_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa39_or0 = s_CSAwallace_rca24_csa21_csa_component_fa39_and0 | s_CSAwallace_rca24_csa21_csa_component_fa39_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa40_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa40_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa40_and0 = s_CSAwallace_rca24_csa20_csa_component_fa40_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa40_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa40_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa40_and1 = s_CSAwallace_rca24_csa21_csa_component_fa40_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa40_or0 = s_CSAwallace_rca24_csa21_csa_component_fa40_and0 | s_CSAwallace_rca24_csa21_csa_component_fa40_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa41_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa41_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa41_and0 = s_CSAwallace_rca24_csa20_csa_component_fa41_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa41_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa41_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa41_and1 = s_CSAwallace_rca24_csa21_csa_component_fa41_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa41_or0 = s_CSAwallace_rca24_csa21_csa_component_fa41_and0 | s_CSAwallace_rca24_csa21_csa_component_fa41_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa42_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa42_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa42_and0 = s_CSAwallace_rca24_csa20_csa_component_fa42_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa42_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa42_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa42_and1 = s_CSAwallace_rca24_csa21_csa_component_fa42_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa42_or0 = s_CSAwallace_rca24_csa21_csa_component_fa42_and0 | s_CSAwallace_rca24_csa21_csa_component_fa42_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa43_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa43_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa43_and0 = s_CSAwallace_rca24_csa20_csa_component_fa43_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa43_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa43_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa43_and1 = s_CSAwallace_rca24_csa21_csa_component_fa43_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa43_or0 = s_CSAwallace_rca24_csa21_csa_component_fa43_and0 | s_CSAwallace_rca24_csa21_csa_component_fa43_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa44_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa44_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa44_and0 = s_CSAwallace_rca24_csa20_csa_component_fa44_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa44_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa44_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa44_and1 = s_CSAwallace_rca24_csa21_csa_component_fa44_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa44_or0 = s_CSAwallace_rca24_csa21_csa_component_fa44_and0 | s_CSAwallace_rca24_csa21_csa_component_fa44_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa45_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa45_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa44_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa45_and0 = s_CSAwallace_rca24_csa20_csa_component_fa45_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa44_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa45_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa45_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa44_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa45_and1 = s_CSAwallace_rca24_csa21_csa_component_fa45_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa44_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa45_or0 = s_CSAwallace_rca24_csa21_csa_component_fa45_and0 | s_CSAwallace_rca24_csa21_csa_component_fa45_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa46_xor0 = s_CSAwallace_rca24_csa20_csa_component_fa46_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa45_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa46_and0 = s_CSAwallace_rca24_csa20_csa_component_fa46_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa45_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa46_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa46_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa45_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa46_and1 = s_CSAwallace_rca24_csa21_csa_component_fa46_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa45_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa46_or0 = s_CSAwallace_rca24_csa21_csa_component_fa46_and0 | s_CSAwallace_rca24_csa21_csa_component_fa46_and1;
  assign s_CSAwallace_rca24_csa21_csa_component_fa47_xor0 = s_CSAwallace_rca24_csa19_csa_component_fa47_xor1 ^ s_CSAwallace_rca24_csa20_csa_component_fa46_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa47_and0 = s_CSAwallace_rca24_csa19_csa_component_fa47_xor1 & s_CSAwallace_rca24_csa20_csa_component_fa46_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa47_xor1 = s_CSAwallace_rca24_csa21_csa_component_fa47_xor0 ^ s_CSAwallace_rca24_csa19_csa_component_fa46_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa47_and1 = s_CSAwallace_rca24_csa21_csa_component_fa47_xor0 & s_CSAwallace_rca24_csa19_csa_component_fa46_or0;
  assign s_CSAwallace_rca24_csa21_csa_component_fa47_or0 = s_CSAwallace_rca24_csa21_csa_component_fa47_and0 | s_CSAwallace_rca24_csa21_csa_component_fa47_and1;
  assign s_CSAwallace_rca24_u_rca48_fa8_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa8_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_u_rca48_fa8_and0 = s_CSAwallace_rca24_csa21_csa_component_fa8_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa7_and0;
  assign s_CSAwallace_rca24_u_rca48_fa9_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa9_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa8_and0;
  assign s_CSAwallace_rca24_u_rca48_fa9_and0 = s_CSAwallace_rca24_csa21_csa_component_fa9_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa8_and0;
  assign s_CSAwallace_rca24_u_rca48_fa9_xor1 = s_CSAwallace_rca24_u_rca48_fa9_xor0 ^ s_CSAwallace_rca24_u_rca48_fa8_and0;
  assign s_CSAwallace_rca24_u_rca48_fa9_and1 = s_CSAwallace_rca24_u_rca48_fa9_xor0 & s_CSAwallace_rca24_u_rca48_fa8_and0;
  assign s_CSAwallace_rca24_u_rca48_fa9_or0 = s_CSAwallace_rca24_u_rca48_fa9_and0 | s_CSAwallace_rca24_u_rca48_fa9_and1;
  assign s_CSAwallace_rca24_u_rca48_fa10_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa10_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa9_and0;
  assign s_CSAwallace_rca24_u_rca48_fa10_and0 = s_CSAwallace_rca24_csa21_csa_component_fa10_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa9_and0;
  assign s_CSAwallace_rca24_u_rca48_fa10_xor1 = s_CSAwallace_rca24_u_rca48_fa10_xor0 ^ s_CSAwallace_rca24_u_rca48_fa9_or0;
  assign s_CSAwallace_rca24_u_rca48_fa10_and1 = s_CSAwallace_rca24_u_rca48_fa10_xor0 & s_CSAwallace_rca24_u_rca48_fa9_or0;
  assign s_CSAwallace_rca24_u_rca48_fa10_or0 = s_CSAwallace_rca24_u_rca48_fa10_and0 | s_CSAwallace_rca24_u_rca48_fa10_and1;
  assign s_CSAwallace_rca24_u_rca48_fa11_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa11_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa10_and0;
  assign s_CSAwallace_rca24_u_rca48_fa11_and0 = s_CSAwallace_rca24_csa21_csa_component_fa11_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa10_and0;
  assign s_CSAwallace_rca24_u_rca48_fa11_xor1 = s_CSAwallace_rca24_u_rca48_fa11_xor0 ^ s_CSAwallace_rca24_u_rca48_fa10_or0;
  assign s_CSAwallace_rca24_u_rca48_fa11_and1 = s_CSAwallace_rca24_u_rca48_fa11_xor0 & s_CSAwallace_rca24_u_rca48_fa10_or0;
  assign s_CSAwallace_rca24_u_rca48_fa11_or0 = s_CSAwallace_rca24_u_rca48_fa11_and0 | s_CSAwallace_rca24_u_rca48_fa11_and1;
  assign s_CSAwallace_rca24_u_rca48_fa12_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa12_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa11_and0;
  assign s_CSAwallace_rca24_u_rca48_fa12_and0 = s_CSAwallace_rca24_csa21_csa_component_fa12_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa11_and0;
  assign s_CSAwallace_rca24_u_rca48_fa12_xor1 = s_CSAwallace_rca24_u_rca48_fa12_xor0 ^ s_CSAwallace_rca24_u_rca48_fa11_or0;
  assign s_CSAwallace_rca24_u_rca48_fa12_and1 = s_CSAwallace_rca24_u_rca48_fa12_xor0 & s_CSAwallace_rca24_u_rca48_fa11_or0;
  assign s_CSAwallace_rca24_u_rca48_fa12_or0 = s_CSAwallace_rca24_u_rca48_fa12_and0 | s_CSAwallace_rca24_u_rca48_fa12_and1;
  assign s_CSAwallace_rca24_u_rca48_fa13_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa13_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa12_and0;
  assign s_CSAwallace_rca24_u_rca48_fa13_and0 = s_CSAwallace_rca24_csa21_csa_component_fa13_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa12_and0;
  assign s_CSAwallace_rca24_u_rca48_fa13_xor1 = s_CSAwallace_rca24_u_rca48_fa13_xor0 ^ s_CSAwallace_rca24_u_rca48_fa12_or0;
  assign s_CSAwallace_rca24_u_rca48_fa13_and1 = s_CSAwallace_rca24_u_rca48_fa13_xor0 & s_CSAwallace_rca24_u_rca48_fa12_or0;
  assign s_CSAwallace_rca24_u_rca48_fa13_or0 = s_CSAwallace_rca24_u_rca48_fa13_and0 | s_CSAwallace_rca24_u_rca48_fa13_and1;
  assign s_CSAwallace_rca24_u_rca48_fa14_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa14_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa13_and0;
  assign s_CSAwallace_rca24_u_rca48_fa14_and0 = s_CSAwallace_rca24_csa21_csa_component_fa14_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa13_and0;
  assign s_CSAwallace_rca24_u_rca48_fa14_xor1 = s_CSAwallace_rca24_u_rca48_fa14_xor0 ^ s_CSAwallace_rca24_u_rca48_fa13_or0;
  assign s_CSAwallace_rca24_u_rca48_fa14_and1 = s_CSAwallace_rca24_u_rca48_fa14_xor0 & s_CSAwallace_rca24_u_rca48_fa13_or0;
  assign s_CSAwallace_rca24_u_rca48_fa14_or0 = s_CSAwallace_rca24_u_rca48_fa14_and0 | s_CSAwallace_rca24_u_rca48_fa14_and1;
  assign s_CSAwallace_rca24_u_rca48_fa15_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa15_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa14_and0;
  assign s_CSAwallace_rca24_u_rca48_fa15_and0 = s_CSAwallace_rca24_csa21_csa_component_fa15_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa14_and0;
  assign s_CSAwallace_rca24_u_rca48_fa15_xor1 = s_CSAwallace_rca24_u_rca48_fa15_xor0 ^ s_CSAwallace_rca24_u_rca48_fa14_or0;
  assign s_CSAwallace_rca24_u_rca48_fa15_and1 = s_CSAwallace_rca24_u_rca48_fa15_xor0 & s_CSAwallace_rca24_u_rca48_fa14_or0;
  assign s_CSAwallace_rca24_u_rca48_fa15_or0 = s_CSAwallace_rca24_u_rca48_fa15_and0 | s_CSAwallace_rca24_u_rca48_fa15_and1;
  assign s_CSAwallace_rca24_u_rca48_fa16_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa16_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa15_and0;
  assign s_CSAwallace_rca24_u_rca48_fa16_and0 = s_CSAwallace_rca24_csa21_csa_component_fa16_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa15_and0;
  assign s_CSAwallace_rca24_u_rca48_fa16_xor1 = s_CSAwallace_rca24_u_rca48_fa16_xor0 ^ s_CSAwallace_rca24_u_rca48_fa15_or0;
  assign s_CSAwallace_rca24_u_rca48_fa16_and1 = s_CSAwallace_rca24_u_rca48_fa16_xor0 & s_CSAwallace_rca24_u_rca48_fa15_or0;
  assign s_CSAwallace_rca24_u_rca48_fa16_or0 = s_CSAwallace_rca24_u_rca48_fa16_and0 | s_CSAwallace_rca24_u_rca48_fa16_and1;
  assign s_CSAwallace_rca24_u_rca48_fa17_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa17_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_u_rca48_fa17_and0 = s_CSAwallace_rca24_csa21_csa_component_fa17_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa16_and0;
  assign s_CSAwallace_rca24_u_rca48_fa17_xor1 = s_CSAwallace_rca24_u_rca48_fa17_xor0 ^ s_CSAwallace_rca24_u_rca48_fa16_or0;
  assign s_CSAwallace_rca24_u_rca48_fa17_and1 = s_CSAwallace_rca24_u_rca48_fa17_xor0 & s_CSAwallace_rca24_u_rca48_fa16_or0;
  assign s_CSAwallace_rca24_u_rca48_fa17_or0 = s_CSAwallace_rca24_u_rca48_fa17_and0 | s_CSAwallace_rca24_u_rca48_fa17_and1;
  assign s_CSAwallace_rca24_u_rca48_fa18_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa18_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa17_and0;
  assign s_CSAwallace_rca24_u_rca48_fa18_and0 = s_CSAwallace_rca24_csa21_csa_component_fa18_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa17_and0;
  assign s_CSAwallace_rca24_u_rca48_fa18_xor1 = s_CSAwallace_rca24_u_rca48_fa18_xor0 ^ s_CSAwallace_rca24_u_rca48_fa17_or0;
  assign s_CSAwallace_rca24_u_rca48_fa18_and1 = s_CSAwallace_rca24_u_rca48_fa18_xor0 & s_CSAwallace_rca24_u_rca48_fa17_or0;
  assign s_CSAwallace_rca24_u_rca48_fa18_or0 = s_CSAwallace_rca24_u_rca48_fa18_and0 | s_CSAwallace_rca24_u_rca48_fa18_and1;
  assign s_CSAwallace_rca24_u_rca48_fa19_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa19_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa18_and0;
  assign s_CSAwallace_rca24_u_rca48_fa19_and0 = s_CSAwallace_rca24_csa21_csa_component_fa19_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa18_and0;
  assign s_CSAwallace_rca24_u_rca48_fa19_xor1 = s_CSAwallace_rca24_u_rca48_fa19_xor0 ^ s_CSAwallace_rca24_u_rca48_fa18_or0;
  assign s_CSAwallace_rca24_u_rca48_fa19_and1 = s_CSAwallace_rca24_u_rca48_fa19_xor0 & s_CSAwallace_rca24_u_rca48_fa18_or0;
  assign s_CSAwallace_rca24_u_rca48_fa19_or0 = s_CSAwallace_rca24_u_rca48_fa19_and0 | s_CSAwallace_rca24_u_rca48_fa19_and1;
  assign s_CSAwallace_rca24_u_rca48_fa20_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa20_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa19_and0;
  assign s_CSAwallace_rca24_u_rca48_fa20_and0 = s_CSAwallace_rca24_csa21_csa_component_fa20_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa19_and0;
  assign s_CSAwallace_rca24_u_rca48_fa20_xor1 = s_CSAwallace_rca24_u_rca48_fa20_xor0 ^ s_CSAwallace_rca24_u_rca48_fa19_or0;
  assign s_CSAwallace_rca24_u_rca48_fa20_and1 = s_CSAwallace_rca24_u_rca48_fa20_xor0 & s_CSAwallace_rca24_u_rca48_fa19_or0;
  assign s_CSAwallace_rca24_u_rca48_fa20_or0 = s_CSAwallace_rca24_u_rca48_fa20_and0 | s_CSAwallace_rca24_u_rca48_fa20_and1;
  assign s_CSAwallace_rca24_u_rca48_fa21_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa21_xor0 ^ s_CSAwallace_rca24_csa21_csa_component_fa20_and0;
  assign s_CSAwallace_rca24_u_rca48_fa21_and0 = s_CSAwallace_rca24_csa21_csa_component_fa21_xor0 & s_CSAwallace_rca24_csa21_csa_component_fa20_and0;
  assign s_CSAwallace_rca24_u_rca48_fa21_xor1 = s_CSAwallace_rca24_u_rca48_fa21_xor0 ^ s_CSAwallace_rca24_u_rca48_fa20_or0;
  assign s_CSAwallace_rca24_u_rca48_fa21_and1 = s_CSAwallace_rca24_u_rca48_fa21_xor0 & s_CSAwallace_rca24_u_rca48_fa20_or0;
  assign s_CSAwallace_rca24_u_rca48_fa21_or0 = s_CSAwallace_rca24_u_rca48_fa21_and0 | s_CSAwallace_rca24_u_rca48_fa21_and1;
  assign s_CSAwallace_rca24_u_rca48_fa22_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa22_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa21_and0;
  assign s_CSAwallace_rca24_u_rca48_fa22_and0 = s_CSAwallace_rca24_csa21_csa_component_fa22_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa21_and0;
  assign s_CSAwallace_rca24_u_rca48_fa22_xor1 = s_CSAwallace_rca24_u_rca48_fa22_xor0 ^ s_CSAwallace_rca24_u_rca48_fa21_or0;
  assign s_CSAwallace_rca24_u_rca48_fa22_and1 = s_CSAwallace_rca24_u_rca48_fa22_xor0 & s_CSAwallace_rca24_u_rca48_fa21_or0;
  assign s_CSAwallace_rca24_u_rca48_fa22_or0 = s_CSAwallace_rca24_u_rca48_fa22_and0 | s_CSAwallace_rca24_u_rca48_fa22_and1;
  assign s_CSAwallace_rca24_u_rca48_fa23_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa23_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_u_rca48_fa23_and0 = s_CSAwallace_rca24_csa21_csa_component_fa23_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa22_or0;
  assign s_CSAwallace_rca24_u_rca48_fa23_xor1 = s_CSAwallace_rca24_u_rca48_fa23_xor0 ^ s_CSAwallace_rca24_u_rca48_fa22_or0;
  assign s_CSAwallace_rca24_u_rca48_fa23_and1 = s_CSAwallace_rca24_u_rca48_fa23_xor0 & s_CSAwallace_rca24_u_rca48_fa22_or0;
  assign s_CSAwallace_rca24_u_rca48_fa23_or0 = s_CSAwallace_rca24_u_rca48_fa23_and0 | s_CSAwallace_rca24_u_rca48_fa23_and1;
  assign s_CSAwallace_rca24_u_rca48_fa24_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa24_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_u_rca48_fa24_and0 = s_CSAwallace_rca24_csa21_csa_component_fa24_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa23_or0;
  assign s_CSAwallace_rca24_u_rca48_fa24_xor1 = s_CSAwallace_rca24_u_rca48_fa24_xor0 ^ s_CSAwallace_rca24_u_rca48_fa23_or0;
  assign s_CSAwallace_rca24_u_rca48_fa24_and1 = s_CSAwallace_rca24_u_rca48_fa24_xor0 & s_CSAwallace_rca24_u_rca48_fa23_or0;
  assign s_CSAwallace_rca24_u_rca48_fa24_or0 = s_CSAwallace_rca24_u_rca48_fa24_and0 | s_CSAwallace_rca24_u_rca48_fa24_and1;
  assign s_CSAwallace_rca24_u_rca48_fa25_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa25_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_u_rca48_fa25_and0 = s_CSAwallace_rca24_csa21_csa_component_fa25_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa24_or0;
  assign s_CSAwallace_rca24_u_rca48_fa25_xor1 = s_CSAwallace_rca24_u_rca48_fa25_xor0 ^ s_CSAwallace_rca24_u_rca48_fa24_or0;
  assign s_CSAwallace_rca24_u_rca48_fa25_and1 = s_CSAwallace_rca24_u_rca48_fa25_xor0 & s_CSAwallace_rca24_u_rca48_fa24_or0;
  assign s_CSAwallace_rca24_u_rca48_fa25_or0 = s_CSAwallace_rca24_u_rca48_fa25_and0 | s_CSAwallace_rca24_u_rca48_fa25_and1;
  assign s_CSAwallace_rca24_u_rca48_fa26_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa26_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_u_rca48_fa26_and0 = s_CSAwallace_rca24_csa21_csa_component_fa26_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa25_or0;
  assign s_CSAwallace_rca24_u_rca48_fa26_xor1 = s_CSAwallace_rca24_u_rca48_fa26_xor0 ^ s_CSAwallace_rca24_u_rca48_fa25_or0;
  assign s_CSAwallace_rca24_u_rca48_fa26_and1 = s_CSAwallace_rca24_u_rca48_fa26_xor0 & s_CSAwallace_rca24_u_rca48_fa25_or0;
  assign s_CSAwallace_rca24_u_rca48_fa26_or0 = s_CSAwallace_rca24_u_rca48_fa26_and0 | s_CSAwallace_rca24_u_rca48_fa26_and1;
  assign s_CSAwallace_rca24_u_rca48_fa27_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa27_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_u_rca48_fa27_and0 = s_CSAwallace_rca24_csa21_csa_component_fa27_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa26_or0;
  assign s_CSAwallace_rca24_u_rca48_fa27_xor1 = s_CSAwallace_rca24_u_rca48_fa27_xor0 ^ s_CSAwallace_rca24_u_rca48_fa26_or0;
  assign s_CSAwallace_rca24_u_rca48_fa27_and1 = s_CSAwallace_rca24_u_rca48_fa27_xor0 & s_CSAwallace_rca24_u_rca48_fa26_or0;
  assign s_CSAwallace_rca24_u_rca48_fa27_or0 = s_CSAwallace_rca24_u_rca48_fa27_and0 | s_CSAwallace_rca24_u_rca48_fa27_and1;
  assign s_CSAwallace_rca24_u_rca48_fa28_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa28_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_u_rca48_fa28_and0 = s_CSAwallace_rca24_csa21_csa_component_fa28_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa27_or0;
  assign s_CSAwallace_rca24_u_rca48_fa28_xor1 = s_CSAwallace_rca24_u_rca48_fa28_xor0 ^ s_CSAwallace_rca24_u_rca48_fa27_or0;
  assign s_CSAwallace_rca24_u_rca48_fa28_and1 = s_CSAwallace_rca24_u_rca48_fa28_xor0 & s_CSAwallace_rca24_u_rca48_fa27_or0;
  assign s_CSAwallace_rca24_u_rca48_fa28_or0 = s_CSAwallace_rca24_u_rca48_fa28_and0 | s_CSAwallace_rca24_u_rca48_fa28_and1;
  assign s_CSAwallace_rca24_u_rca48_fa29_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa29_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_u_rca48_fa29_and0 = s_CSAwallace_rca24_csa21_csa_component_fa29_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa28_or0;
  assign s_CSAwallace_rca24_u_rca48_fa29_xor1 = s_CSAwallace_rca24_u_rca48_fa29_xor0 ^ s_CSAwallace_rca24_u_rca48_fa28_or0;
  assign s_CSAwallace_rca24_u_rca48_fa29_and1 = s_CSAwallace_rca24_u_rca48_fa29_xor0 & s_CSAwallace_rca24_u_rca48_fa28_or0;
  assign s_CSAwallace_rca24_u_rca48_fa29_or0 = s_CSAwallace_rca24_u_rca48_fa29_and0 | s_CSAwallace_rca24_u_rca48_fa29_and1;
  assign s_CSAwallace_rca24_u_rca48_fa30_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa30_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_u_rca48_fa30_and0 = s_CSAwallace_rca24_csa21_csa_component_fa30_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa29_or0;
  assign s_CSAwallace_rca24_u_rca48_fa30_xor1 = s_CSAwallace_rca24_u_rca48_fa30_xor0 ^ s_CSAwallace_rca24_u_rca48_fa29_or0;
  assign s_CSAwallace_rca24_u_rca48_fa30_and1 = s_CSAwallace_rca24_u_rca48_fa30_xor0 & s_CSAwallace_rca24_u_rca48_fa29_or0;
  assign s_CSAwallace_rca24_u_rca48_fa30_or0 = s_CSAwallace_rca24_u_rca48_fa30_and0 | s_CSAwallace_rca24_u_rca48_fa30_and1;
  assign s_CSAwallace_rca24_u_rca48_fa31_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa31_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_u_rca48_fa31_and0 = s_CSAwallace_rca24_csa21_csa_component_fa31_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa30_or0;
  assign s_CSAwallace_rca24_u_rca48_fa31_xor1 = s_CSAwallace_rca24_u_rca48_fa31_xor0 ^ s_CSAwallace_rca24_u_rca48_fa30_or0;
  assign s_CSAwallace_rca24_u_rca48_fa31_and1 = s_CSAwallace_rca24_u_rca48_fa31_xor0 & s_CSAwallace_rca24_u_rca48_fa30_or0;
  assign s_CSAwallace_rca24_u_rca48_fa31_or0 = s_CSAwallace_rca24_u_rca48_fa31_and0 | s_CSAwallace_rca24_u_rca48_fa31_and1;
  assign s_CSAwallace_rca24_u_rca48_fa32_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa32_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_u_rca48_fa32_and0 = s_CSAwallace_rca24_csa21_csa_component_fa32_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa31_or0;
  assign s_CSAwallace_rca24_u_rca48_fa32_xor1 = s_CSAwallace_rca24_u_rca48_fa32_xor0 ^ s_CSAwallace_rca24_u_rca48_fa31_or0;
  assign s_CSAwallace_rca24_u_rca48_fa32_and1 = s_CSAwallace_rca24_u_rca48_fa32_xor0 & s_CSAwallace_rca24_u_rca48_fa31_or0;
  assign s_CSAwallace_rca24_u_rca48_fa32_or0 = s_CSAwallace_rca24_u_rca48_fa32_and0 | s_CSAwallace_rca24_u_rca48_fa32_and1;
  assign s_CSAwallace_rca24_u_rca48_fa33_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa33_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_u_rca48_fa33_and0 = s_CSAwallace_rca24_csa21_csa_component_fa33_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa32_or0;
  assign s_CSAwallace_rca24_u_rca48_fa33_xor1 = s_CSAwallace_rca24_u_rca48_fa33_xor0 ^ s_CSAwallace_rca24_u_rca48_fa32_or0;
  assign s_CSAwallace_rca24_u_rca48_fa33_and1 = s_CSAwallace_rca24_u_rca48_fa33_xor0 & s_CSAwallace_rca24_u_rca48_fa32_or0;
  assign s_CSAwallace_rca24_u_rca48_fa33_or0 = s_CSAwallace_rca24_u_rca48_fa33_and0 | s_CSAwallace_rca24_u_rca48_fa33_and1;
  assign s_CSAwallace_rca24_u_rca48_fa34_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa34_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_u_rca48_fa34_and0 = s_CSAwallace_rca24_csa21_csa_component_fa34_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa33_or0;
  assign s_CSAwallace_rca24_u_rca48_fa34_xor1 = s_CSAwallace_rca24_u_rca48_fa34_xor0 ^ s_CSAwallace_rca24_u_rca48_fa33_or0;
  assign s_CSAwallace_rca24_u_rca48_fa34_and1 = s_CSAwallace_rca24_u_rca48_fa34_xor0 & s_CSAwallace_rca24_u_rca48_fa33_or0;
  assign s_CSAwallace_rca24_u_rca48_fa34_or0 = s_CSAwallace_rca24_u_rca48_fa34_and0 | s_CSAwallace_rca24_u_rca48_fa34_and1;
  assign s_CSAwallace_rca24_u_rca48_fa35_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa35_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_u_rca48_fa35_and0 = s_CSAwallace_rca24_csa21_csa_component_fa35_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa34_or0;
  assign s_CSAwallace_rca24_u_rca48_fa35_xor1 = s_CSAwallace_rca24_u_rca48_fa35_xor0 ^ s_CSAwallace_rca24_u_rca48_fa34_or0;
  assign s_CSAwallace_rca24_u_rca48_fa35_and1 = s_CSAwallace_rca24_u_rca48_fa35_xor0 & s_CSAwallace_rca24_u_rca48_fa34_or0;
  assign s_CSAwallace_rca24_u_rca48_fa35_or0 = s_CSAwallace_rca24_u_rca48_fa35_and0 | s_CSAwallace_rca24_u_rca48_fa35_and1;
  assign s_CSAwallace_rca24_u_rca48_fa36_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa36_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_u_rca48_fa36_and0 = s_CSAwallace_rca24_csa21_csa_component_fa36_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa35_or0;
  assign s_CSAwallace_rca24_u_rca48_fa36_xor1 = s_CSAwallace_rca24_u_rca48_fa36_xor0 ^ s_CSAwallace_rca24_u_rca48_fa35_or0;
  assign s_CSAwallace_rca24_u_rca48_fa36_and1 = s_CSAwallace_rca24_u_rca48_fa36_xor0 & s_CSAwallace_rca24_u_rca48_fa35_or0;
  assign s_CSAwallace_rca24_u_rca48_fa36_or0 = s_CSAwallace_rca24_u_rca48_fa36_and0 | s_CSAwallace_rca24_u_rca48_fa36_and1;
  assign s_CSAwallace_rca24_u_rca48_fa37_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa37_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_u_rca48_fa37_and0 = s_CSAwallace_rca24_csa21_csa_component_fa37_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa36_or0;
  assign s_CSAwallace_rca24_u_rca48_fa37_xor1 = s_CSAwallace_rca24_u_rca48_fa37_xor0 ^ s_CSAwallace_rca24_u_rca48_fa36_or0;
  assign s_CSAwallace_rca24_u_rca48_fa37_and1 = s_CSAwallace_rca24_u_rca48_fa37_xor0 & s_CSAwallace_rca24_u_rca48_fa36_or0;
  assign s_CSAwallace_rca24_u_rca48_fa37_or0 = s_CSAwallace_rca24_u_rca48_fa37_and0 | s_CSAwallace_rca24_u_rca48_fa37_and1;
  assign s_CSAwallace_rca24_u_rca48_fa38_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa38_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_u_rca48_fa38_and0 = s_CSAwallace_rca24_csa21_csa_component_fa38_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa37_or0;
  assign s_CSAwallace_rca24_u_rca48_fa38_xor1 = s_CSAwallace_rca24_u_rca48_fa38_xor0 ^ s_CSAwallace_rca24_u_rca48_fa37_or0;
  assign s_CSAwallace_rca24_u_rca48_fa38_and1 = s_CSAwallace_rca24_u_rca48_fa38_xor0 & s_CSAwallace_rca24_u_rca48_fa37_or0;
  assign s_CSAwallace_rca24_u_rca48_fa38_or0 = s_CSAwallace_rca24_u_rca48_fa38_and0 | s_CSAwallace_rca24_u_rca48_fa38_and1;
  assign s_CSAwallace_rca24_u_rca48_fa39_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa39_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_u_rca48_fa39_and0 = s_CSAwallace_rca24_csa21_csa_component_fa39_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa38_or0;
  assign s_CSAwallace_rca24_u_rca48_fa39_xor1 = s_CSAwallace_rca24_u_rca48_fa39_xor0 ^ s_CSAwallace_rca24_u_rca48_fa38_or0;
  assign s_CSAwallace_rca24_u_rca48_fa39_and1 = s_CSAwallace_rca24_u_rca48_fa39_xor0 & s_CSAwallace_rca24_u_rca48_fa38_or0;
  assign s_CSAwallace_rca24_u_rca48_fa39_or0 = s_CSAwallace_rca24_u_rca48_fa39_and0 | s_CSAwallace_rca24_u_rca48_fa39_and1;
  assign s_CSAwallace_rca24_u_rca48_fa40_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa40_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_u_rca48_fa40_and0 = s_CSAwallace_rca24_csa21_csa_component_fa40_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa39_or0;
  assign s_CSAwallace_rca24_u_rca48_fa40_xor1 = s_CSAwallace_rca24_u_rca48_fa40_xor0 ^ s_CSAwallace_rca24_u_rca48_fa39_or0;
  assign s_CSAwallace_rca24_u_rca48_fa40_and1 = s_CSAwallace_rca24_u_rca48_fa40_xor0 & s_CSAwallace_rca24_u_rca48_fa39_or0;
  assign s_CSAwallace_rca24_u_rca48_fa40_or0 = s_CSAwallace_rca24_u_rca48_fa40_and0 | s_CSAwallace_rca24_u_rca48_fa40_and1;
  assign s_CSAwallace_rca24_u_rca48_fa41_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa41_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_u_rca48_fa41_and0 = s_CSAwallace_rca24_csa21_csa_component_fa41_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa40_or0;
  assign s_CSAwallace_rca24_u_rca48_fa41_xor1 = s_CSAwallace_rca24_u_rca48_fa41_xor0 ^ s_CSAwallace_rca24_u_rca48_fa40_or0;
  assign s_CSAwallace_rca24_u_rca48_fa41_and1 = s_CSAwallace_rca24_u_rca48_fa41_xor0 & s_CSAwallace_rca24_u_rca48_fa40_or0;
  assign s_CSAwallace_rca24_u_rca48_fa41_or0 = s_CSAwallace_rca24_u_rca48_fa41_and0 | s_CSAwallace_rca24_u_rca48_fa41_and1;
  assign s_CSAwallace_rca24_u_rca48_fa42_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa42_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_u_rca48_fa42_and0 = s_CSAwallace_rca24_csa21_csa_component_fa42_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa41_or0;
  assign s_CSAwallace_rca24_u_rca48_fa42_xor1 = s_CSAwallace_rca24_u_rca48_fa42_xor0 ^ s_CSAwallace_rca24_u_rca48_fa41_or0;
  assign s_CSAwallace_rca24_u_rca48_fa42_and1 = s_CSAwallace_rca24_u_rca48_fa42_xor0 & s_CSAwallace_rca24_u_rca48_fa41_or0;
  assign s_CSAwallace_rca24_u_rca48_fa42_or0 = s_CSAwallace_rca24_u_rca48_fa42_and0 | s_CSAwallace_rca24_u_rca48_fa42_and1;
  assign s_CSAwallace_rca24_u_rca48_fa43_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa43_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_u_rca48_fa43_and0 = s_CSAwallace_rca24_csa21_csa_component_fa43_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa42_or0;
  assign s_CSAwallace_rca24_u_rca48_fa43_xor1 = s_CSAwallace_rca24_u_rca48_fa43_xor0 ^ s_CSAwallace_rca24_u_rca48_fa42_or0;
  assign s_CSAwallace_rca24_u_rca48_fa43_and1 = s_CSAwallace_rca24_u_rca48_fa43_xor0 & s_CSAwallace_rca24_u_rca48_fa42_or0;
  assign s_CSAwallace_rca24_u_rca48_fa43_or0 = s_CSAwallace_rca24_u_rca48_fa43_and0 | s_CSAwallace_rca24_u_rca48_fa43_and1;
  assign s_CSAwallace_rca24_u_rca48_fa44_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa44_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_u_rca48_fa44_and0 = s_CSAwallace_rca24_csa21_csa_component_fa44_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa43_or0;
  assign s_CSAwallace_rca24_u_rca48_fa44_xor1 = s_CSAwallace_rca24_u_rca48_fa44_xor0 ^ s_CSAwallace_rca24_u_rca48_fa43_or0;
  assign s_CSAwallace_rca24_u_rca48_fa44_and1 = s_CSAwallace_rca24_u_rca48_fa44_xor0 & s_CSAwallace_rca24_u_rca48_fa43_or0;
  assign s_CSAwallace_rca24_u_rca48_fa44_or0 = s_CSAwallace_rca24_u_rca48_fa44_and0 | s_CSAwallace_rca24_u_rca48_fa44_and1;
  assign s_CSAwallace_rca24_u_rca48_fa45_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa45_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa44_or0;
  assign s_CSAwallace_rca24_u_rca48_fa45_and0 = s_CSAwallace_rca24_csa21_csa_component_fa45_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa44_or0;
  assign s_CSAwallace_rca24_u_rca48_fa45_xor1 = s_CSAwallace_rca24_u_rca48_fa45_xor0 ^ s_CSAwallace_rca24_u_rca48_fa44_or0;
  assign s_CSAwallace_rca24_u_rca48_fa45_and1 = s_CSAwallace_rca24_u_rca48_fa45_xor0 & s_CSAwallace_rca24_u_rca48_fa44_or0;
  assign s_CSAwallace_rca24_u_rca48_fa45_or0 = s_CSAwallace_rca24_u_rca48_fa45_and0 | s_CSAwallace_rca24_u_rca48_fa45_and1;
  assign s_CSAwallace_rca24_u_rca48_fa46_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa46_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa45_or0;
  assign s_CSAwallace_rca24_u_rca48_fa46_and0 = s_CSAwallace_rca24_csa21_csa_component_fa46_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa45_or0;
  assign s_CSAwallace_rca24_u_rca48_fa46_xor1 = s_CSAwallace_rca24_u_rca48_fa46_xor0 ^ s_CSAwallace_rca24_u_rca48_fa45_or0;
  assign s_CSAwallace_rca24_u_rca48_fa46_and1 = s_CSAwallace_rca24_u_rca48_fa46_xor0 & s_CSAwallace_rca24_u_rca48_fa45_or0;
  assign s_CSAwallace_rca24_u_rca48_fa46_or0 = s_CSAwallace_rca24_u_rca48_fa46_and0 | s_CSAwallace_rca24_u_rca48_fa46_and1;
  assign s_CSAwallace_rca24_u_rca48_fa47_xor0 = s_CSAwallace_rca24_csa21_csa_component_fa47_xor1 ^ s_CSAwallace_rca24_csa21_csa_component_fa46_or0;
  assign s_CSAwallace_rca24_u_rca48_fa47_and0 = s_CSAwallace_rca24_csa21_csa_component_fa47_xor1 & s_CSAwallace_rca24_csa21_csa_component_fa46_or0;
  assign s_CSAwallace_rca24_u_rca48_fa47_xor1 = s_CSAwallace_rca24_u_rca48_fa47_xor0 ^ s_CSAwallace_rca24_u_rca48_fa46_or0;
  assign s_CSAwallace_rca24_u_rca48_fa47_and1 = s_CSAwallace_rca24_u_rca48_fa47_xor0 & s_CSAwallace_rca24_u_rca48_fa46_or0;
  assign s_CSAwallace_rca24_u_rca48_fa47_or0 = s_CSAwallace_rca24_u_rca48_fa47_and0 | s_CSAwallace_rca24_u_rca48_fa47_and1;
  assign s_CSAwallace_rca24_xor0 = ~s_CSAwallace_rca24_u_rca48_fa47_xor1;

  assign s_CSAwallace_rca24_out[0] = s_CSAwallace_rca24_and_0_0;
  assign s_CSAwallace_rca24_out[1] = s_CSAwallace_rca24_csa0_csa_component_fa1_xor0;
  assign s_CSAwallace_rca24_out[2] = s_CSAwallace_rca24_csa8_csa_component_fa2_xor0;
  assign s_CSAwallace_rca24_out[3] = s_CSAwallace_rca24_csa13_csa_component_fa3_xor0;
  assign s_CSAwallace_rca24_out[4] = s_CSAwallace_rca24_csa16_csa_component_fa4_xor0;
  assign s_CSAwallace_rca24_out[5] = s_CSAwallace_rca24_csa18_csa_component_fa5_xor0;
  assign s_CSAwallace_rca24_out[6] = s_CSAwallace_rca24_csa20_csa_component_fa6_xor0;
  assign s_CSAwallace_rca24_out[7] = s_CSAwallace_rca24_csa21_csa_component_fa7_xor0;
  assign s_CSAwallace_rca24_out[8] = s_CSAwallace_rca24_u_rca48_fa8_xor0;
  assign s_CSAwallace_rca24_out[9] = s_CSAwallace_rca24_u_rca48_fa9_xor1;
  assign s_CSAwallace_rca24_out[10] = s_CSAwallace_rca24_u_rca48_fa10_xor1;
  assign s_CSAwallace_rca24_out[11] = s_CSAwallace_rca24_u_rca48_fa11_xor1;
  assign s_CSAwallace_rca24_out[12] = s_CSAwallace_rca24_u_rca48_fa12_xor1;
  assign s_CSAwallace_rca24_out[13] = s_CSAwallace_rca24_u_rca48_fa13_xor1;
  assign s_CSAwallace_rca24_out[14] = s_CSAwallace_rca24_u_rca48_fa14_xor1;
  assign s_CSAwallace_rca24_out[15] = s_CSAwallace_rca24_u_rca48_fa15_xor1;
  assign s_CSAwallace_rca24_out[16] = s_CSAwallace_rca24_u_rca48_fa16_xor1;
  assign s_CSAwallace_rca24_out[17] = s_CSAwallace_rca24_u_rca48_fa17_xor1;
  assign s_CSAwallace_rca24_out[18] = s_CSAwallace_rca24_u_rca48_fa18_xor1;
  assign s_CSAwallace_rca24_out[19] = s_CSAwallace_rca24_u_rca48_fa19_xor1;
  assign s_CSAwallace_rca24_out[20] = s_CSAwallace_rca24_u_rca48_fa20_xor1;
  assign s_CSAwallace_rca24_out[21] = s_CSAwallace_rca24_u_rca48_fa21_xor1;
  assign s_CSAwallace_rca24_out[22] = s_CSAwallace_rca24_u_rca48_fa22_xor1;
  assign s_CSAwallace_rca24_out[23] = s_CSAwallace_rca24_u_rca48_fa23_xor1;
  assign s_CSAwallace_rca24_out[24] = s_CSAwallace_rca24_u_rca48_fa24_xor1;
  assign s_CSAwallace_rca24_out[25] = s_CSAwallace_rca24_u_rca48_fa25_xor1;
  assign s_CSAwallace_rca24_out[26] = s_CSAwallace_rca24_u_rca48_fa26_xor1;
  assign s_CSAwallace_rca24_out[27] = s_CSAwallace_rca24_u_rca48_fa27_xor1;
  assign s_CSAwallace_rca24_out[28] = s_CSAwallace_rca24_u_rca48_fa28_xor1;
  assign s_CSAwallace_rca24_out[29] = s_CSAwallace_rca24_u_rca48_fa29_xor1;
  assign s_CSAwallace_rca24_out[30] = s_CSAwallace_rca24_u_rca48_fa30_xor1;
  assign s_CSAwallace_rca24_out[31] = s_CSAwallace_rca24_u_rca48_fa31_xor1;
  assign s_CSAwallace_rca24_out[32] = s_CSAwallace_rca24_u_rca48_fa32_xor1;
  assign s_CSAwallace_rca24_out[33] = s_CSAwallace_rca24_u_rca48_fa33_xor1;
  assign s_CSAwallace_rca24_out[34] = s_CSAwallace_rca24_u_rca48_fa34_xor1;
  assign s_CSAwallace_rca24_out[35] = s_CSAwallace_rca24_u_rca48_fa35_xor1;
  assign s_CSAwallace_rca24_out[36] = s_CSAwallace_rca24_u_rca48_fa36_xor1;
  assign s_CSAwallace_rca24_out[37] = s_CSAwallace_rca24_u_rca48_fa37_xor1;
  assign s_CSAwallace_rca24_out[38] = s_CSAwallace_rca24_u_rca48_fa38_xor1;
  assign s_CSAwallace_rca24_out[39] = s_CSAwallace_rca24_u_rca48_fa39_xor1;
  assign s_CSAwallace_rca24_out[40] = s_CSAwallace_rca24_u_rca48_fa40_xor1;
  assign s_CSAwallace_rca24_out[41] = s_CSAwallace_rca24_u_rca48_fa41_xor1;
  assign s_CSAwallace_rca24_out[42] = s_CSAwallace_rca24_u_rca48_fa42_xor1;
  assign s_CSAwallace_rca24_out[43] = s_CSAwallace_rca24_u_rca48_fa43_xor1;
  assign s_CSAwallace_rca24_out[44] = s_CSAwallace_rca24_u_rca48_fa44_xor1;
  assign s_CSAwallace_rca24_out[45] = s_CSAwallace_rca24_u_rca48_fa45_xor1;
  assign s_CSAwallace_rca24_out[46] = s_CSAwallace_rca24_u_rca48_fa46_xor1;
  assign s_CSAwallace_rca24_out[47] = s_CSAwallace_rca24_xor0;
endmodule