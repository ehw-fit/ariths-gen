module s_csamul_pg_rca4(input [3:0] a, input [3:0] b, output [7:0] s_csamul_pg_rca4_out);
  wire s_csamul_pg_rca4_and0_0;
  wire s_csamul_pg_rca4_and1_0;
  wire s_csamul_pg_rca4_and2_0;
  wire s_csamul_pg_rca4_nand3_0;
  wire s_csamul_pg_rca4_and0_1;
  wire s_csamul_pg_rca4_ha0_1_xor0;
  wire s_csamul_pg_rca4_ha0_1_and0;
  wire s_csamul_pg_rca4_and1_1;
  wire s_csamul_pg_rca4_ha1_1_xor0;
  wire s_csamul_pg_rca4_ha1_1_and0;
  wire s_csamul_pg_rca4_and2_1;
  wire s_csamul_pg_rca4_ha2_1_xor0;
  wire s_csamul_pg_rca4_ha2_1_and0;
  wire s_csamul_pg_rca4_nand3_1;
  wire s_csamul_pg_rca4_ha3_1_xor0;
  wire s_csamul_pg_rca4_and0_2;
  wire s_csamul_pg_rca4_fa0_2_xor0;
  wire s_csamul_pg_rca4_fa0_2_and0;
  wire s_csamul_pg_rca4_fa0_2_xor1;
  wire s_csamul_pg_rca4_fa0_2_and1;
  wire s_csamul_pg_rca4_fa0_2_or0;
  wire s_csamul_pg_rca4_and1_2;
  wire s_csamul_pg_rca4_fa1_2_xor0;
  wire s_csamul_pg_rca4_fa1_2_and0;
  wire s_csamul_pg_rca4_fa1_2_xor1;
  wire s_csamul_pg_rca4_fa1_2_and1;
  wire s_csamul_pg_rca4_fa1_2_or0;
  wire s_csamul_pg_rca4_and2_2;
  wire s_csamul_pg_rca4_fa2_2_xor0;
  wire s_csamul_pg_rca4_fa2_2_and0;
  wire s_csamul_pg_rca4_fa2_2_xor1;
  wire s_csamul_pg_rca4_fa2_2_and1;
  wire s_csamul_pg_rca4_fa2_2_or0;
  wire s_csamul_pg_rca4_nand3_2;
  wire s_csamul_pg_rca4_ha3_2_xor0;
  wire s_csamul_pg_rca4_ha3_2_and0;
  wire s_csamul_pg_rca4_nand0_3;
  wire s_csamul_pg_rca4_fa0_3_xor0;
  wire s_csamul_pg_rca4_fa0_3_and0;
  wire s_csamul_pg_rca4_fa0_3_xor1;
  wire s_csamul_pg_rca4_fa0_3_and1;
  wire s_csamul_pg_rca4_fa0_3_or0;
  wire s_csamul_pg_rca4_nand1_3;
  wire s_csamul_pg_rca4_fa1_3_xor0;
  wire s_csamul_pg_rca4_fa1_3_and0;
  wire s_csamul_pg_rca4_fa1_3_xor1;
  wire s_csamul_pg_rca4_fa1_3_and1;
  wire s_csamul_pg_rca4_fa1_3_or0;
  wire s_csamul_pg_rca4_nand2_3;
  wire s_csamul_pg_rca4_fa2_3_xor0;
  wire s_csamul_pg_rca4_fa2_3_and0;
  wire s_csamul_pg_rca4_fa2_3_xor1;
  wire s_csamul_pg_rca4_fa2_3_and1;
  wire s_csamul_pg_rca4_fa2_3_or0;
  wire s_csamul_pg_rca4_and3_3;
  wire s_csamul_pg_rca4_ha3_3_xor0;
  wire s_csamul_pg_rca4_ha3_3_and0;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa0_xor0;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa0_and0;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa1_xor0;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa1_and0;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa1_xor1;
  wire s_csamul_pg_rca4_u_pg_rca4_and1;
  wire s_csamul_pg_rca4_u_pg_rca4_or1;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa2_xor0;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa2_and0;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa2_xor1;
  wire s_csamul_pg_rca4_u_pg_rca4_and2;
  wire s_csamul_pg_rca4_u_pg_rca4_or2;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa3_xor0;
  wire s_csamul_pg_rca4_u_pg_rca4_pg_fa3_xor1;
  wire s_csamul_pg_rca4_u_pg_rca4_and3;
  wire s_csamul_pg_rca4_u_pg_rca4_or3;

  assign s_csamul_pg_rca4_and0_0 = a[0] & b[0];
  assign s_csamul_pg_rca4_and1_0 = a[1] & b[0];
  assign s_csamul_pg_rca4_and2_0 = a[2] & b[0];
  assign s_csamul_pg_rca4_nand3_0 = ~(a[3] & b[0]);
  assign s_csamul_pg_rca4_and0_1 = a[0] & b[1];
  assign s_csamul_pg_rca4_ha0_1_xor0 = s_csamul_pg_rca4_and0_1 ^ s_csamul_pg_rca4_and1_0;
  assign s_csamul_pg_rca4_ha0_1_and0 = s_csamul_pg_rca4_and0_1 & s_csamul_pg_rca4_and1_0;
  assign s_csamul_pg_rca4_and1_1 = a[1] & b[1];
  assign s_csamul_pg_rca4_ha1_1_xor0 = s_csamul_pg_rca4_and1_1 ^ s_csamul_pg_rca4_and2_0;
  assign s_csamul_pg_rca4_ha1_1_and0 = s_csamul_pg_rca4_and1_1 & s_csamul_pg_rca4_and2_0;
  assign s_csamul_pg_rca4_and2_1 = a[2] & b[1];
  assign s_csamul_pg_rca4_ha2_1_xor0 = s_csamul_pg_rca4_and2_1 ^ s_csamul_pg_rca4_nand3_0;
  assign s_csamul_pg_rca4_ha2_1_and0 = s_csamul_pg_rca4_and2_1 & s_csamul_pg_rca4_nand3_0;
  assign s_csamul_pg_rca4_nand3_1 = ~(a[3] & b[1]);
  assign s_csamul_pg_rca4_ha3_1_xor0 = ~s_csamul_pg_rca4_nand3_1;
  assign s_csamul_pg_rca4_and0_2 = a[0] & b[2];
  assign s_csamul_pg_rca4_fa0_2_xor0 = s_csamul_pg_rca4_and0_2 ^ s_csamul_pg_rca4_ha1_1_xor0;
  assign s_csamul_pg_rca4_fa0_2_and0 = s_csamul_pg_rca4_and0_2 & s_csamul_pg_rca4_ha1_1_xor0;
  assign s_csamul_pg_rca4_fa0_2_xor1 = s_csamul_pg_rca4_fa0_2_xor0 ^ s_csamul_pg_rca4_ha0_1_and0;
  assign s_csamul_pg_rca4_fa0_2_and1 = s_csamul_pg_rca4_fa0_2_xor0 & s_csamul_pg_rca4_ha0_1_and0;
  assign s_csamul_pg_rca4_fa0_2_or0 = s_csamul_pg_rca4_fa0_2_and0 | s_csamul_pg_rca4_fa0_2_and1;
  assign s_csamul_pg_rca4_and1_2 = a[1] & b[2];
  assign s_csamul_pg_rca4_fa1_2_xor0 = s_csamul_pg_rca4_and1_2 ^ s_csamul_pg_rca4_ha2_1_xor0;
  assign s_csamul_pg_rca4_fa1_2_and0 = s_csamul_pg_rca4_and1_2 & s_csamul_pg_rca4_ha2_1_xor0;
  assign s_csamul_pg_rca4_fa1_2_xor1 = s_csamul_pg_rca4_fa1_2_xor0 ^ s_csamul_pg_rca4_ha1_1_and0;
  assign s_csamul_pg_rca4_fa1_2_and1 = s_csamul_pg_rca4_fa1_2_xor0 & s_csamul_pg_rca4_ha1_1_and0;
  assign s_csamul_pg_rca4_fa1_2_or0 = s_csamul_pg_rca4_fa1_2_and0 | s_csamul_pg_rca4_fa1_2_and1;
  assign s_csamul_pg_rca4_and2_2 = a[2] & b[2];
  assign s_csamul_pg_rca4_fa2_2_xor0 = s_csamul_pg_rca4_and2_2 ^ s_csamul_pg_rca4_ha3_1_xor0;
  assign s_csamul_pg_rca4_fa2_2_and0 = s_csamul_pg_rca4_and2_2 & s_csamul_pg_rca4_ha3_1_xor0;
  assign s_csamul_pg_rca4_fa2_2_xor1 = s_csamul_pg_rca4_fa2_2_xor0 ^ s_csamul_pg_rca4_ha2_1_and0;
  assign s_csamul_pg_rca4_fa2_2_and1 = s_csamul_pg_rca4_fa2_2_xor0 & s_csamul_pg_rca4_ha2_1_and0;
  assign s_csamul_pg_rca4_fa2_2_or0 = s_csamul_pg_rca4_fa2_2_and0 | s_csamul_pg_rca4_fa2_2_and1;
  assign s_csamul_pg_rca4_nand3_2 = ~(a[3] & b[2]);
  assign s_csamul_pg_rca4_ha3_2_xor0 = s_csamul_pg_rca4_nand3_2 ^ s_csamul_pg_rca4_nand3_1;
  assign s_csamul_pg_rca4_ha3_2_and0 = s_csamul_pg_rca4_nand3_2 & s_csamul_pg_rca4_nand3_1;
  assign s_csamul_pg_rca4_nand0_3 = ~(a[0] & b[3]);
  assign s_csamul_pg_rca4_fa0_3_xor0 = s_csamul_pg_rca4_nand0_3 ^ s_csamul_pg_rca4_fa1_2_xor1;
  assign s_csamul_pg_rca4_fa0_3_and0 = s_csamul_pg_rca4_nand0_3 & s_csamul_pg_rca4_fa1_2_xor1;
  assign s_csamul_pg_rca4_fa0_3_xor1 = s_csamul_pg_rca4_fa0_3_xor0 ^ s_csamul_pg_rca4_fa0_2_or0;
  assign s_csamul_pg_rca4_fa0_3_and1 = s_csamul_pg_rca4_fa0_3_xor0 & s_csamul_pg_rca4_fa0_2_or0;
  assign s_csamul_pg_rca4_fa0_3_or0 = s_csamul_pg_rca4_fa0_3_and0 | s_csamul_pg_rca4_fa0_3_and1;
  assign s_csamul_pg_rca4_nand1_3 = ~(a[1] & b[3]);
  assign s_csamul_pg_rca4_fa1_3_xor0 = s_csamul_pg_rca4_nand1_3 ^ s_csamul_pg_rca4_fa2_2_xor1;
  assign s_csamul_pg_rca4_fa1_3_and0 = s_csamul_pg_rca4_nand1_3 & s_csamul_pg_rca4_fa2_2_xor1;
  assign s_csamul_pg_rca4_fa1_3_xor1 = s_csamul_pg_rca4_fa1_3_xor0 ^ s_csamul_pg_rca4_fa1_2_or0;
  assign s_csamul_pg_rca4_fa1_3_and1 = s_csamul_pg_rca4_fa1_3_xor0 & s_csamul_pg_rca4_fa1_2_or0;
  assign s_csamul_pg_rca4_fa1_3_or0 = s_csamul_pg_rca4_fa1_3_and0 | s_csamul_pg_rca4_fa1_3_and1;
  assign s_csamul_pg_rca4_nand2_3 = ~(a[2] & b[3]);
  assign s_csamul_pg_rca4_fa2_3_xor0 = s_csamul_pg_rca4_nand2_3 ^ s_csamul_pg_rca4_ha3_2_xor0;
  assign s_csamul_pg_rca4_fa2_3_and0 = s_csamul_pg_rca4_nand2_3 & s_csamul_pg_rca4_ha3_2_xor0;
  assign s_csamul_pg_rca4_fa2_3_xor1 = s_csamul_pg_rca4_fa2_3_xor0 ^ s_csamul_pg_rca4_fa2_2_or0;
  assign s_csamul_pg_rca4_fa2_3_and1 = s_csamul_pg_rca4_fa2_3_xor0 & s_csamul_pg_rca4_fa2_2_or0;
  assign s_csamul_pg_rca4_fa2_3_or0 = s_csamul_pg_rca4_fa2_3_and0 | s_csamul_pg_rca4_fa2_3_and1;
  assign s_csamul_pg_rca4_and3_3 = a[3] & b[3];
  assign s_csamul_pg_rca4_ha3_3_xor0 = s_csamul_pg_rca4_and3_3 ^ s_csamul_pg_rca4_ha3_2_and0;
  assign s_csamul_pg_rca4_ha3_3_and0 = s_csamul_pg_rca4_and3_3 & s_csamul_pg_rca4_ha3_2_and0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa0_xor0 = s_csamul_pg_rca4_fa1_3_xor1 ^ s_csamul_pg_rca4_fa0_3_or0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa0_and0 = s_csamul_pg_rca4_fa1_3_xor1 & s_csamul_pg_rca4_fa0_3_or0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa1_xor0 = s_csamul_pg_rca4_fa2_3_xor1 ^ s_csamul_pg_rca4_fa1_3_or0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa1_and0 = s_csamul_pg_rca4_fa2_3_xor1 & s_csamul_pg_rca4_fa1_3_or0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa1_xor1 = s_csamul_pg_rca4_u_pg_rca4_pg_fa1_xor0 ^ s_csamul_pg_rca4_u_pg_rca4_pg_fa0_and0;
  assign s_csamul_pg_rca4_u_pg_rca4_and1 = s_csamul_pg_rca4_u_pg_rca4_pg_fa0_and0 & s_csamul_pg_rca4_u_pg_rca4_pg_fa1_xor0;
  assign s_csamul_pg_rca4_u_pg_rca4_or1 = s_csamul_pg_rca4_u_pg_rca4_and1 | s_csamul_pg_rca4_u_pg_rca4_pg_fa1_and0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa2_xor0 = s_csamul_pg_rca4_ha3_3_xor0 ^ s_csamul_pg_rca4_fa2_3_or0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa2_and0 = s_csamul_pg_rca4_ha3_3_xor0 & s_csamul_pg_rca4_fa2_3_or0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa2_xor1 = s_csamul_pg_rca4_u_pg_rca4_pg_fa2_xor0 ^ s_csamul_pg_rca4_u_pg_rca4_or1;
  assign s_csamul_pg_rca4_u_pg_rca4_and2 = s_csamul_pg_rca4_u_pg_rca4_or1 & s_csamul_pg_rca4_u_pg_rca4_pg_fa2_xor0;
  assign s_csamul_pg_rca4_u_pg_rca4_or2 = s_csamul_pg_rca4_u_pg_rca4_and2 | s_csamul_pg_rca4_u_pg_rca4_pg_fa2_and0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa3_xor0 = ~s_csamul_pg_rca4_ha3_3_and0;
  assign s_csamul_pg_rca4_u_pg_rca4_pg_fa3_xor1 = s_csamul_pg_rca4_u_pg_rca4_pg_fa3_xor0 ^ s_csamul_pg_rca4_u_pg_rca4_or2;
  assign s_csamul_pg_rca4_u_pg_rca4_and3 = s_csamul_pg_rca4_u_pg_rca4_or2 & s_csamul_pg_rca4_u_pg_rca4_pg_fa3_xor0;
  assign s_csamul_pg_rca4_u_pg_rca4_or3 = s_csamul_pg_rca4_u_pg_rca4_and3 | s_csamul_pg_rca4_ha3_3_and0;

  assign s_csamul_pg_rca4_out[0] = s_csamul_pg_rca4_and0_0;
  assign s_csamul_pg_rca4_out[1] = s_csamul_pg_rca4_ha0_1_xor0;
  assign s_csamul_pg_rca4_out[2] = s_csamul_pg_rca4_fa0_2_xor1;
  assign s_csamul_pg_rca4_out[3] = s_csamul_pg_rca4_fa0_3_xor1;
  assign s_csamul_pg_rca4_out[4] = s_csamul_pg_rca4_u_pg_rca4_pg_fa0_xor0;
  assign s_csamul_pg_rca4_out[5] = s_csamul_pg_rca4_u_pg_rca4_pg_fa1_xor1;
  assign s_csamul_pg_rca4_out[6] = s_csamul_pg_rca4_u_pg_rca4_pg_fa2_xor1;
  assign s_csamul_pg_rca4_out[7] = s_csamul_pg_rca4_u_pg_rca4_pg_fa3_xor1;
endmodule