module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module pg_fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] pg_fa_xor0, output [0:0] pg_fa_and0, output [0:0] pg_fa_xor1);
  xor_gate xor_gate_pg_fa_xor0(a[0], b[0], pg_fa_xor0);
  and_gate and_gate_pg_fa_and0(a[0], b[0], pg_fa_and0);
  xor_gate xor_gate_pg_fa_xor1(pg_fa_xor0[0], cin[0], pg_fa_xor1);
endmodule

module h_s_pg_rca16(input [15:0] a, input [15:0] b, output [16:0] h_s_pg_rca16_out);
  wire [0:0] h_s_pg_rca16_pg_fa0_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa0_and0;
  wire [0:0] h_s_pg_rca16_pg_fa1_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa1_and0;
  wire [0:0] h_s_pg_rca16_pg_fa1_xor1;
  wire [0:0] h_s_pg_rca16_and1;
  wire [0:0] h_s_pg_rca16_or1;
  wire [0:0] h_s_pg_rca16_pg_fa2_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa2_and0;
  wire [0:0] h_s_pg_rca16_pg_fa2_xor1;
  wire [0:0] h_s_pg_rca16_and2;
  wire [0:0] h_s_pg_rca16_or2;
  wire [0:0] h_s_pg_rca16_pg_fa3_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa3_and0;
  wire [0:0] h_s_pg_rca16_pg_fa3_xor1;
  wire [0:0] h_s_pg_rca16_and3;
  wire [0:0] h_s_pg_rca16_or3;
  wire [0:0] h_s_pg_rca16_pg_fa4_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa4_and0;
  wire [0:0] h_s_pg_rca16_pg_fa4_xor1;
  wire [0:0] h_s_pg_rca16_and4;
  wire [0:0] h_s_pg_rca16_or4;
  wire [0:0] h_s_pg_rca16_pg_fa5_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa5_and0;
  wire [0:0] h_s_pg_rca16_pg_fa5_xor1;
  wire [0:0] h_s_pg_rca16_and5;
  wire [0:0] h_s_pg_rca16_or5;
  wire [0:0] h_s_pg_rca16_pg_fa6_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa6_and0;
  wire [0:0] h_s_pg_rca16_pg_fa6_xor1;
  wire [0:0] h_s_pg_rca16_and6;
  wire [0:0] h_s_pg_rca16_or6;
  wire [0:0] h_s_pg_rca16_pg_fa7_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa7_and0;
  wire [0:0] h_s_pg_rca16_pg_fa7_xor1;
  wire [0:0] h_s_pg_rca16_and7;
  wire [0:0] h_s_pg_rca16_or7;
  wire [0:0] h_s_pg_rca16_pg_fa8_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa8_and0;
  wire [0:0] h_s_pg_rca16_pg_fa8_xor1;
  wire [0:0] h_s_pg_rca16_and8;
  wire [0:0] h_s_pg_rca16_or8;
  wire [0:0] h_s_pg_rca16_pg_fa9_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa9_and0;
  wire [0:0] h_s_pg_rca16_pg_fa9_xor1;
  wire [0:0] h_s_pg_rca16_and9;
  wire [0:0] h_s_pg_rca16_or9;
  wire [0:0] h_s_pg_rca16_pg_fa10_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa10_and0;
  wire [0:0] h_s_pg_rca16_pg_fa10_xor1;
  wire [0:0] h_s_pg_rca16_and10;
  wire [0:0] h_s_pg_rca16_or10;
  wire [0:0] h_s_pg_rca16_pg_fa11_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa11_and0;
  wire [0:0] h_s_pg_rca16_pg_fa11_xor1;
  wire [0:0] h_s_pg_rca16_and11;
  wire [0:0] h_s_pg_rca16_or11;
  wire [0:0] h_s_pg_rca16_pg_fa12_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa12_and0;
  wire [0:0] h_s_pg_rca16_pg_fa12_xor1;
  wire [0:0] h_s_pg_rca16_and12;
  wire [0:0] h_s_pg_rca16_or12;
  wire [0:0] h_s_pg_rca16_pg_fa13_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa13_and0;
  wire [0:0] h_s_pg_rca16_pg_fa13_xor1;
  wire [0:0] h_s_pg_rca16_and13;
  wire [0:0] h_s_pg_rca16_or13;
  wire [0:0] h_s_pg_rca16_pg_fa14_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa14_and0;
  wire [0:0] h_s_pg_rca16_pg_fa14_xor1;
  wire [0:0] h_s_pg_rca16_and14;
  wire [0:0] h_s_pg_rca16_or14;
  wire [0:0] h_s_pg_rca16_pg_fa15_xor0;
  wire [0:0] h_s_pg_rca16_pg_fa15_and0;
  wire [0:0] h_s_pg_rca16_pg_fa15_xor1;
  wire [0:0] h_s_pg_rca16_and15;
  wire [0:0] h_s_pg_rca16_or15;
  wire [0:0] h_s_pg_rca16_xor0;
  wire [0:0] h_s_pg_rca16_xor1;

  pg_fa pg_fa_h_s_pg_rca16_pg_fa0_out(a[0], b[0], 1'b0, h_s_pg_rca16_pg_fa0_xor0, h_s_pg_rca16_pg_fa0_and0);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa1_out(a[1], b[1], h_s_pg_rca16_pg_fa0_and0[0], h_s_pg_rca16_pg_fa1_xor0, h_s_pg_rca16_pg_fa1_and0, h_s_pg_rca16_pg_fa1_xor1);
  and_gate and_gate_h_s_pg_rca16_and1(h_s_pg_rca16_pg_fa0_and0[0], h_s_pg_rca16_pg_fa1_xor0[0], h_s_pg_rca16_and1);
  or_gate or_gate_h_s_pg_rca16_or1(h_s_pg_rca16_and1[0], h_s_pg_rca16_pg_fa1_and0[0], h_s_pg_rca16_or1);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa2_out(a[2], b[2], h_s_pg_rca16_or1[0], h_s_pg_rca16_pg_fa2_xor0, h_s_pg_rca16_pg_fa2_and0, h_s_pg_rca16_pg_fa2_xor1);
  and_gate and_gate_h_s_pg_rca16_and2(h_s_pg_rca16_or1[0], h_s_pg_rca16_pg_fa2_xor0[0], h_s_pg_rca16_and2);
  or_gate or_gate_h_s_pg_rca16_or2(h_s_pg_rca16_and2[0], h_s_pg_rca16_pg_fa2_and0[0], h_s_pg_rca16_or2);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa3_out(a[3], b[3], h_s_pg_rca16_or2[0], h_s_pg_rca16_pg_fa3_xor0, h_s_pg_rca16_pg_fa3_and0, h_s_pg_rca16_pg_fa3_xor1);
  and_gate and_gate_h_s_pg_rca16_and3(h_s_pg_rca16_or2[0], h_s_pg_rca16_pg_fa3_xor0[0], h_s_pg_rca16_and3);
  or_gate or_gate_h_s_pg_rca16_or3(h_s_pg_rca16_and3[0], h_s_pg_rca16_pg_fa3_and0[0], h_s_pg_rca16_or3);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa4_out(a[4], b[4], h_s_pg_rca16_or3[0], h_s_pg_rca16_pg_fa4_xor0, h_s_pg_rca16_pg_fa4_and0, h_s_pg_rca16_pg_fa4_xor1);
  and_gate and_gate_h_s_pg_rca16_and4(h_s_pg_rca16_or3[0], h_s_pg_rca16_pg_fa4_xor0[0], h_s_pg_rca16_and4);
  or_gate or_gate_h_s_pg_rca16_or4(h_s_pg_rca16_and4[0], h_s_pg_rca16_pg_fa4_and0[0], h_s_pg_rca16_or4);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa5_out(a[5], b[5], h_s_pg_rca16_or4[0], h_s_pg_rca16_pg_fa5_xor0, h_s_pg_rca16_pg_fa5_and0, h_s_pg_rca16_pg_fa5_xor1);
  and_gate and_gate_h_s_pg_rca16_and5(h_s_pg_rca16_or4[0], h_s_pg_rca16_pg_fa5_xor0[0], h_s_pg_rca16_and5);
  or_gate or_gate_h_s_pg_rca16_or5(h_s_pg_rca16_and5[0], h_s_pg_rca16_pg_fa5_and0[0], h_s_pg_rca16_or5);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa6_out(a[6], b[6], h_s_pg_rca16_or5[0], h_s_pg_rca16_pg_fa6_xor0, h_s_pg_rca16_pg_fa6_and0, h_s_pg_rca16_pg_fa6_xor1);
  and_gate and_gate_h_s_pg_rca16_and6(h_s_pg_rca16_or5[0], h_s_pg_rca16_pg_fa6_xor0[0], h_s_pg_rca16_and6);
  or_gate or_gate_h_s_pg_rca16_or6(h_s_pg_rca16_and6[0], h_s_pg_rca16_pg_fa6_and0[0], h_s_pg_rca16_or6);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa7_out(a[7], b[7], h_s_pg_rca16_or6[0], h_s_pg_rca16_pg_fa7_xor0, h_s_pg_rca16_pg_fa7_and0, h_s_pg_rca16_pg_fa7_xor1);
  and_gate and_gate_h_s_pg_rca16_and7(h_s_pg_rca16_or6[0], h_s_pg_rca16_pg_fa7_xor0[0], h_s_pg_rca16_and7);
  or_gate or_gate_h_s_pg_rca16_or7(h_s_pg_rca16_and7[0], h_s_pg_rca16_pg_fa7_and0[0], h_s_pg_rca16_or7);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa8_out(a[8], b[8], h_s_pg_rca16_or7[0], h_s_pg_rca16_pg_fa8_xor0, h_s_pg_rca16_pg_fa8_and0, h_s_pg_rca16_pg_fa8_xor1);
  and_gate and_gate_h_s_pg_rca16_and8(h_s_pg_rca16_or7[0], h_s_pg_rca16_pg_fa8_xor0[0], h_s_pg_rca16_and8);
  or_gate or_gate_h_s_pg_rca16_or8(h_s_pg_rca16_and8[0], h_s_pg_rca16_pg_fa8_and0[0], h_s_pg_rca16_or8);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa9_out(a[9], b[9], h_s_pg_rca16_or8[0], h_s_pg_rca16_pg_fa9_xor0, h_s_pg_rca16_pg_fa9_and0, h_s_pg_rca16_pg_fa9_xor1);
  and_gate and_gate_h_s_pg_rca16_and9(h_s_pg_rca16_or8[0], h_s_pg_rca16_pg_fa9_xor0[0], h_s_pg_rca16_and9);
  or_gate or_gate_h_s_pg_rca16_or9(h_s_pg_rca16_and9[0], h_s_pg_rca16_pg_fa9_and0[0], h_s_pg_rca16_or9);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa10_out(a[10], b[10], h_s_pg_rca16_or9[0], h_s_pg_rca16_pg_fa10_xor0, h_s_pg_rca16_pg_fa10_and0, h_s_pg_rca16_pg_fa10_xor1);
  and_gate and_gate_h_s_pg_rca16_and10(h_s_pg_rca16_or9[0], h_s_pg_rca16_pg_fa10_xor0[0], h_s_pg_rca16_and10);
  or_gate or_gate_h_s_pg_rca16_or10(h_s_pg_rca16_and10[0], h_s_pg_rca16_pg_fa10_and0[0], h_s_pg_rca16_or10);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa11_out(a[11], b[11], h_s_pg_rca16_or10[0], h_s_pg_rca16_pg_fa11_xor0, h_s_pg_rca16_pg_fa11_and0, h_s_pg_rca16_pg_fa11_xor1);
  and_gate and_gate_h_s_pg_rca16_and11(h_s_pg_rca16_or10[0], h_s_pg_rca16_pg_fa11_xor0[0], h_s_pg_rca16_and11);
  or_gate or_gate_h_s_pg_rca16_or11(h_s_pg_rca16_and11[0], h_s_pg_rca16_pg_fa11_and0[0], h_s_pg_rca16_or11);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa12_out(a[12], b[12], h_s_pg_rca16_or11[0], h_s_pg_rca16_pg_fa12_xor0, h_s_pg_rca16_pg_fa12_and0, h_s_pg_rca16_pg_fa12_xor1);
  and_gate and_gate_h_s_pg_rca16_and12(h_s_pg_rca16_or11[0], h_s_pg_rca16_pg_fa12_xor0[0], h_s_pg_rca16_and12);
  or_gate or_gate_h_s_pg_rca16_or12(h_s_pg_rca16_and12[0], h_s_pg_rca16_pg_fa12_and0[0], h_s_pg_rca16_or12);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa13_out(a[13], b[13], h_s_pg_rca16_or12[0], h_s_pg_rca16_pg_fa13_xor0, h_s_pg_rca16_pg_fa13_and0, h_s_pg_rca16_pg_fa13_xor1);
  and_gate and_gate_h_s_pg_rca16_and13(h_s_pg_rca16_or12[0], h_s_pg_rca16_pg_fa13_xor0[0], h_s_pg_rca16_and13);
  or_gate or_gate_h_s_pg_rca16_or13(h_s_pg_rca16_and13[0], h_s_pg_rca16_pg_fa13_and0[0], h_s_pg_rca16_or13);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa14_out(a[14], b[14], h_s_pg_rca16_or13[0], h_s_pg_rca16_pg_fa14_xor0, h_s_pg_rca16_pg_fa14_and0, h_s_pg_rca16_pg_fa14_xor1);
  and_gate and_gate_h_s_pg_rca16_and14(h_s_pg_rca16_or13[0], h_s_pg_rca16_pg_fa14_xor0[0], h_s_pg_rca16_and14);
  or_gate or_gate_h_s_pg_rca16_or14(h_s_pg_rca16_and14[0], h_s_pg_rca16_pg_fa14_and0[0], h_s_pg_rca16_or14);
  pg_fa pg_fa_h_s_pg_rca16_pg_fa15_out(a[15], b[15], h_s_pg_rca16_or14[0], h_s_pg_rca16_pg_fa15_xor0, h_s_pg_rca16_pg_fa15_and0, h_s_pg_rca16_pg_fa15_xor1);
  and_gate and_gate_h_s_pg_rca16_and15(h_s_pg_rca16_or14[0], h_s_pg_rca16_pg_fa15_xor0[0], h_s_pg_rca16_and15);
  or_gate or_gate_h_s_pg_rca16_or15(h_s_pg_rca16_and15[0], h_s_pg_rca16_pg_fa15_and0[0], h_s_pg_rca16_or15);
  xor_gate xor_gate_h_s_pg_rca16_xor0(a[15], b[15], h_s_pg_rca16_xor0);
  xor_gate xor_gate_h_s_pg_rca16_xor1(h_s_pg_rca16_xor0[0], h_s_pg_rca16_or15[0], h_s_pg_rca16_xor1);

  assign h_s_pg_rca16_out[0] = h_s_pg_rca16_pg_fa0_xor0[0];
  assign h_s_pg_rca16_out[1] = h_s_pg_rca16_pg_fa1_xor1[0];
  assign h_s_pg_rca16_out[2] = h_s_pg_rca16_pg_fa2_xor1[0];
  assign h_s_pg_rca16_out[3] = h_s_pg_rca16_pg_fa3_xor1[0];
  assign h_s_pg_rca16_out[4] = h_s_pg_rca16_pg_fa4_xor1[0];
  assign h_s_pg_rca16_out[5] = h_s_pg_rca16_pg_fa5_xor1[0];
  assign h_s_pg_rca16_out[6] = h_s_pg_rca16_pg_fa6_xor1[0];
  assign h_s_pg_rca16_out[7] = h_s_pg_rca16_pg_fa7_xor1[0];
  assign h_s_pg_rca16_out[8] = h_s_pg_rca16_pg_fa8_xor1[0];
  assign h_s_pg_rca16_out[9] = h_s_pg_rca16_pg_fa9_xor1[0];
  assign h_s_pg_rca16_out[10] = h_s_pg_rca16_pg_fa10_xor1[0];
  assign h_s_pg_rca16_out[11] = h_s_pg_rca16_pg_fa11_xor1[0];
  assign h_s_pg_rca16_out[12] = h_s_pg_rca16_pg_fa12_xor1[0];
  assign h_s_pg_rca16_out[13] = h_s_pg_rca16_pg_fa13_xor1[0];
  assign h_s_pg_rca16_out[14] = h_s_pg_rca16_pg_fa14_xor1[0];
  assign h_s_pg_rca16_out[15] = h_s_pg_rca16_pg_fa15_xor1[0];
  assign h_s_pg_rca16_out[16] = h_s_pg_rca16_xor1[0];
endmodule