module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module u_cska22(input [21:0] a, input [21:0] b, output [22:0] u_cska22_out);
  wire [0:0] u_cska22_xor0;
  wire [0:0] u_cska22_ha0_xor0;
  wire [0:0] u_cska22_ha0_and0;
  wire [0:0] u_cska22_xor1;
  wire [0:0] u_cska22_fa0_xor1;
  wire [0:0] u_cska22_fa0_or0;
  wire [0:0] u_cska22_xor2;
  wire [0:0] u_cska22_fa1_xor1;
  wire [0:0] u_cska22_fa1_or0;
  wire [0:0] u_cska22_xor3;
  wire [0:0] u_cska22_fa2_xor1;
  wire [0:0] u_cska22_fa2_or0;
  wire [0:0] u_cska22_and_propagate00;
  wire [0:0] u_cska22_and_propagate01;
  wire [0:0] u_cska22_and_propagate02;
  wire [0:0] u_cska22_mux2to10_and1;
  wire [0:0] u_cska22_xor4;
  wire [0:0] u_cska22_fa3_xor1;
  wire [0:0] u_cska22_fa3_or0;
  wire [0:0] u_cska22_xor5;
  wire [0:0] u_cska22_fa4_xor1;
  wire [0:0] u_cska22_fa4_or0;
  wire [0:0] u_cska22_xor6;
  wire [0:0] u_cska22_fa5_xor1;
  wire [0:0] u_cska22_fa5_or0;
  wire [0:0] u_cska22_xor7;
  wire [0:0] u_cska22_fa6_xor1;
  wire [0:0] u_cska22_fa6_or0;
  wire [0:0] u_cska22_and_propagate13;
  wire [0:0] u_cska22_and_propagate14;
  wire [0:0] u_cska22_and_propagate15;
  wire [0:0] u_cska22_mux2to11_xor0;
  wire [0:0] u_cska22_xor8;
  wire [0:0] u_cska22_fa7_xor1;
  wire [0:0] u_cska22_fa7_or0;
  wire [0:0] u_cska22_xor9;
  wire [0:0] u_cska22_fa8_xor1;
  wire [0:0] u_cska22_fa8_or0;
  wire [0:0] u_cska22_xor10;
  wire [0:0] u_cska22_fa9_xor1;
  wire [0:0] u_cska22_fa9_or0;
  wire [0:0] u_cska22_xor11;
  wire [0:0] u_cska22_fa10_xor1;
  wire [0:0] u_cska22_fa10_or0;
  wire [0:0] u_cska22_and_propagate26;
  wire [0:0] u_cska22_and_propagate27;
  wire [0:0] u_cska22_and_propagate28;
  wire [0:0] u_cska22_mux2to12_xor0;
  wire [0:0] u_cska22_xor12;
  wire [0:0] u_cska22_fa11_xor1;
  wire [0:0] u_cska22_fa11_or0;
  wire [0:0] u_cska22_xor13;
  wire [0:0] u_cska22_fa12_xor1;
  wire [0:0] u_cska22_fa12_or0;
  wire [0:0] u_cska22_xor14;
  wire [0:0] u_cska22_fa13_xor1;
  wire [0:0] u_cska22_fa13_or0;
  wire [0:0] u_cska22_xor15;
  wire [0:0] u_cska22_fa14_xor1;
  wire [0:0] u_cska22_fa14_or0;
  wire [0:0] u_cska22_and_propagate39;
  wire [0:0] u_cska22_and_propagate310;
  wire [0:0] u_cska22_and_propagate311;
  wire [0:0] u_cska22_mux2to13_xor0;
  wire [0:0] u_cska22_xor16;
  wire [0:0] u_cska22_fa15_xor1;
  wire [0:0] u_cska22_fa15_or0;
  wire [0:0] u_cska22_xor17;
  wire [0:0] u_cska22_fa16_xor1;
  wire [0:0] u_cska22_fa16_or0;
  wire [0:0] u_cska22_xor18;
  wire [0:0] u_cska22_fa17_xor1;
  wire [0:0] u_cska22_fa17_or0;
  wire [0:0] u_cska22_xor19;
  wire [0:0] u_cska22_fa18_xor1;
  wire [0:0] u_cska22_fa18_or0;
  wire [0:0] u_cska22_and_propagate412;
  wire [0:0] u_cska22_and_propagate413;
  wire [0:0] u_cska22_and_propagate414;
  wire [0:0] u_cska22_mux2to14_xor0;
  wire [0:0] u_cska22_xor20;
  wire [0:0] u_cska22_fa19_xor1;
  wire [0:0] u_cska22_fa19_or0;
  wire [0:0] u_cska22_xor21;
  wire [0:0] u_cska22_fa20_xor1;
  wire [0:0] u_cska22_fa20_or0;
  wire [0:0] u_cska22_and_propagate515;
  wire [0:0] u_cska22_mux2to15_xor0;

  xor_gate xor_gate_u_cska22_xor0(.a(a[0]), .b(b[0]), .out(u_cska22_xor0));
  ha ha_u_cska22_ha0_out(.a(a[0]), .b(b[0]), .ha_xor0(u_cska22_ha0_xor0), .ha_and0(u_cska22_ha0_and0));
  xor_gate xor_gate_u_cska22_xor1(.a(a[1]), .b(b[1]), .out(u_cska22_xor1));
  fa fa_u_cska22_fa0_out(.a(a[1]), .b(b[1]), .cin(u_cska22_ha0_and0[0]), .fa_xor1(u_cska22_fa0_xor1), .fa_or0(u_cska22_fa0_or0));
  xor_gate xor_gate_u_cska22_xor2(.a(a[2]), .b(b[2]), .out(u_cska22_xor2));
  fa fa_u_cska22_fa1_out(.a(a[2]), .b(b[2]), .cin(u_cska22_fa0_or0[0]), .fa_xor1(u_cska22_fa1_xor1), .fa_or0(u_cska22_fa1_or0));
  xor_gate xor_gate_u_cska22_xor3(.a(a[3]), .b(b[3]), .out(u_cska22_xor3));
  fa fa_u_cska22_fa2_out(.a(a[3]), .b(b[3]), .cin(u_cska22_fa1_or0[0]), .fa_xor1(u_cska22_fa2_xor1), .fa_or0(u_cska22_fa2_or0));
  and_gate and_gate_u_cska22_and_propagate00(.a(u_cska22_xor0[0]), .b(u_cska22_xor2[0]), .out(u_cska22_and_propagate00));
  and_gate and_gate_u_cska22_and_propagate01(.a(u_cska22_xor1[0]), .b(u_cska22_xor3[0]), .out(u_cska22_and_propagate01));
  and_gate and_gate_u_cska22_and_propagate02(.a(u_cska22_and_propagate00[0]), .b(u_cska22_and_propagate01[0]), .out(u_cska22_and_propagate02));
  mux2to1 mux2to1_u_cska22_mux2to10_out(.d0(u_cska22_fa2_or0[0]), .d1(1'b0), .sel(u_cska22_and_propagate02[0]), .mux2to1_xor0(u_cska22_mux2to10_and1));
  xor_gate xor_gate_u_cska22_xor4(.a(a[4]), .b(b[4]), .out(u_cska22_xor4));
  fa fa_u_cska22_fa3_out(.a(a[4]), .b(b[4]), .cin(u_cska22_mux2to10_and1[0]), .fa_xor1(u_cska22_fa3_xor1), .fa_or0(u_cska22_fa3_or0));
  xor_gate xor_gate_u_cska22_xor5(.a(a[5]), .b(b[5]), .out(u_cska22_xor5));
  fa fa_u_cska22_fa4_out(.a(a[5]), .b(b[5]), .cin(u_cska22_fa3_or0[0]), .fa_xor1(u_cska22_fa4_xor1), .fa_or0(u_cska22_fa4_or0));
  xor_gate xor_gate_u_cska22_xor6(.a(a[6]), .b(b[6]), .out(u_cska22_xor6));
  fa fa_u_cska22_fa5_out(.a(a[6]), .b(b[6]), .cin(u_cska22_fa4_or0[0]), .fa_xor1(u_cska22_fa5_xor1), .fa_or0(u_cska22_fa5_or0));
  xor_gate xor_gate_u_cska22_xor7(.a(a[7]), .b(b[7]), .out(u_cska22_xor7));
  fa fa_u_cska22_fa6_out(.a(a[7]), .b(b[7]), .cin(u_cska22_fa5_or0[0]), .fa_xor1(u_cska22_fa6_xor1), .fa_or0(u_cska22_fa6_or0));
  and_gate and_gate_u_cska22_and_propagate13(.a(u_cska22_xor4[0]), .b(u_cska22_xor6[0]), .out(u_cska22_and_propagate13));
  and_gate and_gate_u_cska22_and_propagate14(.a(u_cska22_xor5[0]), .b(u_cska22_xor7[0]), .out(u_cska22_and_propagate14));
  and_gate and_gate_u_cska22_and_propagate15(.a(u_cska22_and_propagate13[0]), .b(u_cska22_and_propagate14[0]), .out(u_cska22_and_propagate15));
  mux2to1 mux2to1_u_cska22_mux2to11_out(.d0(u_cska22_fa6_or0[0]), .d1(u_cska22_mux2to10_and1[0]), .sel(u_cska22_and_propagate15[0]), .mux2to1_xor0(u_cska22_mux2to11_xor0));
  xor_gate xor_gate_u_cska22_xor8(.a(a[8]), .b(b[8]), .out(u_cska22_xor8));
  fa fa_u_cska22_fa7_out(.a(a[8]), .b(b[8]), .cin(u_cska22_mux2to11_xor0[0]), .fa_xor1(u_cska22_fa7_xor1), .fa_or0(u_cska22_fa7_or0));
  xor_gate xor_gate_u_cska22_xor9(.a(a[9]), .b(b[9]), .out(u_cska22_xor9));
  fa fa_u_cska22_fa8_out(.a(a[9]), .b(b[9]), .cin(u_cska22_fa7_or0[0]), .fa_xor1(u_cska22_fa8_xor1), .fa_or0(u_cska22_fa8_or0));
  xor_gate xor_gate_u_cska22_xor10(.a(a[10]), .b(b[10]), .out(u_cska22_xor10));
  fa fa_u_cska22_fa9_out(.a(a[10]), .b(b[10]), .cin(u_cska22_fa8_or0[0]), .fa_xor1(u_cska22_fa9_xor1), .fa_or0(u_cska22_fa9_or0));
  xor_gate xor_gate_u_cska22_xor11(.a(a[11]), .b(b[11]), .out(u_cska22_xor11));
  fa fa_u_cska22_fa10_out(.a(a[11]), .b(b[11]), .cin(u_cska22_fa9_or0[0]), .fa_xor1(u_cska22_fa10_xor1), .fa_or0(u_cska22_fa10_or0));
  and_gate and_gate_u_cska22_and_propagate26(.a(u_cska22_xor8[0]), .b(u_cska22_xor10[0]), .out(u_cska22_and_propagate26));
  and_gate and_gate_u_cska22_and_propagate27(.a(u_cska22_xor9[0]), .b(u_cska22_xor11[0]), .out(u_cska22_and_propagate27));
  and_gate and_gate_u_cska22_and_propagate28(.a(u_cska22_and_propagate26[0]), .b(u_cska22_and_propagate27[0]), .out(u_cska22_and_propagate28));
  mux2to1 mux2to1_u_cska22_mux2to12_out(.d0(u_cska22_fa10_or0[0]), .d1(u_cska22_mux2to11_xor0[0]), .sel(u_cska22_and_propagate28[0]), .mux2to1_xor0(u_cska22_mux2to12_xor0));
  xor_gate xor_gate_u_cska22_xor12(.a(a[12]), .b(b[12]), .out(u_cska22_xor12));
  fa fa_u_cska22_fa11_out(.a(a[12]), .b(b[12]), .cin(u_cska22_mux2to12_xor0[0]), .fa_xor1(u_cska22_fa11_xor1), .fa_or0(u_cska22_fa11_or0));
  xor_gate xor_gate_u_cska22_xor13(.a(a[13]), .b(b[13]), .out(u_cska22_xor13));
  fa fa_u_cska22_fa12_out(.a(a[13]), .b(b[13]), .cin(u_cska22_fa11_or0[0]), .fa_xor1(u_cska22_fa12_xor1), .fa_or0(u_cska22_fa12_or0));
  xor_gate xor_gate_u_cska22_xor14(.a(a[14]), .b(b[14]), .out(u_cska22_xor14));
  fa fa_u_cska22_fa13_out(.a(a[14]), .b(b[14]), .cin(u_cska22_fa12_or0[0]), .fa_xor1(u_cska22_fa13_xor1), .fa_or0(u_cska22_fa13_or0));
  xor_gate xor_gate_u_cska22_xor15(.a(a[15]), .b(b[15]), .out(u_cska22_xor15));
  fa fa_u_cska22_fa14_out(.a(a[15]), .b(b[15]), .cin(u_cska22_fa13_or0[0]), .fa_xor1(u_cska22_fa14_xor1), .fa_or0(u_cska22_fa14_or0));
  and_gate and_gate_u_cska22_and_propagate39(.a(u_cska22_xor12[0]), .b(u_cska22_xor14[0]), .out(u_cska22_and_propagate39));
  and_gate and_gate_u_cska22_and_propagate310(.a(u_cska22_xor13[0]), .b(u_cska22_xor15[0]), .out(u_cska22_and_propagate310));
  and_gate and_gate_u_cska22_and_propagate311(.a(u_cska22_and_propagate39[0]), .b(u_cska22_and_propagate310[0]), .out(u_cska22_and_propagate311));
  mux2to1 mux2to1_u_cska22_mux2to13_out(.d0(u_cska22_fa14_or0[0]), .d1(u_cska22_mux2to12_xor0[0]), .sel(u_cska22_and_propagate311[0]), .mux2to1_xor0(u_cska22_mux2to13_xor0));
  xor_gate xor_gate_u_cska22_xor16(.a(a[16]), .b(b[16]), .out(u_cska22_xor16));
  fa fa_u_cska22_fa15_out(.a(a[16]), .b(b[16]), .cin(u_cska22_mux2to13_xor0[0]), .fa_xor1(u_cska22_fa15_xor1), .fa_or0(u_cska22_fa15_or0));
  xor_gate xor_gate_u_cska22_xor17(.a(a[17]), .b(b[17]), .out(u_cska22_xor17));
  fa fa_u_cska22_fa16_out(.a(a[17]), .b(b[17]), .cin(u_cska22_fa15_or0[0]), .fa_xor1(u_cska22_fa16_xor1), .fa_or0(u_cska22_fa16_or0));
  xor_gate xor_gate_u_cska22_xor18(.a(a[18]), .b(b[18]), .out(u_cska22_xor18));
  fa fa_u_cska22_fa17_out(.a(a[18]), .b(b[18]), .cin(u_cska22_fa16_or0[0]), .fa_xor1(u_cska22_fa17_xor1), .fa_or0(u_cska22_fa17_or0));
  xor_gate xor_gate_u_cska22_xor19(.a(a[19]), .b(b[19]), .out(u_cska22_xor19));
  fa fa_u_cska22_fa18_out(.a(a[19]), .b(b[19]), .cin(u_cska22_fa17_or0[0]), .fa_xor1(u_cska22_fa18_xor1), .fa_or0(u_cska22_fa18_or0));
  and_gate and_gate_u_cska22_and_propagate412(.a(u_cska22_xor16[0]), .b(u_cska22_xor18[0]), .out(u_cska22_and_propagate412));
  and_gate and_gate_u_cska22_and_propagate413(.a(u_cska22_xor17[0]), .b(u_cska22_xor19[0]), .out(u_cska22_and_propagate413));
  and_gate and_gate_u_cska22_and_propagate414(.a(u_cska22_and_propagate412[0]), .b(u_cska22_and_propagate413[0]), .out(u_cska22_and_propagate414));
  mux2to1 mux2to1_u_cska22_mux2to14_out(.d0(u_cska22_fa18_or0[0]), .d1(u_cska22_mux2to13_xor0[0]), .sel(u_cska22_and_propagate414[0]), .mux2to1_xor0(u_cska22_mux2to14_xor0));
  xor_gate xor_gate_u_cska22_xor20(.a(a[20]), .b(b[20]), .out(u_cska22_xor20));
  fa fa_u_cska22_fa19_out(.a(a[20]), .b(b[20]), .cin(u_cska22_mux2to14_xor0[0]), .fa_xor1(u_cska22_fa19_xor1), .fa_or0(u_cska22_fa19_or0));
  xor_gate xor_gate_u_cska22_xor21(.a(a[21]), .b(b[21]), .out(u_cska22_xor21));
  fa fa_u_cska22_fa20_out(.a(a[21]), .b(b[21]), .cin(u_cska22_fa19_or0[0]), .fa_xor1(u_cska22_fa20_xor1), .fa_or0(u_cska22_fa20_or0));
  and_gate and_gate_u_cska22_and_propagate515(.a(u_cska22_xor20[0]), .b(u_cska22_xor21[0]), .out(u_cska22_and_propagate515));
  mux2to1 mux2to1_u_cska22_mux2to15_out(.d0(u_cska22_fa20_or0[0]), .d1(u_cska22_mux2to14_xor0[0]), .sel(u_cska22_and_propagate515[0]), .mux2to1_xor0(u_cska22_mux2to15_xor0));

  assign u_cska22_out[0] = u_cska22_ha0_xor0[0];
  assign u_cska22_out[1] = u_cska22_fa0_xor1[0];
  assign u_cska22_out[2] = u_cska22_fa1_xor1[0];
  assign u_cska22_out[3] = u_cska22_fa2_xor1[0];
  assign u_cska22_out[4] = u_cska22_fa3_xor1[0];
  assign u_cska22_out[5] = u_cska22_fa4_xor1[0];
  assign u_cska22_out[6] = u_cska22_fa5_xor1[0];
  assign u_cska22_out[7] = u_cska22_fa6_xor1[0];
  assign u_cska22_out[8] = u_cska22_fa7_xor1[0];
  assign u_cska22_out[9] = u_cska22_fa8_xor1[0];
  assign u_cska22_out[10] = u_cska22_fa9_xor1[0];
  assign u_cska22_out[11] = u_cska22_fa10_xor1[0];
  assign u_cska22_out[12] = u_cska22_fa11_xor1[0];
  assign u_cska22_out[13] = u_cska22_fa12_xor1[0];
  assign u_cska22_out[14] = u_cska22_fa13_xor1[0];
  assign u_cska22_out[15] = u_cska22_fa14_xor1[0];
  assign u_cska22_out[16] = u_cska22_fa15_xor1[0];
  assign u_cska22_out[17] = u_cska22_fa16_xor1[0];
  assign u_cska22_out[18] = u_cska22_fa17_xor1[0];
  assign u_cska22_out[19] = u_cska22_fa18_xor1[0];
  assign u_cska22_out[20] = u_cska22_fa19_xor1[0];
  assign u_cska22_out[21] = u_cska22_fa20_xor1[0];
  assign u_cska22_out[22] = u_cska22_mux2to15_xor0[0];
endmodule

module s_dadda_cska12(input [11:0] a, input [11:0] b, output [23:0] s_dadda_cska12_out);
  wire [0:0] s_dadda_cska12_and_9_0;
  wire [0:0] s_dadda_cska12_and_8_1;
  wire [0:0] s_dadda_cska12_ha0_xor0;
  wire [0:0] s_dadda_cska12_ha0_and0;
  wire [0:0] s_dadda_cska12_and_10_0;
  wire [0:0] s_dadda_cska12_and_9_1;
  wire [0:0] s_dadda_cska12_fa0_xor1;
  wire [0:0] s_dadda_cska12_fa0_or0;
  wire [0:0] s_dadda_cska12_and_8_2;
  wire [0:0] s_dadda_cska12_and_7_3;
  wire [0:0] s_dadda_cska12_ha1_xor0;
  wire [0:0] s_dadda_cska12_ha1_and0;
  wire [0:0] s_dadda_cska12_nand_11_0;
  wire [0:0] s_dadda_cska12_fa1_xor1;
  wire [0:0] s_dadda_cska12_fa1_or0;
  wire [0:0] s_dadda_cska12_and_10_1;
  wire [0:0] s_dadda_cska12_and_9_2;
  wire [0:0] s_dadda_cska12_and_8_3;
  wire [0:0] s_dadda_cska12_fa2_xor1;
  wire [0:0] s_dadda_cska12_fa2_or0;
  wire [0:0] s_dadda_cska12_and_7_4;
  wire [0:0] s_dadda_cska12_and_6_5;
  wire [0:0] s_dadda_cska12_ha2_xor0;
  wire [0:0] s_dadda_cska12_ha2_and0;
  wire [0:0] s_dadda_cska12_fa3_xor1;
  wire [0:0] s_dadda_cska12_fa3_or0;
  wire [0:0] s_dadda_cska12_nand_11_1;
  wire [0:0] s_dadda_cska12_and_10_2;
  wire [0:0] s_dadda_cska12_fa4_xor1;
  wire [0:0] s_dadda_cska12_fa4_or0;
  wire [0:0] s_dadda_cska12_and_9_3;
  wire [0:0] s_dadda_cska12_and_8_4;
  wire [0:0] s_dadda_cska12_and_7_5;
  wire [0:0] s_dadda_cska12_fa5_xor1;
  wire [0:0] s_dadda_cska12_fa5_or0;
  wire [0:0] s_dadda_cska12_fa6_xor1;
  wire [0:0] s_dadda_cska12_fa6_or0;
  wire [0:0] s_dadda_cska12_nand_11_2;
  wire [0:0] s_dadda_cska12_and_10_3;
  wire [0:0] s_dadda_cska12_and_9_4;
  wire [0:0] s_dadda_cska12_fa7_xor1;
  wire [0:0] s_dadda_cska12_fa7_or0;
  wire [0:0] s_dadda_cska12_nand_11_3;
  wire [0:0] s_dadda_cska12_fa8_xor1;
  wire [0:0] s_dadda_cska12_fa8_or0;
  wire [0:0] s_dadda_cska12_and_4_0;
  wire [0:0] s_dadda_cska12_and_3_1;
  wire [0:0] s_dadda_cska12_ha3_xor0;
  wire [0:0] s_dadda_cska12_ha3_and0;
  wire [0:0] s_dadda_cska12_and_5_0;
  wire [0:0] s_dadda_cska12_and_4_1;
  wire [0:0] s_dadda_cska12_fa9_xor1;
  wire [0:0] s_dadda_cska12_fa9_or0;
  wire [0:0] s_dadda_cska12_and_3_2;
  wire [0:0] s_dadda_cska12_and_2_3;
  wire [0:0] s_dadda_cska12_ha4_xor0;
  wire [0:0] s_dadda_cska12_ha4_and0;
  wire [0:0] s_dadda_cska12_and_6_0;
  wire [0:0] s_dadda_cska12_fa10_xor1;
  wire [0:0] s_dadda_cska12_fa10_or0;
  wire [0:0] s_dadda_cska12_and_5_1;
  wire [0:0] s_dadda_cska12_and_4_2;
  wire [0:0] s_dadda_cska12_and_3_3;
  wire [0:0] s_dadda_cska12_fa11_xor1;
  wire [0:0] s_dadda_cska12_fa11_or0;
  wire [0:0] s_dadda_cska12_and_2_4;
  wire [0:0] s_dadda_cska12_and_1_5;
  wire [0:0] s_dadda_cska12_ha5_xor0;
  wire [0:0] s_dadda_cska12_ha5_and0;
  wire [0:0] s_dadda_cska12_fa12_xor1;
  wire [0:0] s_dadda_cska12_fa12_or0;
  wire [0:0] s_dadda_cska12_and_7_0;
  wire [0:0] s_dadda_cska12_and_6_1;
  wire [0:0] s_dadda_cska12_and_5_2;
  wire [0:0] s_dadda_cska12_fa13_xor1;
  wire [0:0] s_dadda_cska12_fa13_or0;
  wire [0:0] s_dadda_cska12_and_4_3;
  wire [0:0] s_dadda_cska12_and_3_4;
  wire [0:0] s_dadda_cska12_and_2_5;
  wire [0:0] s_dadda_cska12_fa14_xor1;
  wire [0:0] s_dadda_cska12_fa14_or0;
  wire [0:0] s_dadda_cska12_and_1_6;
  wire [0:0] s_dadda_cska12_and_0_7;
  wire [0:0] s_dadda_cska12_ha6_xor0;
  wire [0:0] s_dadda_cska12_ha6_and0;
  wire [0:0] s_dadda_cska12_fa15_xor1;
  wire [0:0] s_dadda_cska12_fa15_or0;
  wire [0:0] s_dadda_cska12_and_8_0;
  wire [0:0] s_dadda_cska12_and_7_1;
  wire [0:0] s_dadda_cska12_fa16_xor1;
  wire [0:0] s_dadda_cska12_fa16_or0;
  wire [0:0] s_dadda_cska12_and_6_2;
  wire [0:0] s_dadda_cska12_and_5_3;
  wire [0:0] s_dadda_cska12_and_4_4;
  wire [0:0] s_dadda_cska12_fa17_xor1;
  wire [0:0] s_dadda_cska12_fa17_or0;
  wire [0:0] s_dadda_cska12_and_3_5;
  wire [0:0] s_dadda_cska12_and_2_6;
  wire [0:0] s_dadda_cska12_and_1_7;
  wire [0:0] s_dadda_cska12_fa18_xor1;
  wire [0:0] s_dadda_cska12_fa18_or0;
  wire [0:0] s_dadda_cska12_and_0_8;
  wire [0:0] s_dadda_cska12_ha7_xor0;
  wire [0:0] s_dadda_cska12_ha7_and0;
  wire [0:0] s_dadda_cska12_fa19_xor1;
  wire [0:0] s_dadda_cska12_fa19_or0;
  wire [0:0] s_dadda_cska12_and_7_2;
  wire [0:0] s_dadda_cska12_fa20_xor1;
  wire [0:0] s_dadda_cska12_fa20_or0;
  wire [0:0] s_dadda_cska12_and_6_3;
  wire [0:0] s_dadda_cska12_and_5_4;
  wire [0:0] s_dadda_cska12_and_4_5;
  wire [0:0] s_dadda_cska12_fa21_xor1;
  wire [0:0] s_dadda_cska12_fa21_or0;
  wire [0:0] s_dadda_cska12_and_3_6;
  wire [0:0] s_dadda_cska12_and_2_7;
  wire [0:0] s_dadda_cska12_and_1_8;
  wire [0:0] s_dadda_cska12_fa22_xor1;
  wire [0:0] s_dadda_cska12_fa22_or0;
  wire [0:0] s_dadda_cska12_and_0_9;
  wire [0:0] s_dadda_cska12_fa23_xor1;
  wire [0:0] s_dadda_cska12_fa23_or0;
  wire [0:0] s_dadda_cska12_fa24_xor1;
  wire [0:0] s_dadda_cska12_fa24_or0;
  wire [0:0] s_dadda_cska12_and_6_4;
  wire [0:0] s_dadda_cska12_fa25_xor1;
  wire [0:0] s_dadda_cska12_fa25_or0;
  wire [0:0] s_dadda_cska12_and_5_5;
  wire [0:0] s_dadda_cska12_and_4_6;
  wire [0:0] s_dadda_cska12_and_3_7;
  wire [0:0] s_dadda_cska12_fa26_xor1;
  wire [0:0] s_dadda_cska12_fa26_or0;
  wire [0:0] s_dadda_cska12_and_2_8;
  wire [0:0] s_dadda_cska12_and_1_9;
  wire [0:0] s_dadda_cska12_and_0_10;
  wire [0:0] s_dadda_cska12_fa27_xor1;
  wire [0:0] s_dadda_cska12_fa27_or0;
  wire [0:0] s_dadda_cska12_fa28_xor1;
  wire [0:0] s_dadda_cska12_fa28_or0;
  wire [0:0] s_dadda_cska12_fa29_xor1;
  wire [0:0] s_dadda_cska12_fa29_or0;
  wire [0:0] s_dadda_cska12_and_5_6;
  wire [0:0] s_dadda_cska12_fa30_xor1;
  wire [0:0] s_dadda_cska12_fa30_or0;
  wire [0:0] s_dadda_cska12_and_4_7;
  wire [0:0] s_dadda_cska12_and_3_8;
  wire [0:0] s_dadda_cska12_and_2_9;
  wire [0:0] s_dadda_cska12_fa31_xor1;
  wire [0:0] s_dadda_cska12_fa31_or0;
  wire [0:0] s_dadda_cska12_and_1_10;
  wire [0:0] s_dadda_cska12_nand_0_11;
  wire [0:0] s_dadda_cska12_fa32_xor1;
  wire [0:0] s_dadda_cska12_fa32_or0;
  wire [0:0] s_dadda_cska12_fa33_xor1;
  wire [0:0] s_dadda_cska12_fa33_or0;
  wire [0:0] s_dadda_cska12_fa34_xor1;
  wire [0:0] s_dadda_cska12_fa34_or0;
  wire [0:0] s_dadda_cska12_and_6_6;
  wire [0:0] s_dadda_cska12_fa35_xor1;
  wire [0:0] s_dadda_cska12_fa35_or0;
  wire [0:0] s_dadda_cska12_and_5_7;
  wire [0:0] s_dadda_cska12_and_4_8;
  wire [0:0] s_dadda_cska12_and_3_9;
  wire [0:0] s_dadda_cska12_fa36_xor1;
  wire [0:0] s_dadda_cska12_fa36_or0;
  wire [0:0] s_dadda_cska12_and_2_10;
  wire [0:0] s_dadda_cska12_nand_1_11;
  wire [0:0] s_dadda_cska12_fa37_xor1;
  wire [0:0] s_dadda_cska12_fa37_or0;
  wire [0:0] s_dadda_cska12_fa38_xor1;
  wire [0:0] s_dadda_cska12_fa38_or0;
  wire [0:0] s_dadda_cska12_fa39_xor1;
  wire [0:0] s_dadda_cska12_fa39_or0;
  wire [0:0] s_dadda_cska12_and_8_5;
  wire [0:0] s_dadda_cska12_fa40_xor1;
  wire [0:0] s_dadda_cska12_fa40_or0;
  wire [0:0] s_dadda_cska12_and_7_6;
  wire [0:0] s_dadda_cska12_and_6_7;
  wire [0:0] s_dadda_cska12_and_5_8;
  wire [0:0] s_dadda_cska12_fa41_xor1;
  wire [0:0] s_dadda_cska12_fa41_or0;
  wire [0:0] s_dadda_cska12_and_4_9;
  wire [0:0] s_dadda_cska12_and_3_10;
  wire [0:0] s_dadda_cska12_nand_2_11;
  wire [0:0] s_dadda_cska12_fa42_xor1;
  wire [0:0] s_dadda_cska12_fa42_or0;
  wire [0:0] s_dadda_cska12_fa43_xor1;
  wire [0:0] s_dadda_cska12_fa43_or0;
  wire [0:0] s_dadda_cska12_fa44_xor1;
  wire [0:0] s_dadda_cska12_fa44_or0;
  wire [0:0] s_dadda_cska12_and_10_4;
  wire [0:0] s_dadda_cska12_fa45_xor1;
  wire [0:0] s_dadda_cska12_fa45_or0;
  wire [0:0] s_dadda_cska12_and_9_5;
  wire [0:0] s_dadda_cska12_and_8_6;
  wire [0:0] s_dadda_cska12_and_7_7;
  wire [0:0] s_dadda_cska12_fa46_xor1;
  wire [0:0] s_dadda_cska12_fa46_or0;
  wire [0:0] s_dadda_cska12_and_6_8;
  wire [0:0] s_dadda_cska12_and_5_9;
  wire [0:0] s_dadda_cska12_and_4_10;
  wire [0:0] s_dadda_cska12_fa47_xor1;
  wire [0:0] s_dadda_cska12_fa47_or0;
  wire [0:0] s_dadda_cska12_nand_3_11;
  wire [0:0] s_dadda_cska12_fa48_xor1;
  wire [0:0] s_dadda_cska12_fa48_or0;
  wire [0:0] s_dadda_cska12_fa49_xor1;
  wire [0:0] s_dadda_cska12_fa49_or0;
  wire [0:0] s_dadda_cska12_fa50_xor1;
  wire [0:0] s_dadda_cska12_fa50_or0;
  wire [0:0] s_dadda_cska12_nand_11_4;
  wire [0:0] s_dadda_cska12_and_10_5;
  wire [0:0] s_dadda_cska12_and_9_6;
  wire [0:0] s_dadda_cska12_fa51_xor1;
  wire [0:0] s_dadda_cska12_fa51_or0;
  wire [0:0] s_dadda_cska12_and_8_7;
  wire [0:0] s_dadda_cska12_and_7_8;
  wire [0:0] s_dadda_cska12_and_6_9;
  wire [0:0] s_dadda_cska12_fa52_xor1;
  wire [0:0] s_dadda_cska12_fa52_or0;
  wire [0:0] s_dadda_cska12_and_5_10;
  wire [0:0] s_dadda_cska12_nand_4_11;
  wire [0:0] s_dadda_cska12_fa53_xor1;
  wire [0:0] s_dadda_cska12_fa53_or0;
  wire [0:0] s_dadda_cska12_fa54_xor1;
  wire [0:0] s_dadda_cska12_fa54_or0;
  wire [0:0] s_dadda_cska12_nand_11_5;
  wire [0:0] s_dadda_cska12_fa55_xor1;
  wire [0:0] s_dadda_cska12_fa55_or0;
  wire [0:0] s_dadda_cska12_and_10_6;
  wire [0:0] s_dadda_cska12_and_9_7;
  wire [0:0] s_dadda_cska12_and_8_8;
  wire [0:0] s_dadda_cska12_fa56_xor1;
  wire [0:0] s_dadda_cska12_fa56_or0;
  wire [0:0] s_dadda_cska12_and_7_9;
  wire [0:0] s_dadda_cska12_and_6_10;
  wire [0:0] s_dadda_cska12_nand_5_11;
  wire [0:0] s_dadda_cska12_fa57_xor1;
  wire [0:0] s_dadda_cska12_fa57_or0;
  wire [0:0] s_dadda_cska12_fa58_xor1;
  wire [0:0] s_dadda_cska12_fa58_or0;
  wire [0:0] s_dadda_cska12_nand_11_6;
  wire [0:0] s_dadda_cska12_and_10_7;
  wire [0:0] s_dadda_cska12_fa59_xor1;
  wire [0:0] s_dadda_cska12_fa59_or0;
  wire [0:0] s_dadda_cska12_and_9_8;
  wire [0:0] s_dadda_cska12_and_8_9;
  wire [0:0] s_dadda_cska12_and_7_10;
  wire [0:0] s_dadda_cska12_fa60_xor1;
  wire [0:0] s_dadda_cska12_fa60_or0;
  wire [0:0] s_dadda_cska12_fa61_xor1;
  wire [0:0] s_dadda_cska12_fa61_or0;
  wire [0:0] s_dadda_cska12_nand_11_7;
  wire [0:0] s_dadda_cska12_and_10_8;
  wire [0:0] s_dadda_cska12_and_9_9;
  wire [0:0] s_dadda_cska12_fa62_xor1;
  wire [0:0] s_dadda_cska12_fa62_or0;
  wire [0:0] s_dadda_cska12_nand_11_8;
  wire [0:0] s_dadda_cska12_fa63_xor1;
  wire [0:0] s_dadda_cska12_fa63_or0;
  wire [0:0] s_dadda_cska12_and_3_0;
  wire [0:0] s_dadda_cska12_and_2_1;
  wire [0:0] s_dadda_cska12_ha8_xor0;
  wire [0:0] s_dadda_cska12_ha8_and0;
  wire [0:0] s_dadda_cska12_and_2_2;
  wire [0:0] s_dadda_cska12_and_1_3;
  wire [0:0] s_dadda_cska12_fa64_xor1;
  wire [0:0] s_dadda_cska12_fa64_or0;
  wire [0:0] s_dadda_cska12_and_1_4;
  wire [0:0] s_dadda_cska12_and_0_5;
  wire [0:0] s_dadda_cska12_fa65_xor1;
  wire [0:0] s_dadda_cska12_fa65_or0;
  wire [0:0] s_dadda_cska12_and_0_6;
  wire [0:0] s_dadda_cska12_fa66_xor1;
  wire [0:0] s_dadda_cska12_fa66_or0;
  wire [0:0] s_dadda_cska12_fa67_xor1;
  wire [0:0] s_dadda_cska12_fa67_or0;
  wire [0:0] s_dadda_cska12_fa68_xor1;
  wire [0:0] s_dadda_cska12_fa68_or0;
  wire [0:0] s_dadda_cska12_fa69_xor1;
  wire [0:0] s_dadda_cska12_fa69_or0;
  wire [0:0] s_dadda_cska12_fa70_xor1;
  wire [0:0] s_dadda_cska12_fa70_or0;
  wire [0:0] s_dadda_cska12_fa71_xor1;
  wire [0:0] s_dadda_cska12_fa71_or0;
  wire [0:0] s_dadda_cska12_fa72_xor1;
  wire [0:0] s_dadda_cska12_fa72_or0;
  wire [0:0] s_dadda_cska12_fa73_xor1;
  wire [0:0] s_dadda_cska12_fa73_or0;
  wire [0:0] s_dadda_cska12_fa74_xor1;
  wire [0:0] s_dadda_cska12_fa74_or0;
  wire [0:0] s_dadda_cska12_fa75_xor1;
  wire [0:0] s_dadda_cska12_fa75_or0;
  wire [0:0] s_dadda_cska12_fa76_xor1;
  wire [0:0] s_dadda_cska12_fa76_or0;
  wire [0:0] s_dadda_cska12_nand_6_11;
  wire [0:0] s_dadda_cska12_fa77_xor1;
  wire [0:0] s_dadda_cska12_fa77_or0;
  wire [0:0] s_dadda_cska12_and_8_10;
  wire [0:0] s_dadda_cska12_nand_7_11;
  wire [0:0] s_dadda_cska12_fa78_xor1;
  wire [0:0] s_dadda_cska12_fa78_or0;
  wire [0:0] s_dadda_cska12_and_10_9;
  wire [0:0] s_dadda_cska12_and_9_10;
  wire [0:0] s_dadda_cska12_fa79_xor1;
  wire [0:0] s_dadda_cska12_fa79_or0;
  wire [0:0] s_dadda_cska12_nand_11_9;
  wire [0:0] s_dadda_cska12_fa80_xor1;
  wire [0:0] s_dadda_cska12_fa80_or0;
  wire [0:0] s_dadda_cska12_and_2_0;
  wire [0:0] s_dadda_cska12_and_1_1;
  wire [0:0] s_dadda_cska12_ha9_xor0;
  wire [0:0] s_dadda_cska12_ha9_and0;
  wire [0:0] s_dadda_cska12_and_1_2;
  wire [0:0] s_dadda_cska12_and_0_3;
  wire [0:0] s_dadda_cska12_fa81_xor1;
  wire [0:0] s_dadda_cska12_fa81_or0;
  wire [0:0] s_dadda_cska12_and_0_4;
  wire [0:0] s_dadda_cska12_fa82_xor1;
  wire [0:0] s_dadda_cska12_fa82_or0;
  wire [0:0] s_dadda_cska12_fa83_xor1;
  wire [0:0] s_dadda_cska12_fa83_or0;
  wire [0:0] s_dadda_cska12_fa84_xor1;
  wire [0:0] s_dadda_cska12_fa84_or0;
  wire [0:0] s_dadda_cska12_fa85_xor1;
  wire [0:0] s_dadda_cska12_fa85_or0;
  wire [0:0] s_dadda_cska12_fa86_xor1;
  wire [0:0] s_dadda_cska12_fa86_or0;
  wire [0:0] s_dadda_cska12_fa87_xor1;
  wire [0:0] s_dadda_cska12_fa87_or0;
  wire [0:0] s_dadda_cska12_fa88_xor1;
  wire [0:0] s_dadda_cska12_fa88_or0;
  wire [0:0] s_dadda_cska12_fa89_xor1;
  wire [0:0] s_dadda_cska12_fa89_or0;
  wire [0:0] s_dadda_cska12_fa90_xor1;
  wire [0:0] s_dadda_cska12_fa90_or0;
  wire [0:0] s_dadda_cska12_fa91_xor1;
  wire [0:0] s_dadda_cska12_fa91_or0;
  wire [0:0] s_dadda_cska12_fa92_xor1;
  wire [0:0] s_dadda_cska12_fa92_or0;
  wire [0:0] s_dadda_cska12_fa93_xor1;
  wire [0:0] s_dadda_cska12_fa93_or0;
  wire [0:0] s_dadda_cska12_fa94_xor1;
  wire [0:0] s_dadda_cska12_fa94_or0;
  wire [0:0] s_dadda_cska12_fa95_xor1;
  wire [0:0] s_dadda_cska12_fa95_or0;
  wire [0:0] s_dadda_cska12_fa96_xor1;
  wire [0:0] s_dadda_cska12_fa96_or0;
  wire [0:0] s_dadda_cska12_nand_8_11;
  wire [0:0] s_dadda_cska12_fa97_xor1;
  wire [0:0] s_dadda_cska12_fa97_or0;
  wire [0:0] s_dadda_cska12_and_10_10;
  wire [0:0] s_dadda_cska12_nand_9_11;
  wire [0:0] s_dadda_cska12_fa98_xor1;
  wire [0:0] s_dadda_cska12_fa98_or0;
  wire [0:0] s_dadda_cska12_nand_11_10;
  wire [0:0] s_dadda_cska12_fa99_xor1;
  wire [0:0] s_dadda_cska12_fa99_or0;
  wire [0:0] s_dadda_cska12_and_0_0;
  wire [0:0] s_dadda_cska12_and_1_0;
  wire [0:0] s_dadda_cska12_and_0_2;
  wire [0:0] s_dadda_cska12_nand_10_11;
  wire [0:0] s_dadda_cska12_and_0_1;
  wire [0:0] s_dadda_cska12_and_11_11;
  wire [21:0] s_dadda_cska12_u_cska22_a;
  wire [21:0] s_dadda_cska12_u_cska22_b;
  wire [22:0] s_dadda_cska12_u_cska22_out;
  wire [0:0] s_dadda_cska12_xor0;

  and_gate and_gate_s_dadda_cska12_and_9_0(.a(a[9]), .b(b[0]), .out(s_dadda_cska12_and_9_0));
  and_gate and_gate_s_dadda_cska12_and_8_1(.a(a[8]), .b(b[1]), .out(s_dadda_cska12_and_8_1));
  ha ha_s_dadda_cska12_ha0_out(.a(s_dadda_cska12_and_9_0[0]), .b(s_dadda_cska12_and_8_1[0]), .ha_xor0(s_dadda_cska12_ha0_xor0), .ha_and0(s_dadda_cska12_ha0_and0));
  and_gate and_gate_s_dadda_cska12_and_10_0(.a(a[10]), .b(b[0]), .out(s_dadda_cska12_and_10_0));
  and_gate and_gate_s_dadda_cska12_and_9_1(.a(a[9]), .b(b[1]), .out(s_dadda_cska12_and_9_1));
  fa fa_s_dadda_cska12_fa0_out(.a(s_dadda_cska12_ha0_and0[0]), .b(s_dadda_cska12_and_10_0[0]), .cin(s_dadda_cska12_and_9_1[0]), .fa_xor1(s_dadda_cska12_fa0_xor1), .fa_or0(s_dadda_cska12_fa0_or0));
  and_gate and_gate_s_dadda_cska12_and_8_2(.a(a[8]), .b(b[2]), .out(s_dadda_cska12_and_8_2));
  and_gate and_gate_s_dadda_cska12_and_7_3(.a(a[7]), .b(b[3]), .out(s_dadda_cska12_and_7_3));
  ha ha_s_dadda_cska12_ha1_out(.a(s_dadda_cska12_and_8_2[0]), .b(s_dadda_cska12_and_7_3[0]), .ha_xor0(s_dadda_cska12_ha1_xor0), .ha_and0(s_dadda_cska12_ha1_and0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_0(.a(a[11]), .b(b[0]), .out(s_dadda_cska12_nand_11_0));
  fa fa_s_dadda_cska12_fa1_out(.a(s_dadda_cska12_ha1_and0[0]), .b(s_dadda_cska12_fa0_or0[0]), .cin(s_dadda_cska12_nand_11_0[0]), .fa_xor1(s_dadda_cska12_fa1_xor1), .fa_or0(s_dadda_cska12_fa1_or0));
  and_gate and_gate_s_dadda_cska12_and_10_1(.a(a[10]), .b(b[1]), .out(s_dadda_cska12_and_10_1));
  and_gate and_gate_s_dadda_cska12_and_9_2(.a(a[9]), .b(b[2]), .out(s_dadda_cska12_and_9_2));
  and_gate and_gate_s_dadda_cska12_and_8_3(.a(a[8]), .b(b[3]), .out(s_dadda_cska12_and_8_3));
  fa fa_s_dadda_cska12_fa2_out(.a(s_dadda_cska12_and_10_1[0]), .b(s_dadda_cska12_and_9_2[0]), .cin(s_dadda_cska12_and_8_3[0]), .fa_xor1(s_dadda_cska12_fa2_xor1), .fa_or0(s_dadda_cska12_fa2_or0));
  and_gate and_gate_s_dadda_cska12_and_7_4(.a(a[7]), .b(b[4]), .out(s_dadda_cska12_and_7_4));
  and_gate and_gate_s_dadda_cska12_and_6_5(.a(a[6]), .b(b[5]), .out(s_dadda_cska12_and_6_5));
  ha ha_s_dadda_cska12_ha2_out(.a(s_dadda_cska12_and_7_4[0]), .b(s_dadda_cska12_and_6_5[0]), .ha_xor0(s_dadda_cska12_ha2_xor0), .ha_and0(s_dadda_cska12_ha2_and0));
  fa fa_s_dadda_cska12_fa3_out(.a(s_dadda_cska12_ha2_and0[0]), .b(s_dadda_cska12_fa2_or0[0]), .cin(s_dadda_cska12_fa1_or0[0]), .fa_xor1(s_dadda_cska12_fa3_xor1), .fa_or0(s_dadda_cska12_fa3_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_1(.a(a[11]), .b(b[1]), .out(s_dadda_cska12_nand_11_1));
  and_gate and_gate_s_dadda_cska12_and_10_2(.a(a[10]), .b(b[2]), .out(s_dadda_cska12_and_10_2));
  fa fa_s_dadda_cska12_fa4_out(.a(1'b1), .b(s_dadda_cska12_nand_11_1[0]), .cin(s_dadda_cska12_and_10_2[0]), .fa_xor1(s_dadda_cska12_fa4_xor1), .fa_or0(s_dadda_cska12_fa4_or0));
  and_gate and_gate_s_dadda_cska12_and_9_3(.a(a[9]), .b(b[3]), .out(s_dadda_cska12_and_9_3));
  and_gate and_gate_s_dadda_cska12_and_8_4(.a(a[8]), .b(b[4]), .out(s_dadda_cska12_and_8_4));
  and_gate and_gate_s_dadda_cska12_and_7_5(.a(a[7]), .b(b[5]), .out(s_dadda_cska12_and_7_5));
  fa fa_s_dadda_cska12_fa5_out(.a(s_dadda_cska12_and_9_3[0]), .b(s_dadda_cska12_and_8_4[0]), .cin(s_dadda_cska12_and_7_5[0]), .fa_xor1(s_dadda_cska12_fa5_xor1), .fa_or0(s_dadda_cska12_fa5_or0));
  fa fa_s_dadda_cska12_fa6_out(.a(s_dadda_cska12_fa5_or0[0]), .b(s_dadda_cska12_fa4_or0[0]), .cin(s_dadda_cska12_fa3_or0[0]), .fa_xor1(s_dadda_cska12_fa6_xor1), .fa_or0(s_dadda_cska12_fa6_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_2(.a(a[11]), .b(b[2]), .out(s_dadda_cska12_nand_11_2));
  and_gate and_gate_s_dadda_cska12_and_10_3(.a(a[10]), .b(b[3]), .out(s_dadda_cska12_and_10_3));
  and_gate and_gate_s_dadda_cska12_and_9_4(.a(a[9]), .b(b[4]), .out(s_dadda_cska12_and_9_4));
  fa fa_s_dadda_cska12_fa7_out(.a(s_dadda_cska12_nand_11_2[0]), .b(s_dadda_cska12_and_10_3[0]), .cin(s_dadda_cska12_and_9_4[0]), .fa_xor1(s_dadda_cska12_fa7_xor1), .fa_or0(s_dadda_cska12_fa7_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_3(.a(a[11]), .b(b[3]), .out(s_dadda_cska12_nand_11_3));
  fa fa_s_dadda_cska12_fa8_out(.a(s_dadda_cska12_fa7_or0[0]), .b(s_dadda_cska12_fa6_or0[0]), .cin(s_dadda_cska12_nand_11_3[0]), .fa_xor1(s_dadda_cska12_fa8_xor1), .fa_or0(s_dadda_cska12_fa8_or0));
  and_gate and_gate_s_dadda_cska12_and_4_0(.a(a[4]), .b(b[0]), .out(s_dadda_cska12_and_4_0));
  and_gate and_gate_s_dadda_cska12_and_3_1(.a(a[3]), .b(b[1]), .out(s_dadda_cska12_and_3_1));
  ha ha_s_dadda_cska12_ha3_out(.a(s_dadda_cska12_and_4_0[0]), .b(s_dadda_cska12_and_3_1[0]), .ha_xor0(s_dadda_cska12_ha3_xor0), .ha_and0(s_dadda_cska12_ha3_and0));
  and_gate and_gate_s_dadda_cska12_and_5_0(.a(a[5]), .b(b[0]), .out(s_dadda_cska12_and_5_0));
  and_gate and_gate_s_dadda_cska12_and_4_1(.a(a[4]), .b(b[1]), .out(s_dadda_cska12_and_4_1));
  fa fa_s_dadda_cska12_fa9_out(.a(s_dadda_cska12_ha3_and0[0]), .b(s_dadda_cska12_and_5_0[0]), .cin(s_dadda_cska12_and_4_1[0]), .fa_xor1(s_dadda_cska12_fa9_xor1), .fa_or0(s_dadda_cska12_fa9_or0));
  and_gate and_gate_s_dadda_cska12_and_3_2(.a(a[3]), .b(b[2]), .out(s_dadda_cska12_and_3_2));
  and_gate and_gate_s_dadda_cska12_and_2_3(.a(a[2]), .b(b[3]), .out(s_dadda_cska12_and_2_3));
  ha ha_s_dadda_cska12_ha4_out(.a(s_dadda_cska12_and_3_2[0]), .b(s_dadda_cska12_and_2_3[0]), .ha_xor0(s_dadda_cska12_ha4_xor0), .ha_and0(s_dadda_cska12_ha4_and0));
  and_gate and_gate_s_dadda_cska12_and_6_0(.a(a[6]), .b(b[0]), .out(s_dadda_cska12_and_6_0));
  fa fa_s_dadda_cska12_fa10_out(.a(s_dadda_cska12_ha4_and0[0]), .b(s_dadda_cska12_fa9_or0[0]), .cin(s_dadda_cska12_and_6_0[0]), .fa_xor1(s_dadda_cska12_fa10_xor1), .fa_or0(s_dadda_cska12_fa10_or0));
  and_gate and_gate_s_dadda_cska12_and_5_1(.a(a[5]), .b(b[1]), .out(s_dadda_cska12_and_5_1));
  and_gate and_gate_s_dadda_cska12_and_4_2(.a(a[4]), .b(b[2]), .out(s_dadda_cska12_and_4_2));
  and_gate and_gate_s_dadda_cska12_and_3_3(.a(a[3]), .b(b[3]), .out(s_dadda_cska12_and_3_3));
  fa fa_s_dadda_cska12_fa11_out(.a(s_dadda_cska12_and_5_1[0]), .b(s_dadda_cska12_and_4_2[0]), .cin(s_dadda_cska12_and_3_3[0]), .fa_xor1(s_dadda_cska12_fa11_xor1), .fa_or0(s_dadda_cska12_fa11_or0));
  and_gate and_gate_s_dadda_cska12_and_2_4(.a(a[2]), .b(b[4]), .out(s_dadda_cska12_and_2_4));
  and_gate and_gate_s_dadda_cska12_and_1_5(.a(a[1]), .b(b[5]), .out(s_dadda_cska12_and_1_5));
  ha ha_s_dadda_cska12_ha5_out(.a(s_dadda_cska12_and_2_4[0]), .b(s_dadda_cska12_and_1_5[0]), .ha_xor0(s_dadda_cska12_ha5_xor0), .ha_and0(s_dadda_cska12_ha5_and0));
  fa fa_s_dadda_cska12_fa12_out(.a(s_dadda_cska12_ha5_and0[0]), .b(s_dadda_cska12_fa11_or0[0]), .cin(s_dadda_cska12_fa10_or0[0]), .fa_xor1(s_dadda_cska12_fa12_xor1), .fa_or0(s_dadda_cska12_fa12_or0));
  and_gate and_gate_s_dadda_cska12_and_7_0(.a(a[7]), .b(b[0]), .out(s_dadda_cska12_and_7_0));
  and_gate and_gate_s_dadda_cska12_and_6_1(.a(a[6]), .b(b[1]), .out(s_dadda_cska12_and_6_1));
  and_gate and_gate_s_dadda_cska12_and_5_2(.a(a[5]), .b(b[2]), .out(s_dadda_cska12_and_5_2));
  fa fa_s_dadda_cska12_fa13_out(.a(s_dadda_cska12_and_7_0[0]), .b(s_dadda_cska12_and_6_1[0]), .cin(s_dadda_cska12_and_5_2[0]), .fa_xor1(s_dadda_cska12_fa13_xor1), .fa_or0(s_dadda_cska12_fa13_or0));
  and_gate and_gate_s_dadda_cska12_and_4_3(.a(a[4]), .b(b[3]), .out(s_dadda_cska12_and_4_3));
  and_gate and_gate_s_dadda_cska12_and_3_4(.a(a[3]), .b(b[4]), .out(s_dadda_cska12_and_3_4));
  and_gate and_gate_s_dadda_cska12_and_2_5(.a(a[2]), .b(b[5]), .out(s_dadda_cska12_and_2_5));
  fa fa_s_dadda_cska12_fa14_out(.a(s_dadda_cska12_and_4_3[0]), .b(s_dadda_cska12_and_3_4[0]), .cin(s_dadda_cska12_and_2_5[0]), .fa_xor1(s_dadda_cska12_fa14_xor1), .fa_or0(s_dadda_cska12_fa14_or0));
  and_gate and_gate_s_dadda_cska12_and_1_6(.a(a[1]), .b(b[6]), .out(s_dadda_cska12_and_1_6));
  and_gate and_gate_s_dadda_cska12_and_0_7(.a(a[0]), .b(b[7]), .out(s_dadda_cska12_and_0_7));
  ha ha_s_dadda_cska12_ha6_out(.a(s_dadda_cska12_and_1_6[0]), .b(s_dadda_cska12_and_0_7[0]), .ha_xor0(s_dadda_cska12_ha6_xor0), .ha_and0(s_dadda_cska12_ha6_and0));
  fa fa_s_dadda_cska12_fa15_out(.a(s_dadda_cska12_ha6_and0[0]), .b(s_dadda_cska12_fa14_or0[0]), .cin(s_dadda_cska12_fa13_or0[0]), .fa_xor1(s_dadda_cska12_fa15_xor1), .fa_or0(s_dadda_cska12_fa15_or0));
  and_gate and_gate_s_dadda_cska12_and_8_0(.a(a[8]), .b(b[0]), .out(s_dadda_cska12_and_8_0));
  and_gate and_gate_s_dadda_cska12_and_7_1(.a(a[7]), .b(b[1]), .out(s_dadda_cska12_and_7_1));
  fa fa_s_dadda_cska12_fa16_out(.a(s_dadda_cska12_fa12_or0[0]), .b(s_dadda_cska12_and_8_0[0]), .cin(s_dadda_cska12_and_7_1[0]), .fa_xor1(s_dadda_cska12_fa16_xor1), .fa_or0(s_dadda_cska12_fa16_or0));
  and_gate and_gate_s_dadda_cska12_and_6_2(.a(a[6]), .b(b[2]), .out(s_dadda_cska12_and_6_2));
  and_gate and_gate_s_dadda_cska12_and_5_3(.a(a[5]), .b(b[3]), .out(s_dadda_cska12_and_5_3));
  and_gate and_gate_s_dadda_cska12_and_4_4(.a(a[4]), .b(b[4]), .out(s_dadda_cska12_and_4_4));
  fa fa_s_dadda_cska12_fa17_out(.a(s_dadda_cska12_and_6_2[0]), .b(s_dadda_cska12_and_5_3[0]), .cin(s_dadda_cska12_and_4_4[0]), .fa_xor1(s_dadda_cska12_fa17_xor1), .fa_or0(s_dadda_cska12_fa17_or0));
  and_gate and_gate_s_dadda_cska12_and_3_5(.a(a[3]), .b(b[5]), .out(s_dadda_cska12_and_3_5));
  and_gate and_gate_s_dadda_cska12_and_2_6(.a(a[2]), .b(b[6]), .out(s_dadda_cska12_and_2_6));
  and_gate and_gate_s_dadda_cska12_and_1_7(.a(a[1]), .b(b[7]), .out(s_dadda_cska12_and_1_7));
  fa fa_s_dadda_cska12_fa18_out(.a(s_dadda_cska12_and_3_5[0]), .b(s_dadda_cska12_and_2_6[0]), .cin(s_dadda_cska12_and_1_7[0]), .fa_xor1(s_dadda_cska12_fa18_xor1), .fa_or0(s_dadda_cska12_fa18_or0));
  and_gate and_gate_s_dadda_cska12_and_0_8(.a(a[0]), .b(b[8]), .out(s_dadda_cska12_and_0_8));
  ha ha_s_dadda_cska12_ha7_out(.a(s_dadda_cska12_and_0_8[0]), .b(s_dadda_cska12_fa15_xor1[0]), .ha_xor0(s_dadda_cska12_ha7_xor0), .ha_and0(s_dadda_cska12_ha7_and0));
  fa fa_s_dadda_cska12_fa19_out(.a(s_dadda_cska12_ha7_and0[0]), .b(s_dadda_cska12_fa18_or0[0]), .cin(s_dadda_cska12_fa17_or0[0]), .fa_xor1(s_dadda_cska12_fa19_xor1), .fa_or0(s_dadda_cska12_fa19_or0));
  and_gate and_gate_s_dadda_cska12_and_7_2(.a(a[7]), .b(b[2]), .out(s_dadda_cska12_and_7_2));
  fa fa_s_dadda_cska12_fa20_out(.a(s_dadda_cska12_fa16_or0[0]), .b(s_dadda_cska12_fa15_or0[0]), .cin(s_dadda_cska12_and_7_2[0]), .fa_xor1(s_dadda_cska12_fa20_xor1), .fa_or0(s_dadda_cska12_fa20_or0));
  and_gate and_gate_s_dadda_cska12_and_6_3(.a(a[6]), .b(b[3]), .out(s_dadda_cska12_and_6_3));
  and_gate and_gate_s_dadda_cska12_and_5_4(.a(a[5]), .b(b[4]), .out(s_dadda_cska12_and_5_4));
  and_gate and_gate_s_dadda_cska12_and_4_5(.a(a[4]), .b(b[5]), .out(s_dadda_cska12_and_4_5));
  fa fa_s_dadda_cska12_fa21_out(.a(s_dadda_cska12_and_6_3[0]), .b(s_dadda_cska12_and_5_4[0]), .cin(s_dadda_cska12_and_4_5[0]), .fa_xor1(s_dadda_cska12_fa21_xor1), .fa_or0(s_dadda_cska12_fa21_or0));
  and_gate and_gate_s_dadda_cska12_and_3_6(.a(a[3]), .b(b[6]), .out(s_dadda_cska12_and_3_6));
  and_gate and_gate_s_dadda_cska12_and_2_7(.a(a[2]), .b(b[7]), .out(s_dadda_cska12_and_2_7));
  and_gate and_gate_s_dadda_cska12_and_1_8(.a(a[1]), .b(b[8]), .out(s_dadda_cska12_and_1_8));
  fa fa_s_dadda_cska12_fa22_out(.a(s_dadda_cska12_and_3_6[0]), .b(s_dadda_cska12_and_2_7[0]), .cin(s_dadda_cska12_and_1_8[0]), .fa_xor1(s_dadda_cska12_fa22_xor1), .fa_or0(s_dadda_cska12_fa22_or0));
  and_gate and_gate_s_dadda_cska12_and_0_9(.a(a[0]), .b(b[9]), .out(s_dadda_cska12_and_0_9));
  fa fa_s_dadda_cska12_fa23_out(.a(s_dadda_cska12_and_0_9[0]), .b(s_dadda_cska12_ha0_xor0[0]), .cin(s_dadda_cska12_fa19_xor1[0]), .fa_xor1(s_dadda_cska12_fa23_xor1), .fa_or0(s_dadda_cska12_fa23_or0));
  fa fa_s_dadda_cska12_fa24_out(.a(s_dadda_cska12_fa23_or0[0]), .b(s_dadda_cska12_fa22_or0[0]), .cin(s_dadda_cska12_fa21_or0[0]), .fa_xor1(s_dadda_cska12_fa24_xor1), .fa_or0(s_dadda_cska12_fa24_or0));
  and_gate and_gate_s_dadda_cska12_and_6_4(.a(a[6]), .b(b[4]), .out(s_dadda_cska12_and_6_4));
  fa fa_s_dadda_cska12_fa25_out(.a(s_dadda_cska12_fa20_or0[0]), .b(s_dadda_cska12_fa19_or0[0]), .cin(s_dadda_cska12_and_6_4[0]), .fa_xor1(s_dadda_cska12_fa25_xor1), .fa_or0(s_dadda_cska12_fa25_or0));
  and_gate and_gate_s_dadda_cska12_and_5_5(.a(a[5]), .b(b[5]), .out(s_dadda_cska12_and_5_5));
  and_gate and_gate_s_dadda_cska12_and_4_6(.a(a[4]), .b(b[6]), .out(s_dadda_cska12_and_4_6));
  and_gate and_gate_s_dadda_cska12_and_3_7(.a(a[3]), .b(b[7]), .out(s_dadda_cska12_and_3_7));
  fa fa_s_dadda_cska12_fa26_out(.a(s_dadda_cska12_and_5_5[0]), .b(s_dadda_cska12_and_4_6[0]), .cin(s_dadda_cska12_and_3_7[0]), .fa_xor1(s_dadda_cska12_fa26_xor1), .fa_or0(s_dadda_cska12_fa26_or0));
  and_gate and_gate_s_dadda_cska12_and_2_8(.a(a[2]), .b(b[8]), .out(s_dadda_cska12_and_2_8));
  and_gate and_gate_s_dadda_cska12_and_1_9(.a(a[1]), .b(b[9]), .out(s_dadda_cska12_and_1_9));
  and_gate and_gate_s_dadda_cska12_and_0_10(.a(a[0]), .b(b[10]), .out(s_dadda_cska12_and_0_10));
  fa fa_s_dadda_cska12_fa27_out(.a(s_dadda_cska12_and_2_8[0]), .b(s_dadda_cska12_and_1_9[0]), .cin(s_dadda_cska12_and_0_10[0]), .fa_xor1(s_dadda_cska12_fa27_xor1), .fa_or0(s_dadda_cska12_fa27_or0));
  fa fa_s_dadda_cska12_fa28_out(.a(s_dadda_cska12_fa0_xor1[0]), .b(s_dadda_cska12_ha1_xor0[0]), .cin(s_dadda_cska12_fa24_xor1[0]), .fa_xor1(s_dadda_cska12_fa28_xor1), .fa_or0(s_dadda_cska12_fa28_or0));
  fa fa_s_dadda_cska12_fa29_out(.a(s_dadda_cska12_fa28_or0[0]), .b(s_dadda_cska12_fa27_or0[0]), .cin(s_dadda_cska12_fa26_or0[0]), .fa_xor1(s_dadda_cska12_fa29_xor1), .fa_or0(s_dadda_cska12_fa29_or0));
  and_gate and_gate_s_dadda_cska12_and_5_6(.a(a[5]), .b(b[6]), .out(s_dadda_cska12_and_5_6));
  fa fa_s_dadda_cska12_fa30_out(.a(s_dadda_cska12_fa25_or0[0]), .b(s_dadda_cska12_fa24_or0[0]), .cin(s_dadda_cska12_and_5_6[0]), .fa_xor1(s_dadda_cska12_fa30_xor1), .fa_or0(s_dadda_cska12_fa30_or0));
  and_gate and_gate_s_dadda_cska12_and_4_7(.a(a[4]), .b(b[7]), .out(s_dadda_cska12_and_4_7));
  and_gate and_gate_s_dadda_cska12_and_3_8(.a(a[3]), .b(b[8]), .out(s_dadda_cska12_and_3_8));
  and_gate and_gate_s_dadda_cska12_and_2_9(.a(a[2]), .b(b[9]), .out(s_dadda_cska12_and_2_9));
  fa fa_s_dadda_cska12_fa31_out(.a(s_dadda_cska12_and_4_7[0]), .b(s_dadda_cska12_and_3_8[0]), .cin(s_dadda_cska12_and_2_9[0]), .fa_xor1(s_dadda_cska12_fa31_xor1), .fa_or0(s_dadda_cska12_fa31_or0));
  and_gate and_gate_s_dadda_cska12_and_1_10(.a(a[1]), .b(b[10]), .out(s_dadda_cska12_and_1_10));
  nand_gate nand_gate_s_dadda_cska12_nand_0_11(.a(a[0]), .b(b[11]), .out(s_dadda_cska12_nand_0_11));
  fa fa_s_dadda_cska12_fa32_out(.a(s_dadda_cska12_and_1_10[0]), .b(s_dadda_cska12_nand_0_11[0]), .cin(s_dadda_cska12_fa1_xor1[0]), .fa_xor1(s_dadda_cska12_fa32_xor1), .fa_or0(s_dadda_cska12_fa32_or0));
  fa fa_s_dadda_cska12_fa33_out(.a(s_dadda_cska12_fa2_xor1[0]), .b(s_dadda_cska12_ha2_xor0[0]), .cin(s_dadda_cska12_fa29_xor1[0]), .fa_xor1(s_dadda_cska12_fa33_xor1), .fa_or0(s_dadda_cska12_fa33_or0));
  fa fa_s_dadda_cska12_fa34_out(.a(s_dadda_cska12_fa33_or0[0]), .b(s_dadda_cska12_fa32_or0[0]), .cin(s_dadda_cska12_fa31_or0[0]), .fa_xor1(s_dadda_cska12_fa34_xor1), .fa_or0(s_dadda_cska12_fa34_or0));
  and_gate and_gate_s_dadda_cska12_and_6_6(.a(a[6]), .b(b[6]), .out(s_dadda_cska12_and_6_6));
  fa fa_s_dadda_cska12_fa35_out(.a(s_dadda_cska12_fa30_or0[0]), .b(s_dadda_cska12_fa29_or0[0]), .cin(s_dadda_cska12_and_6_6[0]), .fa_xor1(s_dadda_cska12_fa35_xor1), .fa_or0(s_dadda_cska12_fa35_or0));
  and_gate and_gate_s_dadda_cska12_and_5_7(.a(a[5]), .b(b[7]), .out(s_dadda_cska12_and_5_7));
  and_gate and_gate_s_dadda_cska12_and_4_8(.a(a[4]), .b(b[8]), .out(s_dadda_cska12_and_4_8));
  and_gate and_gate_s_dadda_cska12_and_3_9(.a(a[3]), .b(b[9]), .out(s_dadda_cska12_and_3_9));
  fa fa_s_dadda_cska12_fa36_out(.a(s_dadda_cska12_and_5_7[0]), .b(s_dadda_cska12_and_4_8[0]), .cin(s_dadda_cska12_and_3_9[0]), .fa_xor1(s_dadda_cska12_fa36_xor1), .fa_or0(s_dadda_cska12_fa36_or0));
  and_gate and_gate_s_dadda_cska12_and_2_10(.a(a[2]), .b(b[10]), .out(s_dadda_cska12_and_2_10));
  nand_gate nand_gate_s_dadda_cska12_nand_1_11(.a(a[1]), .b(b[11]), .out(s_dadda_cska12_nand_1_11));
  fa fa_s_dadda_cska12_fa37_out(.a(s_dadda_cska12_and_2_10[0]), .b(s_dadda_cska12_nand_1_11[0]), .cin(s_dadda_cska12_fa3_xor1[0]), .fa_xor1(s_dadda_cska12_fa37_xor1), .fa_or0(s_dadda_cska12_fa37_or0));
  fa fa_s_dadda_cska12_fa38_out(.a(s_dadda_cska12_fa4_xor1[0]), .b(s_dadda_cska12_fa5_xor1[0]), .cin(s_dadda_cska12_fa34_xor1[0]), .fa_xor1(s_dadda_cska12_fa38_xor1), .fa_or0(s_dadda_cska12_fa38_or0));
  fa fa_s_dadda_cska12_fa39_out(.a(s_dadda_cska12_fa38_or0[0]), .b(s_dadda_cska12_fa37_or0[0]), .cin(s_dadda_cska12_fa36_or0[0]), .fa_xor1(s_dadda_cska12_fa39_xor1), .fa_or0(s_dadda_cska12_fa39_or0));
  and_gate and_gate_s_dadda_cska12_and_8_5(.a(a[8]), .b(b[5]), .out(s_dadda_cska12_and_8_5));
  fa fa_s_dadda_cska12_fa40_out(.a(s_dadda_cska12_fa35_or0[0]), .b(s_dadda_cska12_fa34_or0[0]), .cin(s_dadda_cska12_and_8_5[0]), .fa_xor1(s_dadda_cska12_fa40_xor1), .fa_or0(s_dadda_cska12_fa40_or0));
  and_gate and_gate_s_dadda_cska12_and_7_6(.a(a[7]), .b(b[6]), .out(s_dadda_cska12_and_7_6));
  and_gate and_gate_s_dadda_cska12_and_6_7(.a(a[6]), .b(b[7]), .out(s_dadda_cska12_and_6_7));
  and_gate and_gate_s_dadda_cska12_and_5_8(.a(a[5]), .b(b[8]), .out(s_dadda_cska12_and_5_8));
  fa fa_s_dadda_cska12_fa41_out(.a(s_dadda_cska12_and_7_6[0]), .b(s_dadda_cska12_and_6_7[0]), .cin(s_dadda_cska12_and_5_8[0]), .fa_xor1(s_dadda_cska12_fa41_xor1), .fa_or0(s_dadda_cska12_fa41_or0));
  and_gate and_gate_s_dadda_cska12_and_4_9(.a(a[4]), .b(b[9]), .out(s_dadda_cska12_and_4_9));
  and_gate and_gate_s_dadda_cska12_and_3_10(.a(a[3]), .b(b[10]), .out(s_dadda_cska12_and_3_10));
  nand_gate nand_gate_s_dadda_cska12_nand_2_11(.a(a[2]), .b(b[11]), .out(s_dadda_cska12_nand_2_11));
  fa fa_s_dadda_cska12_fa42_out(.a(s_dadda_cska12_and_4_9[0]), .b(s_dadda_cska12_and_3_10[0]), .cin(s_dadda_cska12_nand_2_11[0]), .fa_xor1(s_dadda_cska12_fa42_xor1), .fa_or0(s_dadda_cska12_fa42_or0));
  fa fa_s_dadda_cska12_fa43_out(.a(s_dadda_cska12_fa6_xor1[0]), .b(s_dadda_cska12_fa7_xor1[0]), .cin(s_dadda_cska12_fa39_xor1[0]), .fa_xor1(s_dadda_cska12_fa43_xor1), .fa_or0(s_dadda_cska12_fa43_or0));
  fa fa_s_dadda_cska12_fa44_out(.a(s_dadda_cska12_fa43_or0[0]), .b(s_dadda_cska12_fa42_or0[0]), .cin(s_dadda_cska12_fa41_or0[0]), .fa_xor1(s_dadda_cska12_fa44_xor1), .fa_or0(s_dadda_cska12_fa44_or0));
  and_gate and_gate_s_dadda_cska12_and_10_4(.a(a[10]), .b(b[4]), .out(s_dadda_cska12_and_10_4));
  fa fa_s_dadda_cska12_fa45_out(.a(s_dadda_cska12_fa40_or0[0]), .b(s_dadda_cska12_fa39_or0[0]), .cin(s_dadda_cska12_and_10_4[0]), .fa_xor1(s_dadda_cska12_fa45_xor1), .fa_or0(s_dadda_cska12_fa45_or0));
  and_gate and_gate_s_dadda_cska12_and_9_5(.a(a[9]), .b(b[5]), .out(s_dadda_cska12_and_9_5));
  and_gate and_gate_s_dadda_cska12_and_8_6(.a(a[8]), .b(b[6]), .out(s_dadda_cska12_and_8_6));
  and_gate and_gate_s_dadda_cska12_and_7_7(.a(a[7]), .b(b[7]), .out(s_dadda_cska12_and_7_7));
  fa fa_s_dadda_cska12_fa46_out(.a(s_dadda_cska12_and_9_5[0]), .b(s_dadda_cska12_and_8_6[0]), .cin(s_dadda_cska12_and_7_7[0]), .fa_xor1(s_dadda_cska12_fa46_xor1), .fa_or0(s_dadda_cska12_fa46_or0));
  and_gate and_gate_s_dadda_cska12_and_6_8(.a(a[6]), .b(b[8]), .out(s_dadda_cska12_and_6_8));
  and_gate and_gate_s_dadda_cska12_and_5_9(.a(a[5]), .b(b[9]), .out(s_dadda_cska12_and_5_9));
  and_gate and_gate_s_dadda_cska12_and_4_10(.a(a[4]), .b(b[10]), .out(s_dadda_cska12_and_4_10));
  fa fa_s_dadda_cska12_fa47_out(.a(s_dadda_cska12_and_6_8[0]), .b(s_dadda_cska12_and_5_9[0]), .cin(s_dadda_cska12_and_4_10[0]), .fa_xor1(s_dadda_cska12_fa47_xor1), .fa_or0(s_dadda_cska12_fa47_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_3_11(.a(a[3]), .b(b[11]), .out(s_dadda_cska12_nand_3_11));
  fa fa_s_dadda_cska12_fa48_out(.a(s_dadda_cska12_nand_3_11[0]), .b(s_dadda_cska12_fa8_xor1[0]), .cin(s_dadda_cska12_fa44_xor1[0]), .fa_xor1(s_dadda_cska12_fa48_xor1), .fa_or0(s_dadda_cska12_fa48_or0));
  fa fa_s_dadda_cska12_fa49_out(.a(s_dadda_cska12_fa48_or0[0]), .b(s_dadda_cska12_fa47_or0[0]), .cin(s_dadda_cska12_fa46_or0[0]), .fa_xor1(s_dadda_cska12_fa49_xor1), .fa_or0(s_dadda_cska12_fa49_or0));
  fa fa_s_dadda_cska12_fa50_out(.a(s_dadda_cska12_fa45_or0[0]), .b(s_dadda_cska12_fa44_or0[0]), .cin(s_dadda_cska12_fa8_or0[0]), .fa_xor1(s_dadda_cska12_fa50_xor1), .fa_or0(s_dadda_cska12_fa50_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_4(.a(a[11]), .b(b[4]), .out(s_dadda_cska12_nand_11_4));
  and_gate and_gate_s_dadda_cska12_and_10_5(.a(a[10]), .b(b[5]), .out(s_dadda_cska12_and_10_5));
  and_gate and_gate_s_dadda_cska12_and_9_6(.a(a[9]), .b(b[6]), .out(s_dadda_cska12_and_9_6));
  fa fa_s_dadda_cska12_fa51_out(.a(s_dadda_cska12_nand_11_4[0]), .b(s_dadda_cska12_and_10_5[0]), .cin(s_dadda_cska12_and_9_6[0]), .fa_xor1(s_dadda_cska12_fa51_xor1), .fa_or0(s_dadda_cska12_fa51_or0));
  and_gate and_gate_s_dadda_cska12_and_8_7(.a(a[8]), .b(b[7]), .out(s_dadda_cska12_and_8_7));
  and_gate and_gate_s_dadda_cska12_and_7_8(.a(a[7]), .b(b[8]), .out(s_dadda_cska12_and_7_8));
  and_gate and_gate_s_dadda_cska12_and_6_9(.a(a[6]), .b(b[9]), .out(s_dadda_cska12_and_6_9));
  fa fa_s_dadda_cska12_fa52_out(.a(s_dadda_cska12_and_8_7[0]), .b(s_dadda_cska12_and_7_8[0]), .cin(s_dadda_cska12_and_6_9[0]), .fa_xor1(s_dadda_cska12_fa52_xor1), .fa_or0(s_dadda_cska12_fa52_or0));
  and_gate and_gate_s_dadda_cska12_and_5_10(.a(a[5]), .b(b[10]), .out(s_dadda_cska12_and_5_10));
  nand_gate nand_gate_s_dadda_cska12_nand_4_11(.a(a[4]), .b(b[11]), .out(s_dadda_cska12_nand_4_11));
  fa fa_s_dadda_cska12_fa53_out(.a(s_dadda_cska12_and_5_10[0]), .b(s_dadda_cska12_nand_4_11[0]), .cin(s_dadda_cska12_fa49_xor1[0]), .fa_xor1(s_dadda_cska12_fa53_xor1), .fa_or0(s_dadda_cska12_fa53_or0));
  fa fa_s_dadda_cska12_fa54_out(.a(s_dadda_cska12_fa53_or0[0]), .b(s_dadda_cska12_fa52_or0[0]), .cin(s_dadda_cska12_fa51_or0[0]), .fa_xor1(s_dadda_cska12_fa54_xor1), .fa_or0(s_dadda_cska12_fa54_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_5(.a(a[11]), .b(b[5]), .out(s_dadda_cska12_nand_11_5));
  fa fa_s_dadda_cska12_fa55_out(.a(s_dadda_cska12_fa50_or0[0]), .b(s_dadda_cska12_fa49_or0[0]), .cin(s_dadda_cska12_nand_11_5[0]), .fa_xor1(s_dadda_cska12_fa55_xor1), .fa_or0(s_dadda_cska12_fa55_or0));
  and_gate and_gate_s_dadda_cska12_and_10_6(.a(a[10]), .b(b[6]), .out(s_dadda_cska12_and_10_6));
  and_gate and_gate_s_dadda_cska12_and_9_7(.a(a[9]), .b(b[7]), .out(s_dadda_cska12_and_9_7));
  and_gate and_gate_s_dadda_cska12_and_8_8(.a(a[8]), .b(b[8]), .out(s_dadda_cska12_and_8_8));
  fa fa_s_dadda_cska12_fa56_out(.a(s_dadda_cska12_and_10_6[0]), .b(s_dadda_cska12_and_9_7[0]), .cin(s_dadda_cska12_and_8_8[0]), .fa_xor1(s_dadda_cska12_fa56_xor1), .fa_or0(s_dadda_cska12_fa56_or0));
  and_gate and_gate_s_dadda_cska12_and_7_9(.a(a[7]), .b(b[9]), .out(s_dadda_cska12_and_7_9));
  and_gate and_gate_s_dadda_cska12_and_6_10(.a(a[6]), .b(b[10]), .out(s_dadda_cska12_and_6_10));
  nand_gate nand_gate_s_dadda_cska12_nand_5_11(.a(a[5]), .b(b[11]), .out(s_dadda_cska12_nand_5_11));
  fa fa_s_dadda_cska12_fa57_out(.a(s_dadda_cska12_and_7_9[0]), .b(s_dadda_cska12_and_6_10[0]), .cin(s_dadda_cska12_nand_5_11[0]), .fa_xor1(s_dadda_cska12_fa57_xor1), .fa_or0(s_dadda_cska12_fa57_or0));
  fa fa_s_dadda_cska12_fa58_out(.a(s_dadda_cska12_fa57_or0[0]), .b(s_dadda_cska12_fa56_or0[0]), .cin(s_dadda_cska12_fa55_or0[0]), .fa_xor1(s_dadda_cska12_fa58_xor1), .fa_or0(s_dadda_cska12_fa58_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_6(.a(a[11]), .b(b[6]), .out(s_dadda_cska12_nand_11_6));
  and_gate and_gate_s_dadda_cska12_and_10_7(.a(a[10]), .b(b[7]), .out(s_dadda_cska12_and_10_7));
  fa fa_s_dadda_cska12_fa59_out(.a(s_dadda_cska12_fa54_or0[0]), .b(s_dadda_cska12_nand_11_6[0]), .cin(s_dadda_cska12_and_10_7[0]), .fa_xor1(s_dadda_cska12_fa59_xor1), .fa_or0(s_dadda_cska12_fa59_or0));
  and_gate and_gate_s_dadda_cska12_and_9_8(.a(a[9]), .b(b[8]), .out(s_dadda_cska12_and_9_8));
  and_gate and_gate_s_dadda_cska12_and_8_9(.a(a[8]), .b(b[9]), .out(s_dadda_cska12_and_8_9));
  and_gate and_gate_s_dadda_cska12_and_7_10(.a(a[7]), .b(b[10]), .out(s_dadda_cska12_and_7_10));
  fa fa_s_dadda_cska12_fa60_out(.a(s_dadda_cska12_and_9_8[0]), .b(s_dadda_cska12_and_8_9[0]), .cin(s_dadda_cska12_and_7_10[0]), .fa_xor1(s_dadda_cska12_fa60_xor1), .fa_or0(s_dadda_cska12_fa60_or0));
  fa fa_s_dadda_cska12_fa61_out(.a(s_dadda_cska12_fa60_or0[0]), .b(s_dadda_cska12_fa59_or0[0]), .cin(s_dadda_cska12_fa58_or0[0]), .fa_xor1(s_dadda_cska12_fa61_xor1), .fa_or0(s_dadda_cska12_fa61_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_7(.a(a[11]), .b(b[7]), .out(s_dadda_cska12_nand_11_7));
  and_gate and_gate_s_dadda_cska12_and_10_8(.a(a[10]), .b(b[8]), .out(s_dadda_cska12_and_10_8));
  and_gate and_gate_s_dadda_cska12_and_9_9(.a(a[9]), .b(b[9]), .out(s_dadda_cska12_and_9_9));
  fa fa_s_dadda_cska12_fa62_out(.a(s_dadda_cska12_nand_11_7[0]), .b(s_dadda_cska12_and_10_8[0]), .cin(s_dadda_cska12_and_9_9[0]), .fa_xor1(s_dadda_cska12_fa62_xor1), .fa_or0(s_dadda_cska12_fa62_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_8(.a(a[11]), .b(b[8]), .out(s_dadda_cska12_nand_11_8));
  fa fa_s_dadda_cska12_fa63_out(.a(s_dadda_cska12_fa62_or0[0]), .b(s_dadda_cska12_fa61_or0[0]), .cin(s_dadda_cska12_nand_11_8[0]), .fa_xor1(s_dadda_cska12_fa63_xor1), .fa_or0(s_dadda_cska12_fa63_or0));
  and_gate and_gate_s_dadda_cska12_and_3_0(.a(a[3]), .b(b[0]), .out(s_dadda_cska12_and_3_0));
  and_gate and_gate_s_dadda_cska12_and_2_1(.a(a[2]), .b(b[1]), .out(s_dadda_cska12_and_2_1));
  ha ha_s_dadda_cska12_ha8_out(.a(s_dadda_cska12_and_3_0[0]), .b(s_dadda_cska12_and_2_1[0]), .ha_xor0(s_dadda_cska12_ha8_xor0), .ha_and0(s_dadda_cska12_ha8_and0));
  and_gate and_gate_s_dadda_cska12_and_2_2(.a(a[2]), .b(b[2]), .out(s_dadda_cska12_and_2_2));
  and_gate and_gate_s_dadda_cska12_and_1_3(.a(a[1]), .b(b[3]), .out(s_dadda_cska12_and_1_3));
  fa fa_s_dadda_cska12_fa64_out(.a(s_dadda_cska12_ha8_and0[0]), .b(s_dadda_cska12_and_2_2[0]), .cin(s_dadda_cska12_and_1_3[0]), .fa_xor1(s_dadda_cska12_fa64_xor1), .fa_or0(s_dadda_cska12_fa64_or0));
  and_gate and_gate_s_dadda_cska12_and_1_4(.a(a[1]), .b(b[4]), .out(s_dadda_cska12_and_1_4));
  and_gate and_gate_s_dadda_cska12_and_0_5(.a(a[0]), .b(b[5]), .out(s_dadda_cska12_and_0_5));
  fa fa_s_dadda_cska12_fa65_out(.a(s_dadda_cska12_fa64_or0[0]), .b(s_dadda_cska12_and_1_4[0]), .cin(s_dadda_cska12_and_0_5[0]), .fa_xor1(s_dadda_cska12_fa65_xor1), .fa_or0(s_dadda_cska12_fa65_or0));
  and_gate and_gate_s_dadda_cska12_and_0_6(.a(a[0]), .b(b[6]), .out(s_dadda_cska12_and_0_6));
  fa fa_s_dadda_cska12_fa66_out(.a(s_dadda_cska12_fa65_or0[0]), .b(s_dadda_cska12_and_0_6[0]), .cin(s_dadda_cska12_fa10_xor1[0]), .fa_xor1(s_dadda_cska12_fa66_xor1), .fa_or0(s_dadda_cska12_fa66_or0));
  fa fa_s_dadda_cska12_fa67_out(.a(s_dadda_cska12_fa66_or0[0]), .b(s_dadda_cska12_fa12_xor1[0]), .cin(s_dadda_cska12_fa13_xor1[0]), .fa_xor1(s_dadda_cska12_fa67_xor1), .fa_or0(s_dadda_cska12_fa67_or0));
  fa fa_s_dadda_cska12_fa68_out(.a(s_dadda_cska12_fa67_or0[0]), .b(s_dadda_cska12_fa16_xor1[0]), .cin(s_dadda_cska12_fa17_xor1[0]), .fa_xor1(s_dadda_cska12_fa68_xor1), .fa_or0(s_dadda_cska12_fa68_or0));
  fa fa_s_dadda_cska12_fa69_out(.a(s_dadda_cska12_fa68_or0[0]), .b(s_dadda_cska12_fa20_xor1[0]), .cin(s_dadda_cska12_fa21_xor1[0]), .fa_xor1(s_dadda_cska12_fa69_xor1), .fa_or0(s_dadda_cska12_fa69_or0));
  fa fa_s_dadda_cska12_fa70_out(.a(s_dadda_cska12_fa69_or0[0]), .b(s_dadda_cska12_fa25_xor1[0]), .cin(s_dadda_cska12_fa26_xor1[0]), .fa_xor1(s_dadda_cska12_fa70_xor1), .fa_or0(s_dadda_cska12_fa70_or0));
  fa fa_s_dadda_cska12_fa71_out(.a(s_dadda_cska12_fa70_or0[0]), .b(s_dadda_cska12_fa30_xor1[0]), .cin(s_dadda_cska12_fa31_xor1[0]), .fa_xor1(s_dadda_cska12_fa71_xor1), .fa_or0(s_dadda_cska12_fa71_or0));
  fa fa_s_dadda_cska12_fa72_out(.a(s_dadda_cska12_fa71_or0[0]), .b(s_dadda_cska12_fa35_xor1[0]), .cin(s_dadda_cska12_fa36_xor1[0]), .fa_xor1(s_dadda_cska12_fa72_xor1), .fa_or0(s_dadda_cska12_fa72_or0));
  fa fa_s_dadda_cska12_fa73_out(.a(s_dadda_cska12_fa72_or0[0]), .b(s_dadda_cska12_fa40_xor1[0]), .cin(s_dadda_cska12_fa41_xor1[0]), .fa_xor1(s_dadda_cska12_fa73_xor1), .fa_or0(s_dadda_cska12_fa73_or0));
  fa fa_s_dadda_cska12_fa74_out(.a(s_dadda_cska12_fa73_or0[0]), .b(s_dadda_cska12_fa45_xor1[0]), .cin(s_dadda_cska12_fa46_xor1[0]), .fa_xor1(s_dadda_cska12_fa74_xor1), .fa_or0(s_dadda_cska12_fa74_or0));
  fa fa_s_dadda_cska12_fa75_out(.a(s_dadda_cska12_fa74_or0[0]), .b(s_dadda_cska12_fa50_xor1[0]), .cin(s_dadda_cska12_fa51_xor1[0]), .fa_xor1(s_dadda_cska12_fa75_xor1), .fa_or0(s_dadda_cska12_fa75_or0));
  fa fa_s_dadda_cska12_fa76_out(.a(s_dadda_cska12_fa75_or0[0]), .b(s_dadda_cska12_fa54_xor1[0]), .cin(s_dadda_cska12_fa55_xor1[0]), .fa_xor1(s_dadda_cska12_fa76_xor1), .fa_or0(s_dadda_cska12_fa76_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_6_11(.a(a[6]), .b(b[11]), .out(s_dadda_cska12_nand_6_11));
  fa fa_s_dadda_cska12_fa77_out(.a(s_dadda_cska12_fa76_or0[0]), .b(s_dadda_cska12_nand_6_11[0]), .cin(s_dadda_cska12_fa58_xor1[0]), .fa_xor1(s_dadda_cska12_fa77_xor1), .fa_or0(s_dadda_cska12_fa77_or0));
  and_gate and_gate_s_dadda_cska12_and_8_10(.a(a[8]), .b(b[10]), .out(s_dadda_cska12_and_8_10));
  nand_gate nand_gate_s_dadda_cska12_nand_7_11(.a(a[7]), .b(b[11]), .out(s_dadda_cska12_nand_7_11));
  fa fa_s_dadda_cska12_fa78_out(.a(s_dadda_cska12_fa77_or0[0]), .b(s_dadda_cska12_and_8_10[0]), .cin(s_dadda_cska12_nand_7_11[0]), .fa_xor1(s_dadda_cska12_fa78_xor1), .fa_or0(s_dadda_cska12_fa78_or0));
  and_gate and_gate_s_dadda_cska12_and_10_9(.a(a[10]), .b(b[9]), .out(s_dadda_cska12_and_10_9));
  and_gate and_gate_s_dadda_cska12_and_9_10(.a(a[9]), .b(b[10]), .out(s_dadda_cska12_and_9_10));
  fa fa_s_dadda_cska12_fa79_out(.a(s_dadda_cska12_fa78_or0[0]), .b(s_dadda_cska12_and_10_9[0]), .cin(s_dadda_cska12_and_9_10[0]), .fa_xor1(s_dadda_cska12_fa79_xor1), .fa_or0(s_dadda_cska12_fa79_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_9(.a(a[11]), .b(b[9]), .out(s_dadda_cska12_nand_11_9));
  fa fa_s_dadda_cska12_fa80_out(.a(s_dadda_cska12_fa79_or0[0]), .b(s_dadda_cska12_fa63_or0[0]), .cin(s_dadda_cska12_nand_11_9[0]), .fa_xor1(s_dadda_cska12_fa80_xor1), .fa_or0(s_dadda_cska12_fa80_or0));
  and_gate and_gate_s_dadda_cska12_and_2_0(.a(a[2]), .b(b[0]), .out(s_dadda_cska12_and_2_0));
  and_gate and_gate_s_dadda_cska12_and_1_1(.a(a[1]), .b(b[1]), .out(s_dadda_cska12_and_1_1));
  ha ha_s_dadda_cska12_ha9_out(.a(s_dadda_cska12_and_2_0[0]), .b(s_dadda_cska12_and_1_1[0]), .ha_xor0(s_dadda_cska12_ha9_xor0), .ha_and0(s_dadda_cska12_ha9_and0));
  and_gate and_gate_s_dadda_cska12_and_1_2(.a(a[1]), .b(b[2]), .out(s_dadda_cska12_and_1_2));
  and_gate and_gate_s_dadda_cska12_and_0_3(.a(a[0]), .b(b[3]), .out(s_dadda_cska12_and_0_3));
  fa fa_s_dadda_cska12_fa81_out(.a(s_dadda_cska12_ha9_and0[0]), .b(s_dadda_cska12_and_1_2[0]), .cin(s_dadda_cska12_and_0_3[0]), .fa_xor1(s_dadda_cska12_fa81_xor1), .fa_or0(s_dadda_cska12_fa81_or0));
  and_gate and_gate_s_dadda_cska12_and_0_4(.a(a[0]), .b(b[4]), .out(s_dadda_cska12_and_0_4));
  fa fa_s_dadda_cska12_fa82_out(.a(s_dadda_cska12_fa81_or0[0]), .b(s_dadda_cska12_and_0_4[0]), .cin(s_dadda_cska12_ha3_xor0[0]), .fa_xor1(s_dadda_cska12_fa82_xor1), .fa_or0(s_dadda_cska12_fa82_or0));
  fa fa_s_dadda_cska12_fa83_out(.a(s_dadda_cska12_fa82_or0[0]), .b(s_dadda_cska12_fa9_xor1[0]), .cin(s_dadda_cska12_ha4_xor0[0]), .fa_xor1(s_dadda_cska12_fa83_xor1), .fa_or0(s_dadda_cska12_fa83_or0));
  fa fa_s_dadda_cska12_fa84_out(.a(s_dadda_cska12_fa83_or0[0]), .b(s_dadda_cska12_fa11_xor1[0]), .cin(s_dadda_cska12_ha5_xor0[0]), .fa_xor1(s_dadda_cska12_fa84_xor1), .fa_or0(s_dadda_cska12_fa84_or0));
  fa fa_s_dadda_cska12_fa85_out(.a(s_dadda_cska12_fa84_or0[0]), .b(s_dadda_cska12_fa14_xor1[0]), .cin(s_dadda_cska12_ha6_xor0[0]), .fa_xor1(s_dadda_cska12_fa85_xor1), .fa_or0(s_dadda_cska12_fa85_or0));
  fa fa_s_dadda_cska12_fa86_out(.a(s_dadda_cska12_fa85_or0[0]), .b(s_dadda_cska12_fa18_xor1[0]), .cin(s_dadda_cska12_ha7_xor0[0]), .fa_xor1(s_dadda_cska12_fa86_xor1), .fa_or0(s_dadda_cska12_fa86_or0));
  fa fa_s_dadda_cska12_fa87_out(.a(s_dadda_cska12_fa86_or0[0]), .b(s_dadda_cska12_fa22_xor1[0]), .cin(s_dadda_cska12_fa23_xor1[0]), .fa_xor1(s_dadda_cska12_fa87_xor1), .fa_or0(s_dadda_cska12_fa87_or0));
  fa fa_s_dadda_cska12_fa88_out(.a(s_dadda_cska12_fa87_or0[0]), .b(s_dadda_cska12_fa27_xor1[0]), .cin(s_dadda_cska12_fa28_xor1[0]), .fa_xor1(s_dadda_cska12_fa88_xor1), .fa_or0(s_dadda_cska12_fa88_or0));
  fa fa_s_dadda_cska12_fa89_out(.a(s_dadda_cska12_fa88_or0[0]), .b(s_dadda_cska12_fa32_xor1[0]), .cin(s_dadda_cska12_fa33_xor1[0]), .fa_xor1(s_dadda_cska12_fa89_xor1), .fa_or0(s_dadda_cska12_fa89_or0));
  fa fa_s_dadda_cska12_fa90_out(.a(s_dadda_cska12_fa89_or0[0]), .b(s_dadda_cska12_fa37_xor1[0]), .cin(s_dadda_cska12_fa38_xor1[0]), .fa_xor1(s_dadda_cska12_fa90_xor1), .fa_or0(s_dadda_cska12_fa90_or0));
  fa fa_s_dadda_cska12_fa91_out(.a(s_dadda_cska12_fa90_or0[0]), .b(s_dadda_cska12_fa42_xor1[0]), .cin(s_dadda_cska12_fa43_xor1[0]), .fa_xor1(s_dadda_cska12_fa91_xor1), .fa_or0(s_dadda_cska12_fa91_or0));
  fa fa_s_dadda_cska12_fa92_out(.a(s_dadda_cska12_fa91_or0[0]), .b(s_dadda_cska12_fa47_xor1[0]), .cin(s_dadda_cska12_fa48_xor1[0]), .fa_xor1(s_dadda_cska12_fa92_xor1), .fa_or0(s_dadda_cska12_fa92_or0));
  fa fa_s_dadda_cska12_fa93_out(.a(s_dadda_cska12_fa92_or0[0]), .b(s_dadda_cska12_fa52_xor1[0]), .cin(s_dadda_cska12_fa53_xor1[0]), .fa_xor1(s_dadda_cska12_fa93_xor1), .fa_or0(s_dadda_cska12_fa93_or0));
  fa fa_s_dadda_cska12_fa94_out(.a(s_dadda_cska12_fa93_or0[0]), .b(s_dadda_cska12_fa56_xor1[0]), .cin(s_dadda_cska12_fa57_xor1[0]), .fa_xor1(s_dadda_cska12_fa94_xor1), .fa_or0(s_dadda_cska12_fa94_or0));
  fa fa_s_dadda_cska12_fa95_out(.a(s_dadda_cska12_fa94_or0[0]), .b(s_dadda_cska12_fa59_xor1[0]), .cin(s_dadda_cska12_fa60_xor1[0]), .fa_xor1(s_dadda_cska12_fa95_xor1), .fa_or0(s_dadda_cska12_fa95_or0));
  fa fa_s_dadda_cska12_fa96_out(.a(s_dadda_cska12_fa95_or0[0]), .b(s_dadda_cska12_fa61_xor1[0]), .cin(s_dadda_cska12_fa62_xor1[0]), .fa_xor1(s_dadda_cska12_fa96_xor1), .fa_or0(s_dadda_cska12_fa96_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_8_11(.a(a[8]), .b(b[11]), .out(s_dadda_cska12_nand_8_11));
  fa fa_s_dadda_cska12_fa97_out(.a(s_dadda_cska12_fa96_or0[0]), .b(s_dadda_cska12_nand_8_11[0]), .cin(s_dadda_cska12_fa63_xor1[0]), .fa_xor1(s_dadda_cska12_fa97_xor1), .fa_or0(s_dadda_cska12_fa97_or0));
  and_gate and_gate_s_dadda_cska12_and_10_10(.a(a[10]), .b(b[10]), .out(s_dadda_cska12_and_10_10));
  nand_gate nand_gate_s_dadda_cska12_nand_9_11(.a(a[9]), .b(b[11]), .out(s_dadda_cska12_nand_9_11));
  fa fa_s_dadda_cska12_fa98_out(.a(s_dadda_cska12_fa97_or0[0]), .b(s_dadda_cska12_and_10_10[0]), .cin(s_dadda_cska12_nand_9_11[0]), .fa_xor1(s_dadda_cska12_fa98_xor1), .fa_or0(s_dadda_cska12_fa98_or0));
  nand_gate nand_gate_s_dadda_cska12_nand_11_10(.a(a[11]), .b(b[10]), .out(s_dadda_cska12_nand_11_10));
  fa fa_s_dadda_cska12_fa99_out(.a(s_dadda_cska12_fa98_or0[0]), .b(s_dadda_cska12_fa80_or0[0]), .cin(s_dadda_cska12_nand_11_10[0]), .fa_xor1(s_dadda_cska12_fa99_xor1), .fa_or0(s_dadda_cska12_fa99_or0));
  and_gate and_gate_s_dadda_cska12_and_0_0(.a(a[0]), .b(b[0]), .out(s_dadda_cska12_and_0_0));
  and_gate and_gate_s_dadda_cska12_and_1_0(.a(a[1]), .b(b[0]), .out(s_dadda_cska12_and_1_0));
  and_gate and_gate_s_dadda_cska12_and_0_2(.a(a[0]), .b(b[2]), .out(s_dadda_cska12_and_0_2));
  nand_gate nand_gate_s_dadda_cska12_nand_10_11(.a(a[10]), .b(b[11]), .out(s_dadda_cska12_nand_10_11));
  and_gate and_gate_s_dadda_cska12_and_0_1(.a(a[0]), .b(b[1]), .out(s_dadda_cska12_and_0_1));
  and_gate and_gate_s_dadda_cska12_and_11_11(.a(a[11]), .b(b[11]), .out(s_dadda_cska12_and_11_11));
  assign s_dadda_cska12_u_cska22_a[0] = s_dadda_cska12_and_1_0[0];
  assign s_dadda_cska12_u_cska22_a[1] = s_dadda_cska12_and_0_2[0];
  assign s_dadda_cska12_u_cska22_a[2] = s_dadda_cska12_ha8_xor0[0];
  assign s_dadda_cska12_u_cska22_a[3] = s_dadda_cska12_fa64_xor1[0];
  assign s_dadda_cska12_u_cska22_a[4] = s_dadda_cska12_fa65_xor1[0];
  assign s_dadda_cska12_u_cska22_a[5] = s_dadda_cska12_fa66_xor1[0];
  assign s_dadda_cska12_u_cska22_a[6] = s_dadda_cska12_fa67_xor1[0];
  assign s_dadda_cska12_u_cska22_a[7] = s_dadda_cska12_fa68_xor1[0];
  assign s_dadda_cska12_u_cska22_a[8] = s_dadda_cska12_fa69_xor1[0];
  assign s_dadda_cska12_u_cska22_a[9] = s_dadda_cska12_fa70_xor1[0];
  assign s_dadda_cska12_u_cska22_a[10] = s_dadda_cska12_fa71_xor1[0];
  assign s_dadda_cska12_u_cska22_a[11] = s_dadda_cska12_fa72_xor1[0];
  assign s_dadda_cska12_u_cska22_a[12] = s_dadda_cska12_fa73_xor1[0];
  assign s_dadda_cska12_u_cska22_a[13] = s_dadda_cska12_fa74_xor1[0];
  assign s_dadda_cska12_u_cska22_a[14] = s_dadda_cska12_fa75_xor1[0];
  assign s_dadda_cska12_u_cska22_a[15] = s_dadda_cska12_fa76_xor1[0];
  assign s_dadda_cska12_u_cska22_a[16] = s_dadda_cska12_fa77_xor1[0];
  assign s_dadda_cska12_u_cska22_a[17] = s_dadda_cska12_fa78_xor1[0];
  assign s_dadda_cska12_u_cska22_a[18] = s_dadda_cska12_fa79_xor1[0];
  assign s_dadda_cska12_u_cska22_a[19] = s_dadda_cska12_fa80_xor1[0];
  assign s_dadda_cska12_u_cska22_a[20] = s_dadda_cska12_nand_10_11[0];
  assign s_dadda_cska12_u_cska22_a[21] = s_dadda_cska12_fa99_or0[0];
  assign s_dadda_cska12_u_cska22_b[0] = s_dadda_cska12_and_0_1[0];
  assign s_dadda_cska12_u_cska22_b[1] = s_dadda_cska12_ha9_xor0[0];
  assign s_dadda_cska12_u_cska22_b[2] = s_dadda_cska12_fa81_xor1[0];
  assign s_dadda_cska12_u_cska22_b[3] = s_dadda_cska12_fa82_xor1[0];
  assign s_dadda_cska12_u_cska22_b[4] = s_dadda_cska12_fa83_xor1[0];
  assign s_dadda_cska12_u_cska22_b[5] = s_dadda_cska12_fa84_xor1[0];
  assign s_dadda_cska12_u_cska22_b[6] = s_dadda_cska12_fa85_xor1[0];
  assign s_dadda_cska12_u_cska22_b[7] = s_dadda_cska12_fa86_xor1[0];
  assign s_dadda_cska12_u_cska22_b[8] = s_dadda_cska12_fa87_xor1[0];
  assign s_dadda_cska12_u_cska22_b[9] = s_dadda_cska12_fa88_xor1[0];
  assign s_dadda_cska12_u_cska22_b[10] = s_dadda_cska12_fa89_xor1[0];
  assign s_dadda_cska12_u_cska22_b[11] = s_dadda_cska12_fa90_xor1[0];
  assign s_dadda_cska12_u_cska22_b[12] = s_dadda_cska12_fa91_xor1[0];
  assign s_dadda_cska12_u_cska22_b[13] = s_dadda_cska12_fa92_xor1[0];
  assign s_dadda_cska12_u_cska22_b[14] = s_dadda_cska12_fa93_xor1[0];
  assign s_dadda_cska12_u_cska22_b[15] = s_dadda_cska12_fa94_xor1[0];
  assign s_dadda_cska12_u_cska22_b[16] = s_dadda_cska12_fa95_xor1[0];
  assign s_dadda_cska12_u_cska22_b[17] = s_dadda_cska12_fa96_xor1[0];
  assign s_dadda_cska12_u_cska22_b[18] = s_dadda_cska12_fa97_xor1[0];
  assign s_dadda_cska12_u_cska22_b[19] = s_dadda_cska12_fa98_xor1[0];
  assign s_dadda_cska12_u_cska22_b[20] = s_dadda_cska12_fa99_xor1[0];
  assign s_dadda_cska12_u_cska22_b[21] = s_dadda_cska12_and_11_11[0];
  u_cska22 u_cska22_s_dadda_cska12_u_cska22_out(.a(s_dadda_cska12_u_cska22_a), .b(s_dadda_cska12_u_cska22_b), .u_cska22_out(s_dadda_cska12_u_cska22_out));
  not_gate not_gate_s_dadda_cska12_xor0(.a(s_dadda_cska12_u_cska22_out[22]), .out(s_dadda_cska12_xor0));

  assign s_dadda_cska12_out[0] = s_dadda_cska12_and_0_0[0];
  assign s_dadda_cska12_out[1] = s_dadda_cska12_u_cska22_out[0];
  assign s_dadda_cska12_out[2] = s_dadda_cska12_u_cska22_out[1];
  assign s_dadda_cska12_out[3] = s_dadda_cska12_u_cska22_out[2];
  assign s_dadda_cska12_out[4] = s_dadda_cska12_u_cska22_out[3];
  assign s_dadda_cska12_out[5] = s_dadda_cska12_u_cska22_out[4];
  assign s_dadda_cska12_out[6] = s_dadda_cska12_u_cska22_out[5];
  assign s_dadda_cska12_out[7] = s_dadda_cska12_u_cska22_out[6];
  assign s_dadda_cska12_out[8] = s_dadda_cska12_u_cska22_out[7];
  assign s_dadda_cska12_out[9] = s_dadda_cska12_u_cska22_out[8];
  assign s_dadda_cska12_out[10] = s_dadda_cska12_u_cska22_out[9];
  assign s_dadda_cska12_out[11] = s_dadda_cska12_u_cska22_out[10];
  assign s_dadda_cska12_out[12] = s_dadda_cska12_u_cska22_out[11];
  assign s_dadda_cska12_out[13] = s_dadda_cska12_u_cska22_out[12];
  assign s_dadda_cska12_out[14] = s_dadda_cska12_u_cska22_out[13];
  assign s_dadda_cska12_out[15] = s_dadda_cska12_u_cska22_out[14];
  assign s_dadda_cska12_out[16] = s_dadda_cska12_u_cska22_out[15];
  assign s_dadda_cska12_out[17] = s_dadda_cska12_u_cska22_out[16];
  assign s_dadda_cska12_out[18] = s_dadda_cska12_u_cska22_out[17];
  assign s_dadda_cska12_out[19] = s_dadda_cska12_u_cska22_out[18];
  assign s_dadda_cska12_out[20] = s_dadda_cska12_u_cska22_out[19];
  assign s_dadda_cska12_out[21] = s_dadda_cska12_u_cska22_out[20];
  assign s_dadda_cska12_out[22] = s_dadda_cska12_u_cska22_out[21];
  assign s_dadda_cska12_out[23] = s_dadda_cska12_xor0[0];
endmodule