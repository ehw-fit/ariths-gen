module s_CSAwallace_cska12(input [11:0] a, input [11:0] b, output [23:0] s_CSAwallace_cska12_out);
  wire s_CSAwallace_cska12_and_0_0;
  wire s_CSAwallace_cska12_and_1_0;
  wire s_CSAwallace_cska12_and_2_0;
  wire s_CSAwallace_cska12_and_3_0;
  wire s_CSAwallace_cska12_and_4_0;
  wire s_CSAwallace_cska12_and_5_0;
  wire s_CSAwallace_cska12_and_6_0;
  wire s_CSAwallace_cska12_and_7_0;
  wire s_CSAwallace_cska12_and_8_0;
  wire s_CSAwallace_cska12_and_9_0;
  wire s_CSAwallace_cska12_and_10_0;
  wire s_CSAwallace_cska12_nand_11_0;
  wire s_CSAwallace_cska12_and_0_1;
  wire s_CSAwallace_cska12_and_1_1;
  wire s_CSAwallace_cska12_and_2_1;
  wire s_CSAwallace_cska12_and_3_1;
  wire s_CSAwallace_cska12_and_4_1;
  wire s_CSAwallace_cska12_and_5_1;
  wire s_CSAwallace_cska12_and_6_1;
  wire s_CSAwallace_cska12_and_7_1;
  wire s_CSAwallace_cska12_and_8_1;
  wire s_CSAwallace_cska12_and_9_1;
  wire s_CSAwallace_cska12_and_10_1;
  wire s_CSAwallace_cska12_nand_11_1;
  wire s_CSAwallace_cska12_and_0_2;
  wire s_CSAwallace_cska12_and_1_2;
  wire s_CSAwallace_cska12_and_2_2;
  wire s_CSAwallace_cska12_and_3_2;
  wire s_CSAwallace_cska12_and_4_2;
  wire s_CSAwallace_cska12_and_5_2;
  wire s_CSAwallace_cska12_and_6_2;
  wire s_CSAwallace_cska12_and_7_2;
  wire s_CSAwallace_cska12_and_8_2;
  wire s_CSAwallace_cska12_and_9_2;
  wire s_CSAwallace_cska12_and_10_2;
  wire s_CSAwallace_cska12_nand_11_2;
  wire s_CSAwallace_cska12_and_0_3;
  wire s_CSAwallace_cska12_and_1_3;
  wire s_CSAwallace_cska12_and_2_3;
  wire s_CSAwallace_cska12_and_3_3;
  wire s_CSAwallace_cska12_and_4_3;
  wire s_CSAwallace_cska12_and_5_3;
  wire s_CSAwallace_cska12_and_6_3;
  wire s_CSAwallace_cska12_and_7_3;
  wire s_CSAwallace_cska12_and_8_3;
  wire s_CSAwallace_cska12_and_9_3;
  wire s_CSAwallace_cska12_and_10_3;
  wire s_CSAwallace_cska12_nand_11_3;
  wire s_CSAwallace_cska12_and_0_4;
  wire s_CSAwallace_cska12_and_1_4;
  wire s_CSAwallace_cska12_and_2_4;
  wire s_CSAwallace_cska12_and_3_4;
  wire s_CSAwallace_cska12_and_4_4;
  wire s_CSAwallace_cska12_and_5_4;
  wire s_CSAwallace_cska12_and_6_4;
  wire s_CSAwallace_cska12_and_7_4;
  wire s_CSAwallace_cska12_and_8_4;
  wire s_CSAwallace_cska12_and_9_4;
  wire s_CSAwallace_cska12_and_10_4;
  wire s_CSAwallace_cska12_nand_11_4;
  wire s_CSAwallace_cska12_and_0_5;
  wire s_CSAwallace_cska12_and_1_5;
  wire s_CSAwallace_cska12_and_2_5;
  wire s_CSAwallace_cska12_and_3_5;
  wire s_CSAwallace_cska12_and_4_5;
  wire s_CSAwallace_cska12_and_5_5;
  wire s_CSAwallace_cska12_and_6_5;
  wire s_CSAwallace_cska12_and_7_5;
  wire s_CSAwallace_cska12_and_8_5;
  wire s_CSAwallace_cska12_and_9_5;
  wire s_CSAwallace_cska12_and_10_5;
  wire s_CSAwallace_cska12_nand_11_5;
  wire s_CSAwallace_cska12_and_0_6;
  wire s_CSAwallace_cska12_and_1_6;
  wire s_CSAwallace_cska12_and_2_6;
  wire s_CSAwallace_cska12_and_3_6;
  wire s_CSAwallace_cska12_and_4_6;
  wire s_CSAwallace_cska12_and_5_6;
  wire s_CSAwallace_cska12_and_6_6;
  wire s_CSAwallace_cska12_and_7_6;
  wire s_CSAwallace_cska12_and_8_6;
  wire s_CSAwallace_cska12_and_9_6;
  wire s_CSAwallace_cska12_and_10_6;
  wire s_CSAwallace_cska12_nand_11_6;
  wire s_CSAwallace_cska12_and_0_7;
  wire s_CSAwallace_cska12_and_1_7;
  wire s_CSAwallace_cska12_and_2_7;
  wire s_CSAwallace_cska12_and_3_7;
  wire s_CSAwallace_cska12_and_4_7;
  wire s_CSAwallace_cska12_and_5_7;
  wire s_CSAwallace_cska12_and_6_7;
  wire s_CSAwallace_cska12_and_7_7;
  wire s_CSAwallace_cska12_and_8_7;
  wire s_CSAwallace_cska12_and_9_7;
  wire s_CSAwallace_cska12_and_10_7;
  wire s_CSAwallace_cska12_nand_11_7;
  wire s_CSAwallace_cska12_and_0_8;
  wire s_CSAwallace_cska12_and_1_8;
  wire s_CSAwallace_cska12_and_2_8;
  wire s_CSAwallace_cska12_and_3_8;
  wire s_CSAwallace_cska12_and_4_8;
  wire s_CSAwallace_cska12_and_5_8;
  wire s_CSAwallace_cska12_and_6_8;
  wire s_CSAwallace_cska12_and_7_8;
  wire s_CSAwallace_cska12_and_8_8;
  wire s_CSAwallace_cska12_and_9_8;
  wire s_CSAwallace_cska12_and_10_8;
  wire s_CSAwallace_cska12_nand_11_8;
  wire s_CSAwallace_cska12_and_0_9;
  wire s_CSAwallace_cska12_and_1_9;
  wire s_CSAwallace_cska12_and_2_9;
  wire s_CSAwallace_cska12_and_3_9;
  wire s_CSAwallace_cska12_and_4_9;
  wire s_CSAwallace_cska12_and_5_9;
  wire s_CSAwallace_cska12_and_6_9;
  wire s_CSAwallace_cska12_and_7_9;
  wire s_CSAwallace_cska12_and_8_9;
  wire s_CSAwallace_cska12_and_9_9;
  wire s_CSAwallace_cska12_and_10_9;
  wire s_CSAwallace_cska12_nand_11_9;
  wire s_CSAwallace_cska12_and_0_10;
  wire s_CSAwallace_cska12_and_1_10;
  wire s_CSAwallace_cska12_and_2_10;
  wire s_CSAwallace_cska12_and_3_10;
  wire s_CSAwallace_cska12_and_4_10;
  wire s_CSAwallace_cska12_and_5_10;
  wire s_CSAwallace_cska12_and_6_10;
  wire s_CSAwallace_cska12_and_7_10;
  wire s_CSAwallace_cska12_and_8_10;
  wire s_CSAwallace_cska12_and_9_10;
  wire s_CSAwallace_cska12_and_10_10;
  wire s_CSAwallace_cska12_nand_11_10;
  wire s_CSAwallace_cska12_nand_0_11;
  wire s_CSAwallace_cska12_nand_1_11;
  wire s_CSAwallace_cska12_nand_2_11;
  wire s_CSAwallace_cska12_nand_3_11;
  wire s_CSAwallace_cska12_nand_4_11;
  wire s_CSAwallace_cska12_nand_5_11;
  wire s_CSAwallace_cska12_nand_6_11;
  wire s_CSAwallace_cska12_nand_7_11;
  wire s_CSAwallace_cska12_nand_8_11;
  wire s_CSAwallace_cska12_nand_9_11;
  wire s_CSAwallace_cska12_nand_10_11;
  wire s_CSAwallace_cska12_and_11_11;
  wire s_CSAwallace_cska12_csa0_csa_component_fa1_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa1_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa2_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa2_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa2_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa2_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa2_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa3_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa3_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa3_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa3_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa3_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa4_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa4_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa4_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa4_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa4_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa5_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa5_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa5_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa5_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa5_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa6_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa6_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa6_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa6_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa6_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa7_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa7_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa7_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa7_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa7_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa8_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa8_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa8_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa8_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa8_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa9_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa9_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa9_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa9_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa9_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa10_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa10_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa10_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa0_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa0_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa4_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa4_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa5_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa5_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa5_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa5_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa5_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa6_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa6_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa6_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa6_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa6_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa7_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa7_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa7_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa7_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa7_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa8_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa8_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa8_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa8_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa8_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa9_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa9_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa9_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa9_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa9_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa10_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa10_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa10_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa12_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa13_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa13_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa13_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa13_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa13_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa14_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa14_and0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa14_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa14_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa14_or0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa15_xor0;
  wire s_CSAwallace_cska12_csa1_csa_component_fa15_xor1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa15_and1;
  wire s_CSAwallace_cska12_csa1_csa_component_fa15_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa7_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa7_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa8_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa8_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa8_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa8_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa8_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa9_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa9_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa9_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa9_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa9_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa10_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa10_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa10_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa12_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa13_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa13_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa13_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa13_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa13_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa14_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa14_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa14_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa14_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa14_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa15_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa15_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa15_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa15_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa15_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa16_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa16_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa16_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa16_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa16_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa17_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa17_and0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa17_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa17_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa17_or0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa18_xor0;
  wire s_CSAwallace_cska12_csa2_csa_component_fa18_xor1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa18_and1;
  wire s_CSAwallace_cska12_csa2_csa_component_fa18_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa12_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa13_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa13_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa13_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa13_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa13_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa14_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa14_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa14_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa14_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa14_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa15_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa15_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa15_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa15_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa15_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa16_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa16_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa16_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa16_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa16_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa17_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa17_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa17_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa17_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa17_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa18_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa18_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa18_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa18_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa18_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa19_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa19_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa19_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa19_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa19_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa20_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa20_and0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa20_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa20_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa20_or0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa21_xor0;
  wire s_CSAwallace_cska12_csa3_csa_component_fa21_xor1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa21_and1;
  wire s_CSAwallace_cska12_csa3_csa_component_fa21_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa2_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa2_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa3_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa3_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa3_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa3_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa3_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa4_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa4_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa4_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa4_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa4_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa5_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa5_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa5_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa5_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa5_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa6_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa6_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa6_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa6_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa6_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa7_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa7_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa7_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa7_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa7_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa8_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa8_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa8_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa8_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa8_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa9_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa9_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa9_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa9_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa9_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa10_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa10_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa10_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa12_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa13_xor0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa13_and0;
  wire s_CSAwallace_cska12_csa4_csa_component_fa13_xor1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa13_and1;
  wire s_CSAwallace_cska12_csa4_csa_component_fa13_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa6_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa6_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa7_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa7_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa8_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa8_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa8_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa8_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa8_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa9_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa9_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa9_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa9_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa9_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa10_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa10_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa10_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa12_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa13_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa13_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa13_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa13_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa13_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa14_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa14_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa14_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa14_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa14_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa15_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa15_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa15_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa15_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa15_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa16_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa16_and0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa16_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa16_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa16_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa17_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa17_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa17_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa17_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa18_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa18_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa18_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa18_or0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa19_xor0;
  wire s_CSAwallace_cska12_csa5_csa_component_fa19_xor1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa19_and1;
  wire s_CSAwallace_cska12_csa5_csa_component_fa19_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa3_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa3_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa4_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa4_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa5_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa5_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa5_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa5_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa5_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa6_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa6_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa6_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa6_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa6_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa7_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa7_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa7_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa7_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa7_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa8_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa8_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa8_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa8_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa8_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa9_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa9_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa9_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa9_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa9_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa10_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa10_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa10_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa12_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa13_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa13_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa13_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa13_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa13_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa14_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa14_and0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa14_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa14_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa14_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa15_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa15_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa15_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa15_or0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa16_xor0;
  wire s_CSAwallace_cska12_csa6_csa_component_fa16_xor1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa16_and1;
  wire s_CSAwallace_cska12_csa6_csa_component_fa16_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa9_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa9_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa12_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa13_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa13_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa13_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa13_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa13_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa14_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa14_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa14_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa14_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa14_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa15_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa15_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa15_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa15_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa15_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa16_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa16_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa16_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa16_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa16_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa17_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa17_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa17_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa17_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa17_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa18_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa18_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa18_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa18_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa18_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa19_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa19_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa19_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa19_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa19_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa20_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa20_and0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa20_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa20_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa20_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa21_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa21_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa21_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa21_or0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa22_xor0;
  wire s_CSAwallace_cska12_csa7_csa_component_fa22_xor1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa22_and1;
  wire s_CSAwallace_cska12_csa7_csa_component_fa22_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa4_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa4_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa5_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa5_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa6_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa6_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa7_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa7_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa7_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa7_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa7_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa8_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa8_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa8_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa8_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa8_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa9_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa9_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa9_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa9_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa9_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa10_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa10_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa10_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa12_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa13_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa13_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa13_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa13_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa13_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa14_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa14_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa14_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa14_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa14_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa15_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa15_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa15_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa15_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa15_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa16_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa16_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa16_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa16_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa16_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa17_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa17_and0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa17_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa17_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa17_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa18_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa18_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa18_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa18_or0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa19_xor0;
  wire s_CSAwallace_cska12_csa8_csa_component_fa19_xor1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa19_and1;
  wire s_CSAwallace_cska12_csa8_csa_component_fa19_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa5_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa5_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa6_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa6_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa7_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa7_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa8_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa8_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa9_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa9_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa10_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa10_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa10_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa10_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa10_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa11_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa11_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa11_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa11_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa11_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa12_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa12_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa12_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa12_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa12_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa13_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa13_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa13_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa13_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa13_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa14_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa14_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa14_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa14_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa14_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa15_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa15_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa15_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa15_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa15_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa16_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa16_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa16_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa16_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa16_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa17_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa17_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa17_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa17_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa17_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa18_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa18_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa18_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa18_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa18_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa19_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa19_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa19_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa19_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa19_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa20_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa20_and0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa20_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa20_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa20_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa21_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa21_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa21_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa21_or0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa22_xor0;
  wire s_CSAwallace_cska12_csa9_csa_component_fa22_xor1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa22_and1;
  wire s_CSAwallace_cska12_csa9_csa_component_fa22_or0;
  wire s_CSAwallace_cska12_u_cska24_and_propagate00;
  wire s_CSAwallace_cska12_u_cska24_and_propagate01;
  wire s_CSAwallace_cska12_u_cska24_and_propagate02;
  wire s_CSAwallace_cska12_u_cska24_mux2to10_not0;
  wire s_CSAwallace_cska12_u_cska24_xor6;
  wire s_CSAwallace_cska12_u_cska24_fa5_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa5_and0;
  wire s_CSAwallace_cska12_u_cska24_xor7;
  wire s_CSAwallace_cska12_u_cska24_fa6_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa6_and0;
  wire s_CSAwallace_cska12_u_cska24_fa6_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa6_and1;
  wire s_CSAwallace_cska12_u_cska24_fa6_or0;
  wire s_CSAwallace_cska12_u_cska24_and_propagate13;
  wire s_CSAwallace_cska12_u_cska24_and_propagate14;
  wire s_CSAwallace_cska12_u_cska24_and_propagate15;
  wire s_CSAwallace_cska12_u_cska24_mux2to11_not0;
  wire s_CSAwallace_cska12_u_cska24_mux2to11_and1;
  wire s_CSAwallace_cska12_u_cska24_xor8;
  wire s_CSAwallace_cska12_u_cska24_fa7_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa7_and0;
  wire s_CSAwallace_cska12_u_cska24_fa7_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa7_and1;
  wire s_CSAwallace_cska12_u_cska24_fa7_or0;
  wire s_CSAwallace_cska12_u_cska24_xor9;
  wire s_CSAwallace_cska12_u_cska24_fa8_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa8_and0;
  wire s_CSAwallace_cska12_u_cska24_fa8_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa8_and1;
  wire s_CSAwallace_cska12_u_cska24_fa8_or0;
  wire s_CSAwallace_cska12_u_cska24_xor10;
  wire s_CSAwallace_cska12_u_cska24_fa9_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa9_and0;
  wire s_CSAwallace_cska12_u_cska24_fa9_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa9_and1;
  wire s_CSAwallace_cska12_u_cska24_fa9_or0;
  wire s_CSAwallace_cska12_u_cska24_xor11;
  wire s_CSAwallace_cska12_u_cska24_fa10_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa10_and0;
  wire s_CSAwallace_cska12_u_cska24_fa10_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa10_and1;
  wire s_CSAwallace_cska12_u_cska24_fa10_or0;
  wire s_CSAwallace_cska12_u_cska24_and_propagate26;
  wire s_CSAwallace_cska12_u_cska24_and_propagate27;
  wire s_CSAwallace_cska12_u_cska24_and_propagate28;
  wire s_CSAwallace_cska12_u_cska24_mux2to12_and0;
  wire s_CSAwallace_cska12_u_cska24_mux2to12_not0;
  wire s_CSAwallace_cska12_u_cska24_mux2to12_and1;
  wire s_CSAwallace_cska12_u_cska24_mux2to12_xor0;
  wire s_CSAwallace_cska12_u_cska24_xor12;
  wire s_CSAwallace_cska12_u_cska24_fa11_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa11_and0;
  wire s_CSAwallace_cska12_u_cska24_fa11_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa11_and1;
  wire s_CSAwallace_cska12_u_cska24_fa11_or0;
  wire s_CSAwallace_cska12_u_cska24_xor13;
  wire s_CSAwallace_cska12_u_cska24_fa12_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa12_and0;
  wire s_CSAwallace_cska12_u_cska24_fa12_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa12_and1;
  wire s_CSAwallace_cska12_u_cska24_fa12_or0;
  wire s_CSAwallace_cska12_u_cska24_xor14;
  wire s_CSAwallace_cska12_u_cska24_fa13_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa13_and0;
  wire s_CSAwallace_cska12_u_cska24_fa13_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa13_and1;
  wire s_CSAwallace_cska12_u_cska24_fa13_or0;
  wire s_CSAwallace_cska12_u_cska24_xor15;
  wire s_CSAwallace_cska12_u_cska24_fa14_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa14_and0;
  wire s_CSAwallace_cska12_u_cska24_fa14_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa14_and1;
  wire s_CSAwallace_cska12_u_cska24_fa14_or0;
  wire s_CSAwallace_cska12_u_cska24_and_propagate39;
  wire s_CSAwallace_cska12_u_cska24_and_propagate310;
  wire s_CSAwallace_cska12_u_cska24_and_propagate311;
  wire s_CSAwallace_cska12_u_cska24_mux2to13_and0;
  wire s_CSAwallace_cska12_u_cska24_mux2to13_not0;
  wire s_CSAwallace_cska12_u_cska24_mux2to13_and1;
  wire s_CSAwallace_cska12_u_cska24_mux2to13_xor0;
  wire s_CSAwallace_cska12_u_cska24_xor16;
  wire s_CSAwallace_cska12_u_cska24_fa15_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa15_and0;
  wire s_CSAwallace_cska12_u_cska24_fa15_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa15_and1;
  wire s_CSAwallace_cska12_u_cska24_fa15_or0;
  wire s_CSAwallace_cska12_u_cska24_xor17;
  wire s_CSAwallace_cska12_u_cska24_fa16_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa16_and0;
  wire s_CSAwallace_cska12_u_cska24_fa16_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa16_and1;
  wire s_CSAwallace_cska12_u_cska24_fa16_or0;
  wire s_CSAwallace_cska12_u_cska24_xor18;
  wire s_CSAwallace_cska12_u_cska24_fa17_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa17_and0;
  wire s_CSAwallace_cska12_u_cska24_fa17_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa17_and1;
  wire s_CSAwallace_cska12_u_cska24_fa17_or0;
  wire s_CSAwallace_cska12_u_cska24_xor19;
  wire s_CSAwallace_cska12_u_cska24_fa18_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa18_and0;
  wire s_CSAwallace_cska12_u_cska24_fa18_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa18_and1;
  wire s_CSAwallace_cska12_u_cska24_fa18_or0;
  wire s_CSAwallace_cska12_u_cska24_and_propagate412;
  wire s_CSAwallace_cska12_u_cska24_and_propagate413;
  wire s_CSAwallace_cska12_u_cska24_and_propagate414;
  wire s_CSAwallace_cska12_u_cska24_mux2to14_and0;
  wire s_CSAwallace_cska12_u_cska24_mux2to14_not0;
  wire s_CSAwallace_cska12_u_cska24_mux2to14_and1;
  wire s_CSAwallace_cska12_u_cska24_mux2to14_xor0;
  wire s_CSAwallace_cska12_u_cska24_xor20;
  wire s_CSAwallace_cska12_u_cska24_fa19_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa19_and0;
  wire s_CSAwallace_cska12_u_cska24_fa19_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa19_and1;
  wire s_CSAwallace_cska12_u_cska24_fa19_or0;
  wire s_CSAwallace_cska12_u_cska24_xor21;
  wire s_CSAwallace_cska12_u_cska24_fa20_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa20_and0;
  wire s_CSAwallace_cska12_u_cska24_fa20_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa20_and1;
  wire s_CSAwallace_cska12_u_cska24_fa20_or0;
  wire s_CSAwallace_cska12_u_cska24_xor22;
  wire s_CSAwallace_cska12_u_cska24_fa21_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa21_and0;
  wire s_CSAwallace_cska12_u_cska24_fa21_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa21_and1;
  wire s_CSAwallace_cska12_u_cska24_fa21_or0;
  wire s_CSAwallace_cska12_u_cska24_xor23;
  wire s_CSAwallace_cska12_u_cska24_fa22_xor0;
  wire s_CSAwallace_cska12_u_cska24_fa22_and0;
  wire s_CSAwallace_cska12_u_cska24_fa22_xor1;
  wire s_CSAwallace_cska12_u_cska24_fa22_and1;
  wire s_CSAwallace_cska12_u_cska24_fa22_or0;
  wire s_CSAwallace_cska12_u_cska24_and_propagate515;
  wire s_CSAwallace_cska12_u_cska24_and_propagate516;
  wire s_CSAwallace_cska12_u_cska24_and_propagate517;
  wire s_CSAwallace_cska12_u_cska24_mux2to15_and0;
  wire s_CSAwallace_cska12_u_cska24_mux2to15_not0;
  wire s_CSAwallace_cska12_u_cska24_mux2to15_and1;
  wire s_CSAwallace_cska12_u_cska24_mux2to15_xor0;
  wire s_CSAwallace_cska12_xor0;

  assign s_CSAwallace_cska12_and_0_0 = a[0] & b[0];
  assign s_CSAwallace_cska12_and_1_0 = a[1] & b[0];
  assign s_CSAwallace_cska12_and_2_0 = a[2] & b[0];
  assign s_CSAwallace_cska12_and_3_0 = a[3] & b[0];
  assign s_CSAwallace_cska12_and_4_0 = a[4] & b[0];
  assign s_CSAwallace_cska12_and_5_0 = a[5] & b[0];
  assign s_CSAwallace_cska12_and_6_0 = a[6] & b[0];
  assign s_CSAwallace_cska12_and_7_0 = a[7] & b[0];
  assign s_CSAwallace_cska12_and_8_0 = a[8] & b[0];
  assign s_CSAwallace_cska12_and_9_0 = a[9] & b[0];
  assign s_CSAwallace_cska12_and_10_0 = a[10] & b[0];
  assign s_CSAwallace_cska12_nand_11_0 = ~(a[11] & b[0]);
  assign s_CSAwallace_cska12_and_0_1 = a[0] & b[1];
  assign s_CSAwallace_cska12_and_1_1 = a[1] & b[1];
  assign s_CSAwallace_cska12_and_2_1 = a[2] & b[1];
  assign s_CSAwallace_cska12_and_3_1 = a[3] & b[1];
  assign s_CSAwallace_cska12_and_4_1 = a[4] & b[1];
  assign s_CSAwallace_cska12_and_5_1 = a[5] & b[1];
  assign s_CSAwallace_cska12_and_6_1 = a[6] & b[1];
  assign s_CSAwallace_cska12_and_7_1 = a[7] & b[1];
  assign s_CSAwallace_cska12_and_8_1 = a[8] & b[1];
  assign s_CSAwallace_cska12_and_9_1 = a[9] & b[1];
  assign s_CSAwallace_cska12_and_10_1 = a[10] & b[1];
  assign s_CSAwallace_cska12_nand_11_1 = ~(a[11] & b[1]);
  assign s_CSAwallace_cska12_and_0_2 = a[0] & b[2];
  assign s_CSAwallace_cska12_and_1_2 = a[1] & b[2];
  assign s_CSAwallace_cska12_and_2_2 = a[2] & b[2];
  assign s_CSAwallace_cska12_and_3_2 = a[3] & b[2];
  assign s_CSAwallace_cska12_and_4_2 = a[4] & b[2];
  assign s_CSAwallace_cska12_and_5_2 = a[5] & b[2];
  assign s_CSAwallace_cska12_and_6_2 = a[6] & b[2];
  assign s_CSAwallace_cska12_and_7_2 = a[7] & b[2];
  assign s_CSAwallace_cska12_and_8_2 = a[8] & b[2];
  assign s_CSAwallace_cska12_and_9_2 = a[9] & b[2];
  assign s_CSAwallace_cska12_and_10_2 = a[10] & b[2];
  assign s_CSAwallace_cska12_nand_11_2 = ~(a[11] & b[2]);
  assign s_CSAwallace_cska12_and_0_3 = a[0] & b[3];
  assign s_CSAwallace_cska12_and_1_3 = a[1] & b[3];
  assign s_CSAwallace_cska12_and_2_3 = a[2] & b[3];
  assign s_CSAwallace_cska12_and_3_3 = a[3] & b[3];
  assign s_CSAwallace_cska12_and_4_3 = a[4] & b[3];
  assign s_CSAwallace_cska12_and_5_3 = a[5] & b[3];
  assign s_CSAwallace_cska12_and_6_3 = a[6] & b[3];
  assign s_CSAwallace_cska12_and_7_3 = a[7] & b[3];
  assign s_CSAwallace_cska12_and_8_3 = a[8] & b[3];
  assign s_CSAwallace_cska12_and_9_3 = a[9] & b[3];
  assign s_CSAwallace_cska12_and_10_3 = a[10] & b[3];
  assign s_CSAwallace_cska12_nand_11_3 = ~(a[11] & b[3]);
  assign s_CSAwallace_cska12_and_0_4 = a[0] & b[4];
  assign s_CSAwallace_cska12_and_1_4 = a[1] & b[4];
  assign s_CSAwallace_cska12_and_2_4 = a[2] & b[4];
  assign s_CSAwallace_cska12_and_3_4 = a[3] & b[4];
  assign s_CSAwallace_cska12_and_4_4 = a[4] & b[4];
  assign s_CSAwallace_cska12_and_5_4 = a[5] & b[4];
  assign s_CSAwallace_cska12_and_6_4 = a[6] & b[4];
  assign s_CSAwallace_cska12_and_7_4 = a[7] & b[4];
  assign s_CSAwallace_cska12_and_8_4 = a[8] & b[4];
  assign s_CSAwallace_cska12_and_9_4 = a[9] & b[4];
  assign s_CSAwallace_cska12_and_10_4 = a[10] & b[4];
  assign s_CSAwallace_cska12_nand_11_4 = ~(a[11] & b[4]);
  assign s_CSAwallace_cska12_and_0_5 = a[0] & b[5];
  assign s_CSAwallace_cska12_and_1_5 = a[1] & b[5];
  assign s_CSAwallace_cska12_and_2_5 = a[2] & b[5];
  assign s_CSAwallace_cska12_and_3_5 = a[3] & b[5];
  assign s_CSAwallace_cska12_and_4_5 = a[4] & b[5];
  assign s_CSAwallace_cska12_and_5_5 = a[5] & b[5];
  assign s_CSAwallace_cska12_and_6_5 = a[6] & b[5];
  assign s_CSAwallace_cska12_and_7_5 = a[7] & b[5];
  assign s_CSAwallace_cska12_and_8_5 = a[8] & b[5];
  assign s_CSAwallace_cska12_and_9_5 = a[9] & b[5];
  assign s_CSAwallace_cska12_and_10_5 = a[10] & b[5];
  assign s_CSAwallace_cska12_nand_11_5 = ~(a[11] & b[5]);
  assign s_CSAwallace_cska12_and_0_6 = a[0] & b[6];
  assign s_CSAwallace_cska12_and_1_6 = a[1] & b[6];
  assign s_CSAwallace_cska12_and_2_6 = a[2] & b[6];
  assign s_CSAwallace_cska12_and_3_6 = a[3] & b[6];
  assign s_CSAwallace_cska12_and_4_6 = a[4] & b[6];
  assign s_CSAwallace_cska12_and_5_6 = a[5] & b[6];
  assign s_CSAwallace_cska12_and_6_6 = a[6] & b[6];
  assign s_CSAwallace_cska12_and_7_6 = a[7] & b[6];
  assign s_CSAwallace_cska12_and_8_6 = a[8] & b[6];
  assign s_CSAwallace_cska12_and_9_6 = a[9] & b[6];
  assign s_CSAwallace_cska12_and_10_6 = a[10] & b[6];
  assign s_CSAwallace_cska12_nand_11_6 = ~(a[11] & b[6]);
  assign s_CSAwallace_cska12_and_0_7 = a[0] & b[7];
  assign s_CSAwallace_cska12_and_1_7 = a[1] & b[7];
  assign s_CSAwallace_cska12_and_2_7 = a[2] & b[7];
  assign s_CSAwallace_cska12_and_3_7 = a[3] & b[7];
  assign s_CSAwallace_cska12_and_4_7 = a[4] & b[7];
  assign s_CSAwallace_cska12_and_5_7 = a[5] & b[7];
  assign s_CSAwallace_cska12_and_6_7 = a[6] & b[7];
  assign s_CSAwallace_cska12_and_7_7 = a[7] & b[7];
  assign s_CSAwallace_cska12_and_8_7 = a[8] & b[7];
  assign s_CSAwallace_cska12_and_9_7 = a[9] & b[7];
  assign s_CSAwallace_cska12_and_10_7 = a[10] & b[7];
  assign s_CSAwallace_cska12_nand_11_7 = ~(a[11] & b[7]);
  assign s_CSAwallace_cska12_and_0_8 = a[0] & b[8];
  assign s_CSAwallace_cska12_and_1_8 = a[1] & b[8];
  assign s_CSAwallace_cska12_and_2_8 = a[2] & b[8];
  assign s_CSAwallace_cska12_and_3_8 = a[3] & b[8];
  assign s_CSAwallace_cska12_and_4_8 = a[4] & b[8];
  assign s_CSAwallace_cska12_and_5_8 = a[5] & b[8];
  assign s_CSAwallace_cska12_and_6_8 = a[6] & b[8];
  assign s_CSAwallace_cska12_and_7_8 = a[7] & b[8];
  assign s_CSAwallace_cska12_and_8_8 = a[8] & b[8];
  assign s_CSAwallace_cska12_and_9_8 = a[9] & b[8];
  assign s_CSAwallace_cska12_and_10_8 = a[10] & b[8];
  assign s_CSAwallace_cska12_nand_11_8 = ~(a[11] & b[8]);
  assign s_CSAwallace_cska12_and_0_9 = a[0] & b[9];
  assign s_CSAwallace_cska12_and_1_9 = a[1] & b[9];
  assign s_CSAwallace_cska12_and_2_9 = a[2] & b[9];
  assign s_CSAwallace_cska12_and_3_9 = a[3] & b[9];
  assign s_CSAwallace_cska12_and_4_9 = a[4] & b[9];
  assign s_CSAwallace_cska12_and_5_9 = a[5] & b[9];
  assign s_CSAwallace_cska12_and_6_9 = a[6] & b[9];
  assign s_CSAwallace_cska12_and_7_9 = a[7] & b[9];
  assign s_CSAwallace_cska12_and_8_9 = a[8] & b[9];
  assign s_CSAwallace_cska12_and_9_9 = a[9] & b[9];
  assign s_CSAwallace_cska12_and_10_9 = a[10] & b[9];
  assign s_CSAwallace_cska12_nand_11_9 = ~(a[11] & b[9]);
  assign s_CSAwallace_cska12_and_0_10 = a[0] & b[10];
  assign s_CSAwallace_cska12_and_1_10 = a[1] & b[10];
  assign s_CSAwallace_cska12_and_2_10 = a[2] & b[10];
  assign s_CSAwallace_cska12_and_3_10 = a[3] & b[10];
  assign s_CSAwallace_cska12_and_4_10 = a[4] & b[10];
  assign s_CSAwallace_cska12_and_5_10 = a[5] & b[10];
  assign s_CSAwallace_cska12_and_6_10 = a[6] & b[10];
  assign s_CSAwallace_cska12_and_7_10 = a[7] & b[10];
  assign s_CSAwallace_cska12_and_8_10 = a[8] & b[10];
  assign s_CSAwallace_cska12_and_9_10 = a[9] & b[10];
  assign s_CSAwallace_cska12_and_10_10 = a[10] & b[10];
  assign s_CSAwallace_cska12_nand_11_10 = ~(a[11] & b[10]);
  assign s_CSAwallace_cska12_nand_0_11 = ~(a[0] & b[11]);
  assign s_CSAwallace_cska12_nand_1_11 = ~(a[1] & b[11]);
  assign s_CSAwallace_cska12_nand_2_11 = ~(a[2] & b[11]);
  assign s_CSAwallace_cska12_nand_3_11 = ~(a[3] & b[11]);
  assign s_CSAwallace_cska12_nand_4_11 = ~(a[4] & b[11]);
  assign s_CSAwallace_cska12_nand_5_11 = ~(a[5] & b[11]);
  assign s_CSAwallace_cska12_nand_6_11 = ~(a[6] & b[11]);
  assign s_CSAwallace_cska12_nand_7_11 = ~(a[7] & b[11]);
  assign s_CSAwallace_cska12_nand_8_11 = ~(a[8] & b[11]);
  assign s_CSAwallace_cska12_nand_9_11 = ~(a[9] & b[11]);
  assign s_CSAwallace_cska12_nand_10_11 = ~(a[10] & b[11]);
  assign s_CSAwallace_cska12_and_11_11 = a[11] & b[11];
  assign s_CSAwallace_cska12_csa0_csa_component_fa1_xor0 = s_CSAwallace_cska12_and_1_0 ^ s_CSAwallace_cska12_and_0_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa1_and0 = s_CSAwallace_cska12_and_1_0 & s_CSAwallace_cska12_and_0_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa2_xor0 = s_CSAwallace_cska12_and_2_0 ^ s_CSAwallace_cska12_and_1_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa2_and0 = s_CSAwallace_cska12_and_2_0 & s_CSAwallace_cska12_and_1_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa2_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa2_xor0 ^ s_CSAwallace_cska12_and_0_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa2_and1 = s_CSAwallace_cska12_csa0_csa_component_fa2_xor0 & s_CSAwallace_cska12_and_0_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa2_or0 = s_CSAwallace_cska12_csa0_csa_component_fa2_and0 | s_CSAwallace_cska12_csa0_csa_component_fa2_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa3_xor0 = s_CSAwallace_cska12_and_3_0 ^ s_CSAwallace_cska12_and_2_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa3_and0 = s_CSAwallace_cska12_and_3_0 & s_CSAwallace_cska12_and_2_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa3_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa3_xor0 ^ s_CSAwallace_cska12_and_1_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa3_and1 = s_CSAwallace_cska12_csa0_csa_component_fa3_xor0 & s_CSAwallace_cska12_and_1_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa3_or0 = s_CSAwallace_cska12_csa0_csa_component_fa3_and0 | s_CSAwallace_cska12_csa0_csa_component_fa3_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa4_xor0 = s_CSAwallace_cska12_and_4_0 ^ s_CSAwallace_cska12_and_3_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa4_and0 = s_CSAwallace_cska12_and_4_0 & s_CSAwallace_cska12_and_3_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa4_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa4_xor0 ^ s_CSAwallace_cska12_and_2_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa4_and1 = s_CSAwallace_cska12_csa0_csa_component_fa4_xor0 & s_CSAwallace_cska12_and_2_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa4_or0 = s_CSAwallace_cska12_csa0_csa_component_fa4_and0 | s_CSAwallace_cska12_csa0_csa_component_fa4_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa5_xor0 = s_CSAwallace_cska12_and_5_0 ^ s_CSAwallace_cska12_and_4_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa5_and0 = s_CSAwallace_cska12_and_5_0 & s_CSAwallace_cska12_and_4_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa5_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa5_xor0 ^ s_CSAwallace_cska12_and_3_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa5_and1 = s_CSAwallace_cska12_csa0_csa_component_fa5_xor0 & s_CSAwallace_cska12_and_3_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa5_or0 = s_CSAwallace_cska12_csa0_csa_component_fa5_and0 | s_CSAwallace_cska12_csa0_csa_component_fa5_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa6_xor0 = s_CSAwallace_cska12_and_6_0 ^ s_CSAwallace_cska12_and_5_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa6_and0 = s_CSAwallace_cska12_and_6_0 & s_CSAwallace_cska12_and_5_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa6_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa6_xor0 ^ s_CSAwallace_cska12_and_4_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa6_and1 = s_CSAwallace_cska12_csa0_csa_component_fa6_xor0 & s_CSAwallace_cska12_and_4_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa6_or0 = s_CSAwallace_cska12_csa0_csa_component_fa6_and0 | s_CSAwallace_cska12_csa0_csa_component_fa6_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa7_xor0 = s_CSAwallace_cska12_and_7_0 ^ s_CSAwallace_cska12_and_6_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa7_and0 = s_CSAwallace_cska12_and_7_0 & s_CSAwallace_cska12_and_6_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa7_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa7_xor0 ^ s_CSAwallace_cska12_and_5_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa7_and1 = s_CSAwallace_cska12_csa0_csa_component_fa7_xor0 & s_CSAwallace_cska12_and_5_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa7_or0 = s_CSAwallace_cska12_csa0_csa_component_fa7_and0 | s_CSAwallace_cska12_csa0_csa_component_fa7_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa8_xor0 = s_CSAwallace_cska12_and_8_0 ^ s_CSAwallace_cska12_and_7_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa8_and0 = s_CSAwallace_cska12_and_8_0 & s_CSAwallace_cska12_and_7_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa8_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa8_xor0 ^ s_CSAwallace_cska12_and_6_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa8_and1 = s_CSAwallace_cska12_csa0_csa_component_fa8_xor0 & s_CSAwallace_cska12_and_6_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa8_or0 = s_CSAwallace_cska12_csa0_csa_component_fa8_and0 | s_CSAwallace_cska12_csa0_csa_component_fa8_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa9_xor0 = s_CSAwallace_cska12_and_9_0 ^ s_CSAwallace_cska12_and_8_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa9_and0 = s_CSAwallace_cska12_and_9_0 & s_CSAwallace_cska12_and_8_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa9_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa9_xor0 ^ s_CSAwallace_cska12_and_7_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa9_and1 = s_CSAwallace_cska12_csa0_csa_component_fa9_xor0 & s_CSAwallace_cska12_and_7_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa9_or0 = s_CSAwallace_cska12_csa0_csa_component_fa9_and0 | s_CSAwallace_cska12_csa0_csa_component_fa9_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa10_xor0 = s_CSAwallace_cska12_and_10_0 ^ s_CSAwallace_cska12_and_9_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa10_and0 = s_CSAwallace_cska12_and_10_0 & s_CSAwallace_cska12_and_9_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa10_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa10_xor0 ^ s_CSAwallace_cska12_and_8_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa10_and1 = s_CSAwallace_cska12_csa0_csa_component_fa10_xor0 & s_CSAwallace_cska12_and_8_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa10_or0 = s_CSAwallace_cska12_csa0_csa_component_fa10_and0 | s_CSAwallace_cska12_csa0_csa_component_fa10_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa11_xor0 = s_CSAwallace_cska12_nand_11_0 ^ s_CSAwallace_cska12_and_10_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa11_and0 = s_CSAwallace_cska12_nand_11_0 & s_CSAwallace_cska12_and_10_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_and_9_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa11_and1 = s_CSAwallace_cska12_csa0_csa_component_fa11_xor0 & s_CSAwallace_cska12_and_9_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa11_or0 = s_CSAwallace_cska12_csa0_csa_component_fa11_and0 | s_CSAwallace_cska12_csa0_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa12_xor0 = ~s_CSAwallace_cska12_nand_11_1;
  assign s_CSAwallace_cska12_csa0_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa0_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_and_10_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa12_and1 = s_CSAwallace_cska12_csa0_csa_component_fa12_xor0 & s_CSAwallace_cska12_and_10_2;
  assign s_CSAwallace_cska12_csa0_csa_component_fa12_or0 = s_CSAwallace_cska12_nand_11_1 | s_CSAwallace_cska12_csa0_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa4_xor0 = s_CSAwallace_cska12_and_1_3 ^ s_CSAwallace_cska12_and_0_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa4_and0 = s_CSAwallace_cska12_and_1_3 & s_CSAwallace_cska12_and_0_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa5_xor0 = s_CSAwallace_cska12_and_2_3 ^ s_CSAwallace_cska12_and_1_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa5_and0 = s_CSAwallace_cska12_and_2_3 & s_CSAwallace_cska12_and_1_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa5_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa5_xor0 ^ s_CSAwallace_cska12_and_0_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa5_and1 = s_CSAwallace_cska12_csa1_csa_component_fa5_xor0 & s_CSAwallace_cska12_and_0_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa5_or0 = s_CSAwallace_cska12_csa1_csa_component_fa5_and0 | s_CSAwallace_cska12_csa1_csa_component_fa5_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa6_xor0 = s_CSAwallace_cska12_and_3_3 ^ s_CSAwallace_cska12_and_2_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa6_and0 = s_CSAwallace_cska12_and_3_3 & s_CSAwallace_cska12_and_2_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa6_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa6_xor0 ^ s_CSAwallace_cska12_and_1_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa6_and1 = s_CSAwallace_cska12_csa1_csa_component_fa6_xor0 & s_CSAwallace_cska12_and_1_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa6_or0 = s_CSAwallace_cska12_csa1_csa_component_fa6_and0 | s_CSAwallace_cska12_csa1_csa_component_fa6_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa7_xor0 = s_CSAwallace_cska12_and_4_3 ^ s_CSAwallace_cska12_and_3_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa7_and0 = s_CSAwallace_cska12_and_4_3 & s_CSAwallace_cska12_and_3_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa7_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa7_xor0 ^ s_CSAwallace_cska12_and_2_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa7_and1 = s_CSAwallace_cska12_csa1_csa_component_fa7_xor0 & s_CSAwallace_cska12_and_2_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa7_or0 = s_CSAwallace_cska12_csa1_csa_component_fa7_and0 | s_CSAwallace_cska12_csa1_csa_component_fa7_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa8_xor0 = s_CSAwallace_cska12_and_5_3 ^ s_CSAwallace_cska12_and_4_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa8_and0 = s_CSAwallace_cska12_and_5_3 & s_CSAwallace_cska12_and_4_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa8_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa8_xor0 ^ s_CSAwallace_cska12_and_3_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa8_and1 = s_CSAwallace_cska12_csa1_csa_component_fa8_xor0 & s_CSAwallace_cska12_and_3_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa8_or0 = s_CSAwallace_cska12_csa1_csa_component_fa8_and0 | s_CSAwallace_cska12_csa1_csa_component_fa8_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa9_xor0 = s_CSAwallace_cska12_and_6_3 ^ s_CSAwallace_cska12_and_5_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa9_and0 = s_CSAwallace_cska12_and_6_3 & s_CSAwallace_cska12_and_5_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa9_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa9_xor0 ^ s_CSAwallace_cska12_and_4_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa9_and1 = s_CSAwallace_cska12_csa1_csa_component_fa9_xor0 & s_CSAwallace_cska12_and_4_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa9_or0 = s_CSAwallace_cska12_csa1_csa_component_fa9_and0 | s_CSAwallace_cska12_csa1_csa_component_fa9_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa10_xor0 = s_CSAwallace_cska12_and_7_3 ^ s_CSAwallace_cska12_and_6_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa10_and0 = s_CSAwallace_cska12_and_7_3 & s_CSAwallace_cska12_and_6_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa10_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa10_xor0 ^ s_CSAwallace_cska12_and_5_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa10_and1 = s_CSAwallace_cska12_csa1_csa_component_fa10_xor0 & s_CSAwallace_cska12_and_5_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa10_or0 = s_CSAwallace_cska12_csa1_csa_component_fa10_and0 | s_CSAwallace_cska12_csa1_csa_component_fa10_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa11_xor0 = s_CSAwallace_cska12_and_8_3 ^ s_CSAwallace_cska12_and_7_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa11_and0 = s_CSAwallace_cska12_and_8_3 & s_CSAwallace_cska12_and_7_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_and_6_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa11_and1 = s_CSAwallace_cska12_csa1_csa_component_fa11_xor0 & s_CSAwallace_cska12_and_6_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa11_or0 = s_CSAwallace_cska12_csa1_csa_component_fa11_and0 | s_CSAwallace_cska12_csa1_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa12_xor0 = s_CSAwallace_cska12_and_9_3 ^ s_CSAwallace_cska12_and_8_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa12_and0 = s_CSAwallace_cska12_and_9_3 & s_CSAwallace_cska12_and_8_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_and_7_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa12_and1 = s_CSAwallace_cska12_csa1_csa_component_fa12_xor0 & s_CSAwallace_cska12_and_7_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa12_or0 = s_CSAwallace_cska12_csa1_csa_component_fa12_and0 | s_CSAwallace_cska12_csa1_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa13_xor0 = s_CSAwallace_cska12_and_10_3 ^ s_CSAwallace_cska12_and_9_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa13_and0 = s_CSAwallace_cska12_and_10_3 & s_CSAwallace_cska12_and_9_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa13_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa13_xor0 ^ s_CSAwallace_cska12_and_8_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa13_and1 = s_CSAwallace_cska12_csa1_csa_component_fa13_xor0 & s_CSAwallace_cska12_and_8_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa13_or0 = s_CSAwallace_cska12_csa1_csa_component_fa13_and0 | s_CSAwallace_cska12_csa1_csa_component_fa13_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa14_xor0 = s_CSAwallace_cska12_nand_11_3 ^ s_CSAwallace_cska12_and_10_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa14_and0 = s_CSAwallace_cska12_nand_11_3 & s_CSAwallace_cska12_and_10_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa14_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa14_xor0 ^ s_CSAwallace_cska12_and_9_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa14_and1 = s_CSAwallace_cska12_csa1_csa_component_fa14_xor0 & s_CSAwallace_cska12_and_9_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa14_or0 = s_CSAwallace_cska12_csa1_csa_component_fa14_and0 | s_CSAwallace_cska12_csa1_csa_component_fa14_and1;
  assign s_CSAwallace_cska12_csa1_csa_component_fa15_xor0 = ~s_CSAwallace_cska12_nand_11_4;
  assign s_CSAwallace_cska12_csa1_csa_component_fa15_xor1 = s_CSAwallace_cska12_csa1_csa_component_fa15_xor0 ^ s_CSAwallace_cska12_and_10_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa15_and1 = s_CSAwallace_cska12_csa1_csa_component_fa15_xor0 & s_CSAwallace_cska12_and_10_5;
  assign s_CSAwallace_cska12_csa1_csa_component_fa15_or0 = s_CSAwallace_cska12_nand_11_4 | s_CSAwallace_cska12_csa1_csa_component_fa15_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa7_xor0 = s_CSAwallace_cska12_and_1_6 ^ s_CSAwallace_cska12_and_0_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa7_and0 = s_CSAwallace_cska12_and_1_6 & s_CSAwallace_cska12_and_0_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa8_xor0 = s_CSAwallace_cska12_and_2_6 ^ s_CSAwallace_cska12_and_1_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa8_and0 = s_CSAwallace_cska12_and_2_6 & s_CSAwallace_cska12_and_1_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa8_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa8_xor0 ^ s_CSAwallace_cska12_and_0_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa8_and1 = s_CSAwallace_cska12_csa2_csa_component_fa8_xor0 & s_CSAwallace_cska12_and_0_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa8_or0 = s_CSAwallace_cska12_csa2_csa_component_fa8_and0 | s_CSAwallace_cska12_csa2_csa_component_fa8_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa9_xor0 = s_CSAwallace_cska12_and_3_6 ^ s_CSAwallace_cska12_and_2_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa9_and0 = s_CSAwallace_cska12_and_3_6 & s_CSAwallace_cska12_and_2_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa9_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa9_xor0 ^ s_CSAwallace_cska12_and_1_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa9_and1 = s_CSAwallace_cska12_csa2_csa_component_fa9_xor0 & s_CSAwallace_cska12_and_1_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa9_or0 = s_CSAwallace_cska12_csa2_csa_component_fa9_and0 | s_CSAwallace_cska12_csa2_csa_component_fa9_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa10_xor0 = s_CSAwallace_cska12_and_4_6 ^ s_CSAwallace_cska12_and_3_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa10_and0 = s_CSAwallace_cska12_and_4_6 & s_CSAwallace_cska12_and_3_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa10_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa10_xor0 ^ s_CSAwallace_cska12_and_2_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa10_and1 = s_CSAwallace_cska12_csa2_csa_component_fa10_xor0 & s_CSAwallace_cska12_and_2_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa10_or0 = s_CSAwallace_cska12_csa2_csa_component_fa10_and0 | s_CSAwallace_cska12_csa2_csa_component_fa10_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa11_xor0 = s_CSAwallace_cska12_and_5_6 ^ s_CSAwallace_cska12_and_4_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa11_and0 = s_CSAwallace_cska12_and_5_6 & s_CSAwallace_cska12_and_4_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_and_3_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa11_and1 = s_CSAwallace_cska12_csa2_csa_component_fa11_xor0 & s_CSAwallace_cska12_and_3_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa11_or0 = s_CSAwallace_cska12_csa2_csa_component_fa11_and0 | s_CSAwallace_cska12_csa2_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa12_xor0 = s_CSAwallace_cska12_and_6_6 ^ s_CSAwallace_cska12_and_5_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa12_and0 = s_CSAwallace_cska12_and_6_6 & s_CSAwallace_cska12_and_5_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_and_4_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa12_and1 = s_CSAwallace_cska12_csa2_csa_component_fa12_xor0 & s_CSAwallace_cska12_and_4_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa12_or0 = s_CSAwallace_cska12_csa2_csa_component_fa12_and0 | s_CSAwallace_cska12_csa2_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa13_xor0 = s_CSAwallace_cska12_and_7_6 ^ s_CSAwallace_cska12_and_6_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa13_and0 = s_CSAwallace_cska12_and_7_6 & s_CSAwallace_cska12_and_6_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa13_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa13_xor0 ^ s_CSAwallace_cska12_and_5_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa13_and1 = s_CSAwallace_cska12_csa2_csa_component_fa13_xor0 & s_CSAwallace_cska12_and_5_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa13_or0 = s_CSAwallace_cska12_csa2_csa_component_fa13_and0 | s_CSAwallace_cska12_csa2_csa_component_fa13_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa14_xor0 = s_CSAwallace_cska12_and_8_6 ^ s_CSAwallace_cska12_and_7_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa14_and0 = s_CSAwallace_cska12_and_8_6 & s_CSAwallace_cska12_and_7_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa14_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa14_xor0 ^ s_CSAwallace_cska12_and_6_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa14_and1 = s_CSAwallace_cska12_csa2_csa_component_fa14_xor0 & s_CSAwallace_cska12_and_6_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa14_or0 = s_CSAwallace_cska12_csa2_csa_component_fa14_and0 | s_CSAwallace_cska12_csa2_csa_component_fa14_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa15_xor0 = s_CSAwallace_cska12_and_9_6 ^ s_CSAwallace_cska12_and_8_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa15_and0 = s_CSAwallace_cska12_and_9_6 & s_CSAwallace_cska12_and_8_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa15_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa15_xor0 ^ s_CSAwallace_cska12_and_7_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa15_and1 = s_CSAwallace_cska12_csa2_csa_component_fa15_xor0 & s_CSAwallace_cska12_and_7_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa15_or0 = s_CSAwallace_cska12_csa2_csa_component_fa15_and0 | s_CSAwallace_cska12_csa2_csa_component_fa15_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa16_xor0 = s_CSAwallace_cska12_and_10_6 ^ s_CSAwallace_cska12_and_9_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa16_and0 = s_CSAwallace_cska12_and_10_6 & s_CSAwallace_cska12_and_9_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa16_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa16_xor0 ^ s_CSAwallace_cska12_and_8_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa16_and1 = s_CSAwallace_cska12_csa2_csa_component_fa16_xor0 & s_CSAwallace_cska12_and_8_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa16_or0 = s_CSAwallace_cska12_csa2_csa_component_fa16_and0 | s_CSAwallace_cska12_csa2_csa_component_fa16_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa17_xor0 = s_CSAwallace_cska12_nand_11_6 ^ s_CSAwallace_cska12_and_10_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa17_and0 = s_CSAwallace_cska12_nand_11_6 & s_CSAwallace_cska12_and_10_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa17_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa17_xor0 ^ s_CSAwallace_cska12_and_9_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa17_and1 = s_CSAwallace_cska12_csa2_csa_component_fa17_xor0 & s_CSAwallace_cska12_and_9_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa17_or0 = s_CSAwallace_cska12_csa2_csa_component_fa17_and0 | s_CSAwallace_cska12_csa2_csa_component_fa17_and1;
  assign s_CSAwallace_cska12_csa2_csa_component_fa18_xor0 = ~s_CSAwallace_cska12_nand_11_7;
  assign s_CSAwallace_cska12_csa2_csa_component_fa18_xor1 = s_CSAwallace_cska12_csa2_csa_component_fa18_xor0 ^ s_CSAwallace_cska12_and_10_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa18_and1 = s_CSAwallace_cska12_csa2_csa_component_fa18_xor0 & s_CSAwallace_cska12_and_10_8;
  assign s_CSAwallace_cska12_csa2_csa_component_fa18_or0 = s_CSAwallace_cska12_nand_11_7 | s_CSAwallace_cska12_csa2_csa_component_fa18_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa10_xor0 = s_CSAwallace_cska12_and_1_9 ^ s_CSAwallace_cska12_and_0_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa10_and0 = s_CSAwallace_cska12_and_1_9 & s_CSAwallace_cska12_and_0_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa11_xor0 = s_CSAwallace_cska12_and_2_9 ^ s_CSAwallace_cska12_and_1_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa11_and0 = s_CSAwallace_cska12_and_2_9 & s_CSAwallace_cska12_and_1_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_nand_0_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa11_and1 = s_CSAwallace_cska12_csa3_csa_component_fa11_xor0 & s_CSAwallace_cska12_nand_0_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa11_or0 = s_CSAwallace_cska12_csa3_csa_component_fa11_and0 | s_CSAwallace_cska12_csa3_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa12_xor0 = s_CSAwallace_cska12_and_3_9 ^ s_CSAwallace_cska12_and_2_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa12_and0 = s_CSAwallace_cska12_and_3_9 & s_CSAwallace_cska12_and_2_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_nand_1_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa12_and1 = s_CSAwallace_cska12_csa3_csa_component_fa12_xor0 & s_CSAwallace_cska12_nand_1_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa12_or0 = s_CSAwallace_cska12_csa3_csa_component_fa12_and0 | s_CSAwallace_cska12_csa3_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa13_xor0 = s_CSAwallace_cska12_and_4_9 ^ s_CSAwallace_cska12_and_3_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa13_and0 = s_CSAwallace_cska12_and_4_9 & s_CSAwallace_cska12_and_3_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa13_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa13_xor0 ^ s_CSAwallace_cska12_nand_2_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa13_and1 = s_CSAwallace_cska12_csa3_csa_component_fa13_xor0 & s_CSAwallace_cska12_nand_2_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa13_or0 = s_CSAwallace_cska12_csa3_csa_component_fa13_and0 | s_CSAwallace_cska12_csa3_csa_component_fa13_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa14_xor0 = s_CSAwallace_cska12_and_5_9 ^ s_CSAwallace_cska12_and_4_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa14_and0 = s_CSAwallace_cska12_and_5_9 & s_CSAwallace_cska12_and_4_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa14_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa14_xor0 ^ s_CSAwallace_cska12_nand_3_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa14_and1 = s_CSAwallace_cska12_csa3_csa_component_fa14_xor0 & s_CSAwallace_cska12_nand_3_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa14_or0 = s_CSAwallace_cska12_csa3_csa_component_fa14_and0 | s_CSAwallace_cska12_csa3_csa_component_fa14_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa15_xor0 = s_CSAwallace_cska12_and_6_9 ^ s_CSAwallace_cska12_and_5_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa15_and0 = s_CSAwallace_cska12_and_6_9 & s_CSAwallace_cska12_and_5_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa15_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa15_xor0 ^ s_CSAwallace_cska12_nand_4_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa15_and1 = s_CSAwallace_cska12_csa3_csa_component_fa15_xor0 & s_CSAwallace_cska12_nand_4_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa15_or0 = s_CSAwallace_cska12_csa3_csa_component_fa15_and0 | s_CSAwallace_cska12_csa3_csa_component_fa15_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa16_xor0 = s_CSAwallace_cska12_and_7_9 ^ s_CSAwallace_cska12_and_6_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa16_and0 = s_CSAwallace_cska12_and_7_9 & s_CSAwallace_cska12_and_6_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa16_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa16_xor0 ^ s_CSAwallace_cska12_nand_5_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa16_and1 = s_CSAwallace_cska12_csa3_csa_component_fa16_xor0 & s_CSAwallace_cska12_nand_5_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa16_or0 = s_CSAwallace_cska12_csa3_csa_component_fa16_and0 | s_CSAwallace_cska12_csa3_csa_component_fa16_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa17_xor0 = s_CSAwallace_cska12_and_8_9 ^ s_CSAwallace_cska12_and_7_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa17_and0 = s_CSAwallace_cska12_and_8_9 & s_CSAwallace_cska12_and_7_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa17_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa17_xor0 ^ s_CSAwallace_cska12_nand_6_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa17_and1 = s_CSAwallace_cska12_csa3_csa_component_fa17_xor0 & s_CSAwallace_cska12_nand_6_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa17_or0 = s_CSAwallace_cska12_csa3_csa_component_fa17_and0 | s_CSAwallace_cska12_csa3_csa_component_fa17_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa18_xor0 = s_CSAwallace_cska12_and_9_9 ^ s_CSAwallace_cska12_and_8_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa18_and0 = s_CSAwallace_cska12_and_9_9 & s_CSAwallace_cska12_and_8_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa18_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa18_xor0 ^ s_CSAwallace_cska12_nand_7_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa18_and1 = s_CSAwallace_cska12_csa3_csa_component_fa18_xor0 & s_CSAwallace_cska12_nand_7_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa18_or0 = s_CSAwallace_cska12_csa3_csa_component_fa18_and0 | s_CSAwallace_cska12_csa3_csa_component_fa18_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa19_xor0 = s_CSAwallace_cska12_and_10_9 ^ s_CSAwallace_cska12_and_9_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa19_and0 = s_CSAwallace_cska12_and_10_9 & s_CSAwallace_cska12_and_9_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa19_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa19_xor0 ^ s_CSAwallace_cska12_nand_8_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa19_and1 = s_CSAwallace_cska12_csa3_csa_component_fa19_xor0 & s_CSAwallace_cska12_nand_8_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa19_or0 = s_CSAwallace_cska12_csa3_csa_component_fa19_and0 | s_CSAwallace_cska12_csa3_csa_component_fa19_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa20_xor0 = s_CSAwallace_cska12_nand_11_9 ^ s_CSAwallace_cska12_and_10_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa20_and0 = s_CSAwallace_cska12_nand_11_9 & s_CSAwallace_cska12_and_10_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa20_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa20_xor0 ^ s_CSAwallace_cska12_nand_9_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa20_and1 = s_CSAwallace_cska12_csa3_csa_component_fa20_xor0 & s_CSAwallace_cska12_nand_9_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa20_or0 = s_CSAwallace_cska12_csa3_csa_component_fa20_and0 | s_CSAwallace_cska12_csa3_csa_component_fa20_and1;
  assign s_CSAwallace_cska12_csa3_csa_component_fa21_xor0 = ~s_CSAwallace_cska12_nand_11_10;
  assign s_CSAwallace_cska12_csa3_csa_component_fa21_xor1 = s_CSAwallace_cska12_csa3_csa_component_fa21_xor0 ^ s_CSAwallace_cska12_nand_10_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa21_and1 = s_CSAwallace_cska12_csa3_csa_component_fa21_xor0 & s_CSAwallace_cska12_nand_10_11;
  assign s_CSAwallace_cska12_csa3_csa_component_fa21_or0 = s_CSAwallace_cska12_nand_11_10 | s_CSAwallace_cska12_csa3_csa_component_fa21_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa2_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa2_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa1_and0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa2_and0 = s_CSAwallace_cska12_csa0_csa_component_fa2_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa1_and0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa3_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa3_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa2_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa3_and0 = s_CSAwallace_cska12_csa0_csa_component_fa3_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa2_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa3_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa3_xor0 ^ s_CSAwallace_cska12_and_0_3;
  assign s_CSAwallace_cska12_csa4_csa_component_fa3_and1 = s_CSAwallace_cska12_csa4_csa_component_fa3_xor0 & s_CSAwallace_cska12_and_0_3;
  assign s_CSAwallace_cska12_csa4_csa_component_fa3_or0 = s_CSAwallace_cska12_csa4_csa_component_fa3_and0 | s_CSAwallace_cska12_csa4_csa_component_fa3_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa4_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa4_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa3_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa4_and0 = s_CSAwallace_cska12_csa0_csa_component_fa4_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa3_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa4_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa4_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa4_xor0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa4_and1 = s_CSAwallace_cska12_csa4_csa_component_fa4_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa4_xor0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa4_or0 = s_CSAwallace_cska12_csa4_csa_component_fa4_and0 | s_CSAwallace_cska12_csa4_csa_component_fa4_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa5_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa5_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa4_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa5_and0 = s_CSAwallace_cska12_csa0_csa_component_fa5_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa4_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa5_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa5_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa5_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa5_and1 = s_CSAwallace_cska12_csa4_csa_component_fa5_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa5_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa5_or0 = s_CSAwallace_cska12_csa4_csa_component_fa5_and0 | s_CSAwallace_cska12_csa4_csa_component_fa5_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa6_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa6_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa5_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa6_and0 = s_CSAwallace_cska12_csa0_csa_component_fa6_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa5_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa6_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa6_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa6_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa6_and1 = s_CSAwallace_cska12_csa4_csa_component_fa6_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa6_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa6_or0 = s_CSAwallace_cska12_csa4_csa_component_fa6_and0 | s_CSAwallace_cska12_csa4_csa_component_fa6_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa7_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa7_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa6_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa7_and0 = s_CSAwallace_cska12_csa0_csa_component_fa7_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa6_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa7_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa7_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa7_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa7_and1 = s_CSAwallace_cska12_csa4_csa_component_fa7_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa7_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa7_or0 = s_CSAwallace_cska12_csa4_csa_component_fa7_and0 | s_CSAwallace_cska12_csa4_csa_component_fa7_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa8_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa8_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa7_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa8_and0 = s_CSAwallace_cska12_csa0_csa_component_fa8_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa7_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa8_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa8_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa8_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa8_and1 = s_CSAwallace_cska12_csa4_csa_component_fa8_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa8_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa8_or0 = s_CSAwallace_cska12_csa4_csa_component_fa8_and0 | s_CSAwallace_cska12_csa4_csa_component_fa8_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa9_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa9_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa9_and0 = s_CSAwallace_cska12_csa0_csa_component_fa9_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa9_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa9_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa9_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa9_and1 = s_CSAwallace_cska12_csa4_csa_component_fa9_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa9_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa9_or0 = s_CSAwallace_cska12_csa4_csa_component_fa9_and0 | s_CSAwallace_cska12_csa4_csa_component_fa9_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa10_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa10_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa10_and0 = s_CSAwallace_cska12_csa0_csa_component_fa10_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa10_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa10_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa10_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa10_and1 = s_CSAwallace_cska12_csa4_csa_component_fa10_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa10_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa10_or0 = s_CSAwallace_cska12_csa4_csa_component_fa10_and0 | s_CSAwallace_cska12_csa4_csa_component_fa10_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa11_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa11_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa11_and0 = s_CSAwallace_cska12_csa0_csa_component_fa11_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa11_and1 = s_CSAwallace_cska12_csa4_csa_component_fa11_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa11_or0 = s_CSAwallace_cska12_csa4_csa_component_fa11_and0 | s_CSAwallace_cska12_csa4_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa12_xor0 = s_CSAwallace_cska12_csa0_csa_component_fa12_xor1 ^ s_CSAwallace_cska12_csa0_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa12_and0 = s_CSAwallace_cska12_csa0_csa_component_fa12_xor1 & s_CSAwallace_cska12_csa0_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa12_and1 = s_CSAwallace_cska12_csa4_csa_component_fa12_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa12_or0 = s_CSAwallace_cska12_csa4_csa_component_fa12_and0 | s_CSAwallace_cska12_csa4_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa13_xor0 = s_CSAwallace_cska12_nand_11_2 ^ s_CSAwallace_cska12_csa0_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa13_and0 = s_CSAwallace_cska12_nand_11_2 & s_CSAwallace_cska12_csa0_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa4_csa_component_fa13_xor1 = s_CSAwallace_cska12_csa4_csa_component_fa13_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa13_and1 = s_CSAwallace_cska12_csa4_csa_component_fa13_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa4_csa_component_fa13_or0 = s_CSAwallace_cska12_csa4_csa_component_fa13_and0 | s_CSAwallace_cska12_csa4_csa_component_fa13_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa6_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa5_or0 ^ s_CSAwallace_cska12_and_0_6;
  assign s_CSAwallace_cska12_csa5_csa_component_fa6_and0 = s_CSAwallace_cska12_csa1_csa_component_fa5_or0 & s_CSAwallace_cska12_and_0_6;
  assign s_CSAwallace_cska12_csa5_csa_component_fa7_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa6_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa7_xor0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa7_and0 = s_CSAwallace_cska12_csa1_csa_component_fa6_or0 & s_CSAwallace_cska12_csa2_csa_component_fa7_xor0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa8_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa7_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa8_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa8_and0 = s_CSAwallace_cska12_csa1_csa_component_fa7_or0 & s_CSAwallace_cska12_csa2_csa_component_fa8_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa8_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa8_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa7_and0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa8_and1 = s_CSAwallace_cska12_csa5_csa_component_fa8_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa7_and0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa8_or0 = s_CSAwallace_cska12_csa5_csa_component_fa8_and0 | s_CSAwallace_cska12_csa5_csa_component_fa8_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa9_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa8_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa9_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa9_and0 = s_CSAwallace_cska12_csa1_csa_component_fa8_or0 & s_CSAwallace_cska12_csa2_csa_component_fa9_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa9_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa9_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa9_and1 = s_CSAwallace_cska12_csa5_csa_component_fa9_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa9_or0 = s_CSAwallace_cska12_csa5_csa_component_fa9_and0 | s_CSAwallace_cska12_csa5_csa_component_fa9_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa10_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa9_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa10_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa10_and0 = s_CSAwallace_cska12_csa1_csa_component_fa9_or0 & s_CSAwallace_cska12_csa2_csa_component_fa10_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa10_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa10_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa10_and1 = s_CSAwallace_cska12_csa5_csa_component_fa10_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa10_or0 = s_CSAwallace_cska12_csa5_csa_component_fa10_and0 | s_CSAwallace_cska12_csa5_csa_component_fa10_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa11_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa10_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa11_and0 = s_CSAwallace_cska12_csa1_csa_component_fa10_or0 & s_CSAwallace_cska12_csa2_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa11_and1 = s_CSAwallace_cska12_csa5_csa_component_fa11_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa11_or0 = s_CSAwallace_cska12_csa5_csa_component_fa11_and0 | s_CSAwallace_cska12_csa5_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa12_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa11_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa12_and0 = s_CSAwallace_cska12_csa1_csa_component_fa11_or0 & s_CSAwallace_cska12_csa2_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa12_and1 = s_CSAwallace_cska12_csa5_csa_component_fa12_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa12_or0 = s_CSAwallace_cska12_csa5_csa_component_fa12_and0 | s_CSAwallace_cska12_csa5_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa13_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa12_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa13_and0 = s_CSAwallace_cska12_csa1_csa_component_fa12_or0 & s_CSAwallace_cska12_csa2_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa13_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa13_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa13_and1 = s_CSAwallace_cska12_csa5_csa_component_fa13_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa13_or0 = s_CSAwallace_cska12_csa5_csa_component_fa13_and0 | s_CSAwallace_cska12_csa5_csa_component_fa13_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa14_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa13_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa14_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa14_and0 = s_CSAwallace_cska12_csa1_csa_component_fa13_or0 & s_CSAwallace_cska12_csa2_csa_component_fa14_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa14_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa14_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa14_and1 = s_CSAwallace_cska12_csa5_csa_component_fa14_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa14_or0 = s_CSAwallace_cska12_csa5_csa_component_fa14_and0 | s_CSAwallace_cska12_csa5_csa_component_fa14_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa15_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa14_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa15_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa15_and0 = s_CSAwallace_cska12_csa1_csa_component_fa14_or0 & s_CSAwallace_cska12_csa2_csa_component_fa15_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa15_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa15_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa15_and1 = s_CSAwallace_cska12_csa5_csa_component_fa15_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa15_or0 = s_CSAwallace_cska12_csa5_csa_component_fa15_and0 | s_CSAwallace_cska12_csa5_csa_component_fa15_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa16_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa15_or0 ^ s_CSAwallace_cska12_csa2_csa_component_fa16_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa16_and0 = s_CSAwallace_cska12_csa1_csa_component_fa15_or0 & s_CSAwallace_cska12_csa2_csa_component_fa16_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa16_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa16_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa16_and1 = s_CSAwallace_cska12_csa5_csa_component_fa16_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa16_or0 = s_CSAwallace_cska12_csa5_csa_component_fa16_and0 | s_CSAwallace_cska12_csa5_csa_component_fa16_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa17_xor0 = ~s_CSAwallace_cska12_csa2_csa_component_fa17_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa17_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa17_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa17_and1 = s_CSAwallace_cska12_csa5_csa_component_fa17_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa17_or0 = s_CSAwallace_cska12_csa2_csa_component_fa17_xor1 | s_CSAwallace_cska12_csa5_csa_component_fa17_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa18_xor0 = ~s_CSAwallace_cska12_csa2_csa_component_fa18_xor1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa18_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa18_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa18_and1 = s_CSAwallace_cska12_csa5_csa_component_fa18_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa18_or0 = s_CSAwallace_cska12_csa2_csa_component_fa18_xor1 | s_CSAwallace_cska12_csa5_csa_component_fa18_and1;
  assign s_CSAwallace_cska12_csa5_csa_component_fa19_xor0 = ~s_CSAwallace_cska12_nand_11_8;
  assign s_CSAwallace_cska12_csa5_csa_component_fa19_xor1 = s_CSAwallace_cska12_csa5_csa_component_fa19_xor0 ^ s_CSAwallace_cska12_csa2_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa19_and1 = s_CSAwallace_cska12_csa5_csa_component_fa19_xor0 & s_CSAwallace_cska12_csa2_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_csa5_csa_component_fa19_or0 = s_CSAwallace_cska12_nand_11_8 | s_CSAwallace_cska12_csa5_csa_component_fa19_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa3_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa3_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa2_and0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa3_and0 = s_CSAwallace_cska12_csa4_csa_component_fa3_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa2_and0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa4_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa4_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa3_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa4_and0 = s_CSAwallace_cska12_csa4_csa_component_fa4_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa3_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa5_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa5_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa4_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa5_and0 = s_CSAwallace_cska12_csa4_csa_component_fa5_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa4_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa5_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa5_xor0 ^ s_CSAwallace_cska12_csa1_csa_component_fa4_and0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa5_and1 = s_CSAwallace_cska12_csa6_csa_component_fa5_xor0 & s_CSAwallace_cska12_csa1_csa_component_fa4_and0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa5_or0 = s_CSAwallace_cska12_csa6_csa_component_fa5_and0 | s_CSAwallace_cska12_csa6_csa_component_fa5_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa6_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa6_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa5_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa6_and0 = s_CSAwallace_cska12_csa4_csa_component_fa6_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa5_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa6_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa6_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa6_xor0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa6_and1 = s_CSAwallace_cska12_csa6_csa_component_fa6_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa6_xor0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa6_or0 = s_CSAwallace_cska12_csa6_csa_component_fa6_and0 | s_CSAwallace_cska12_csa6_csa_component_fa6_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa7_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa7_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa6_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa7_and0 = s_CSAwallace_cska12_csa4_csa_component_fa7_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa6_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa7_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa7_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa7_xor0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa7_and1 = s_CSAwallace_cska12_csa6_csa_component_fa7_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa7_xor0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa7_or0 = s_CSAwallace_cska12_csa6_csa_component_fa7_and0 | s_CSAwallace_cska12_csa6_csa_component_fa7_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa8_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa8_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa7_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa8_and0 = s_CSAwallace_cska12_csa4_csa_component_fa8_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa7_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa8_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa8_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa8_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa8_and1 = s_CSAwallace_cska12_csa6_csa_component_fa8_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa8_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa8_or0 = s_CSAwallace_cska12_csa6_csa_component_fa8_and0 | s_CSAwallace_cska12_csa6_csa_component_fa8_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa9_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa9_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa9_and0 = s_CSAwallace_cska12_csa4_csa_component_fa9_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa9_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa9_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa9_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa9_and1 = s_CSAwallace_cska12_csa6_csa_component_fa9_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa9_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa9_or0 = s_CSAwallace_cska12_csa6_csa_component_fa9_and0 | s_CSAwallace_cska12_csa6_csa_component_fa9_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa10_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa10_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa10_and0 = s_CSAwallace_cska12_csa4_csa_component_fa10_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa10_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa10_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa10_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa10_and1 = s_CSAwallace_cska12_csa6_csa_component_fa10_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa10_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa10_or0 = s_CSAwallace_cska12_csa6_csa_component_fa10_and0 | s_CSAwallace_cska12_csa6_csa_component_fa10_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa11_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa11_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa11_and0 = s_CSAwallace_cska12_csa4_csa_component_fa11_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa11_and1 = s_CSAwallace_cska12_csa6_csa_component_fa11_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa11_or0 = s_CSAwallace_cska12_csa6_csa_component_fa11_and0 | s_CSAwallace_cska12_csa6_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa12_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa12_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa12_and0 = s_CSAwallace_cska12_csa4_csa_component_fa12_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa12_and1 = s_CSAwallace_cska12_csa6_csa_component_fa12_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa12_or0 = s_CSAwallace_cska12_csa6_csa_component_fa12_and0 | s_CSAwallace_cska12_csa6_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa13_xor0 = s_CSAwallace_cska12_csa4_csa_component_fa13_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa13_and0 = s_CSAwallace_cska12_csa4_csa_component_fa13_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa13_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa13_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa13_and1 = s_CSAwallace_cska12_csa6_csa_component_fa13_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa13_or0 = s_CSAwallace_cska12_csa6_csa_component_fa13_and0 | s_CSAwallace_cska12_csa6_csa_component_fa13_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa14_xor0 = s_CSAwallace_cska12_csa1_csa_component_fa14_xor1 ^ s_CSAwallace_cska12_csa4_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa14_and0 = s_CSAwallace_cska12_csa1_csa_component_fa14_xor1 & s_CSAwallace_cska12_csa4_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa6_csa_component_fa14_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa14_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa14_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa14_and1 = s_CSAwallace_cska12_csa6_csa_component_fa14_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa14_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa14_or0 = s_CSAwallace_cska12_csa6_csa_component_fa14_and0 | s_CSAwallace_cska12_csa6_csa_component_fa14_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa15_xor0 = ~s_CSAwallace_cska12_csa1_csa_component_fa15_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa15_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa15_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa15_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa15_and1 = s_CSAwallace_cska12_csa6_csa_component_fa15_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa15_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa15_or0 = s_CSAwallace_cska12_csa1_csa_component_fa15_xor1 | s_CSAwallace_cska12_csa6_csa_component_fa15_and1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa16_xor0 = ~s_CSAwallace_cska12_nand_11_5;
  assign s_CSAwallace_cska12_csa6_csa_component_fa16_xor1 = s_CSAwallace_cska12_csa6_csa_component_fa16_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa16_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa16_and1 = s_CSAwallace_cska12_csa6_csa_component_fa16_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa16_xor1;
  assign s_CSAwallace_cska12_csa6_csa_component_fa16_or0 = s_CSAwallace_cska12_nand_11_5 | s_CSAwallace_cska12_csa6_csa_component_fa16_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa9_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa8_or0 ^ s_CSAwallace_cska12_and_0_9;
  assign s_CSAwallace_cska12_csa7_csa_component_fa9_and0 = s_CSAwallace_cska12_csa5_csa_component_fa8_or0 & s_CSAwallace_cska12_and_0_9;
  assign s_CSAwallace_cska12_csa7_csa_component_fa10_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa9_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa10_xor0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa10_and0 = s_CSAwallace_cska12_csa5_csa_component_fa9_or0 & s_CSAwallace_cska12_csa3_csa_component_fa10_xor0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa11_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa10_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa11_and0 = s_CSAwallace_cska12_csa5_csa_component_fa10_or0 & s_CSAwallace_cska12_csa3_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa10_and0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa11_and1 = s_CSAwallace_cska12_csa7_csa_component_fa11_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa10_and0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa11_or0 = s_CSAwallace_cska12_csa7_csa_component_fa11_and0 | s_CSAwallace_cska12_csa7_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa12_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa11_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa12_and0 = s_CSAwallace_cska12_csa5_csa_component_fa11_or0 & s_CSAwallace_cska12_csa3_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa12_and1 = s_CSAwallace_cska12_csa7_csa_component_fa12_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa12_or0 = s_CSAwallace_cska12_csa7_csa_component_fa12_and0 | s_CSAwallace_cska12_csa7_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa13_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa12_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa13_and0 = s_CSAwallace_cska12_csa5_csa_component_fa12_or0 & s_CSAwallace_cska12_csa3_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa13_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa13_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa13_and1 = s_CSAwallace_cska12_csa7_csa_component_fa13_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa13_or0 = s_CSAwallace_cska12_csa7_csa_component_fa13_and0 | s_CSAwallace_cska12_csa7_csa_component_fa13_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa14_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa13_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa14_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa14_and0 = s_CSAwallace_cska12_csa5_csa_component_fa13_or0 & s_CSAwallace_cska12_csa3_csa_component_fa14_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa14_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa14_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa14_and1 = s_CSAwallace_cska12_csa7_csa_component_fa14_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa14_or0 = s_CSAwallace_cska12_csa7_csa_component_fa14_and0 | s_CSAwallace_cska12_csa7_csa_component_fa14_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa15_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa14_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa15_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa15_and0 = s_CSAwallace_cska12_csa5_csa_component_fa14_or0 & s_CSAwallace_cska12_csa3_csa_component_fa15_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa15_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa15_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa15_and1 = s_CSAwallace_cska12_csa7_csa_component_fa15_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa15_or0 = s_CSAwallace_cska12_csa7_csa_component_fa15_and0 | s_CSAwallace_cska12_csa7_csa_component_fa15_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa16_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa15_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa16_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa16_and0 = s_CSAwallace_cska12_csa5_csa_component_fa15_or0 & s_CSAwallace_cska12_csa3_csa_component_fa16_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa16_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa16_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa16_and1 = s_CSAwallace_cska12_csa7_csa_component_fa16_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa16_or0 = s_CSAwallace_cska12_csa7_csa_component_fa16_and0 | s_CSAwallace_cska12_csa7_csa_component_fa16_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa17_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa16_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa17_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa17_and0 = s_CSAwallace_cska12_csa5_csa_component_fa16_or0 & s_CSAwallace_cska12_csa3_csa_component_fa17_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa17_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa17_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa17_and1 = s_CSAwallace_cska12_csa7_csa_component_fa17_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa17_or0 = s_CSAwallace_cska12_csa7_csa_component_fa17_and0 | s_CSAwallace_cska12_csa7_csa_component_fa17_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa18_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa17_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa18_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa18_and0 = s_CSAwallace_cska12_csa5_csa_component_fa17_or0 & s_CSAwallace_cska12_csa3_csa_component_fa18_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa18_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa18_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa18_and1 = s_CSAwallace_cska12_csa7_csa_component_fa18_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa18_or0 = s_CSAwallace_cska12_csa7_csa_component_fa18_and0 | s_CSAwallace_cska12_csa7_csa_component_fa18_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa19_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa18_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa19_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa19_and0 = s_CSAwallace_cska12_csa5_csa_component_fa18_or0 & s_CSAwallace_cska12_csa3_csa_component_fa19_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa19_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa19_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa19_and1 = s_CSAwallace_cska12_csa7_csa_component_fa19_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa19_or0 = s_CSAwallace_cska12_csa7_csa_component_fa19_and0 | s_CSAwallace_cska12_csa7_csa_component_fa19_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa20_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa19_or0 ^ s_CSAwallace_cska12_csa3_csa_component_fa20_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa20_and0 = s_CSAwallace_cska12_csa5_csa_component_fa19_or0 & s_CSAwallace_cska12_csa3_csa_component_fa20_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa20_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa20_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa19_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa20_and1 = s_CSAwallace_cska12_csa7_csa_component_fa20_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa19_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa20_or0 = s_CSAwallace_cska12_csa7_csa_component_fa20_and0 | s_CSAwallace_cska12_csa7_csa_component_fa20_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa21_xor0 = ~s_CSAwallace_cska12_csa3_csa_component_fa21_xor1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa21_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa21_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa20_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa21_and1 = s_CSAwallace_cska12_csa7_csa_component_fa21_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa20_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa21_or0 = s_CSAwallace_cska12_csa3_csa_component_fa21_xor1 | s_CSAwallace_cska12_csa7_csa_component_fa21_and1;
  assign s_CSAwallace_cska12_csa7_csa_component_fa22_xor0 = ~s_CSAwallace_cska12_and_11_11;
  assign s_CSAwallace_cska12_csa7_csa_component_fa22_xor1 = s_CSAwallace_cska12_csa7_csa_component_fa22_xor0 ^ s_CSAwallace_cska12_csa3_csa_component_fa21_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa22_and1 = s_CSAwallace_cska12_csa7_csa_component_fa22_xor0 & s_CSAwallace_cska12_csa3_csa_component_fa21_or0;
  assign s_CSAwallace_cska12_csa7_csa_component_fa22_or0 = s_CSAwallace_cska12_and_11_11 | s_CSAwallace_cska12_csa7_csa_component_fa22_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa4_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa4_xor0 ^ s_CSAwallace_cska12_csa6_csa_component_fa3_and0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa4_and0 = s_CSAwallace_cska12_csa6_csa_component_fa4_xor0 & s_CSAwallace_cska12_csa6_csa_component_fa3_and0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa5_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa5_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa4_and0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa5_and0 = s_CSAwallace_cska12_csa6_csa_component_fa5_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa4_and0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa6_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa6_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa5_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa6_and0 = s_CSAwallace_cska12_csa6_csa_component_fa6_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa5_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa7_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa7_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa6_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa7_and0 = s_CSAwallace_cska12_csa6_csa_component_fa7_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa6_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa7_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa7_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa6_and0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa7_and1 = s_CSAwallace_cska12_csa8_csa_component_fa7_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa6_and0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa7_or0 = s_CSAwallace_cska12_csa8_csa_component_fa7_and0 | s_CSAwallace_cska12_csa8_csa_component_fa7_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa8_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa8_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa7_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa8_and0 = s_CSAwallace_cska12_csa6_csa_component_fa8_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa7_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa8_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa8_xor0 ^ s_CSAwallace_cska12_csa5_csa_component_fa7_and0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa8_and1 = s_CSAwallace_cska12_csa8_csa_component_fa8_xor0 & s_CSAwallace_cska12_csa5_csa_component_fa7_and0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa8_or0 = s_CSAwallace_cska12_csa8_csa_component_fa8_and0 | s_CSAwallace_cska12_csa8_csa_component_fa8_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa9_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa9_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa9_and0 = s_CSAwallace_cska12_csa6_csa_component_fa9_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa9_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa9_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa9_xor0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa9_and1 = s_CSAwallace_cska12_csa8_csa_component_fa9_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa9_xor0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa9_or0 = s_CSAwallace_cska12_csa8_csa_component_fa9_and0 | s_CSAwallace_cska12_csa8_csa_component_fa9_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa10_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa10_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa10_and0 = s_CSAwallace_cska12_csa6_csa_component_fa10_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa10_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa10_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa10_xor0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa10_and1 = s_CSAwallace_cska12_csa8_csa_component_fa10_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa10_xor0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa10_or0 = s_CSAwallace_cska12_csa8_csa_component_fa10_and0 | s_CSAwallace_cska12_csa8_csa_component_fa10_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa11_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa11_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa11_and0 = s_CSAwallace_cska12_csa6_csa_component_fa11_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa11_and1 = s_CSAwallace_cska12_csa8_csa_component_fa11_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa11_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa11_or0 = s_CSAwallace_cska12_csa8_csa_component_fa11_and0 | s_CSAwallace_cska12_csa8_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa12_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa12_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa12_and0 = s_CSAwallace_cska12_csa6_csa_component_fa12_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa12_and1 = s_CSAwallace_cska12_csa8_csa_component_fa12_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa12_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa12_or0 = s_CSAwallace_cska12_csa8_csa_component_fa12_and0 | s_CSAwallace_cska12_csa8_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa13_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa13_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa13_and0 = s_CSAwallace_cska12_csa6_csa_component_fa13_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa13_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa13_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa13_and1 = s_CSAwallace_cska12_csa8_csa_component_fa13_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa13_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa13_or0 = s_CSAwallace_cska12_csa8_csa_component_fa13_and0 | s_CSAwallace_cska12_csa8_csa_component_fa13_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa14_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa14_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa14_and0 = s_CSAwallace_cska12_csa6_csa_component_fa14_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa14_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa14_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa14_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa14_and1 = s_CSAwallace_cska12_csa8_csa_component_fa14_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa14_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa14_or0 = s_CSAwallace_cska12_csa8_csa_component_fa14_and0 | s_CSAwallace_cska12_csa8_csa_component_fa14_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa15_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa15_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa15_and0 = s_CSAwallace_cska12_csa6_csa_component_fa15_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa15_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa15_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa15_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa15_and1 = s_CSAwallace_cska12_csa8_csa_component_fa15_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa15_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa15_or0 = s_CSAwallace_cska12_csa8_csa_component_fa15_and0 | s_CSAwallace_cska12_csa8_csa_component_fa15_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa16_xor0 = s_CSAwallace_cska12_csa6_csa_component_fa16_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa16_and0 = s_CSAwallace_cska12_csa6_csa_component_fa16_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa16_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa16_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa16_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa16_and1 = s_CSAwallace_cska12_csa8_csa_component_fa16_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa16_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa16_or0 = s_CSAwallace_cska12_csa8_csa_component_fa16_and0 | s_CSAwallace_cska12_csa8_csa_component_fa16_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa17_xor0 = s_CSAwallace_cska12_csa5_csa_component_fa17_xor1 ^ s_CSAwallace_cska12_csa6_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa17_and0 = s_CSAwallace_cska12_csa5_csa_component_fa17_xor1 & s_CSAwallace_cska12_csa6_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa8_csa_component_fa17_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa17_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa17_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa17_and1 = s_CSAwallace_cska12_csa8_csa_component_fa17_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa17_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa17_or0 = s_CSAwallace_cska12_csa8_csa_component_fa17_and0 | s_CSAwallace_cska12_csa8_csa_component_fa17_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa18_xor0 = ~s_CSAwallace_cska12_csa5_csa_component_fa18_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa18_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa18_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa18_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa18_and1 = s_CSAwallace_cska12_csa8_csa_component_fa18_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa18_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa18_or0 = s_CSAwallace_cska12_csa5_csa_component_fa18_xor1 | s_CSAwallace_cska12_csa8_csa_component_fa18_and1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa19_xor0 = ~s_CSAwallace_cska12_csa5_csa_component_fa19_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa19_xor1 = s_CSAwallace_cska12_csa8_csa_component_fa19_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa19_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa19_and1 = s_CSAwallace_cska12_csa8_csa_component_fa19_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa19_xor1;
  assign s_CSAwallace_cska12_csa8_csa_component_fa19_or0 = s_CSAwallace_cska12_csa5_csa_component_fa19_xor1 | s_CSAwallace_cska12_csa8_csa_component_fa19_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa5_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa5_xor0 ^ s_CSAwallace_cska12_csa8_csa_component_fa4_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa5_and0 = s_CSAwallace_cska12_csa8_csa_component_fa5_xor0 & s_CSAwallace_cska12_csa8_csa_component_fa4_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa6_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa6_xor0 ^ s_CSAwallace_cska12_csa8_csa_component_fa5_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa6_and0 = s_CSAwallace_cska12_csa8_csa_component_fa6_xor0 & s_CSAwallace_cska12_csa8_csa_component_fa5_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa7_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa7_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa6_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa7_and0 = s_CSAwallace_cska12_csa8_csa_component_fa7_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa6_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa8_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa8_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa7_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa8_and0 = s_CSAwallace_cska12_csa8_csa_component_fa8_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa7_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa9_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa9_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa9_and0 = s_CSAwallace_cska12_csa8_csa_component_fa9_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa8_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa10_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa10_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa10_and0 = s_CSAwallace_cska12_csa8_csa_component_fa10_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa9_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa10_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa10_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa9_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa10_and1 = s_CSAwallace_cska12_csa9_csa_component_fa10_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa9_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa10_or0 = s_CSAwallace_cska12_csa9_csa_component_fa10_and0 | s_CSAwallace_cska12_csa9_csa_component_fa10_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa11_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa11_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa11_and0 = s_CSAwallace_cska12_csa8_csa_component_fa11_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa11_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa11_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa10_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa11_and1 = s_CSAwallace_cska12_csa9_csa_component_fa11_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa10_and0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa11_or0 = s_CSAwallace_cska12_csa9_csa_component_fa11_and0 | s_CSAwallace_cska12_csa9_csa_component_fa11_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa12_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa12_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa12_and0 = s_CSAwallace_cska12_csa8_csa_component_fa12_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa12_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa12_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa12_and1 = s_CSAwallace_cska12_csa9_csa_component_fa12_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa12_or0 = s_CSAwallace_cska12_csa9_csa_component_fa12_and0 | s_CSAwallace_cska12_csa9_csa_component_fa12_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa13_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa13_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa13_and0 = s_CSAwallace_cska12_csa8_csa_component_fa13_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa13_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa13_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa13_and1 = s_CSAwallace_cska12_csa9_csa_component_fa13_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa13_or0 = s_CSAwallace_cska12_csa9_csa_component_fa13_and0 | s_CSAwallace_cska12_csa9_csa_component_fa13_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa14_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa14_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa14_and0 = s_CSAwallace_cska12_csa8_csa_component_fa14_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa14_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa14_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa14_and1 = s_CSAwallace_cska12_csa9_csa_component_fa14_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa14_or0 = s_CSAwallace_cska12_csa9_csa_component_fa14_and0 | s_CSAwallace_cska12_csa9_csa_component_fa14_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa15_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa15_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa15_and0 = s_CSAwallace_cska12_csa8_csa_component_fa15_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa15_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa15_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa15_and1 = s_CSAwallace_cska12_csa9_csa_component_fa15_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa15_or0 = s_CSAwallace_cska12_csa9_csa_component_fa15_and0 | s_CSAwallace_cska12_csa9_csa_component_fa15_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa16_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa16_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa16_and0 = s_CSAwallace_cska12_csa8_csa_component_fa16_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa16_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa16_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa16_and1 = s_CSAwallace_cska12_csa9_csa_component_fa16_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa16_or0 = s_CSAwallace_cska12_csa9_csa_component_fa16_and0 | s_CSAwallace_cska12_csa9_csa_component_fa16_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa17_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa17_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa17_and0 = s_CSAwallace_cska12_csa8_csa_component_fa17_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa17_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa17_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa17_and1 = s_CSAwallace_cska12_csa9_csa_component_fa17_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa17_or0 = s_CSAwallace_cska12_csa9_csa_component_fa17_and0 | s_CSAwallace_cska12_csa9_csa_component_fa17_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa18_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa18_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa18_and0 = s_CSAwallace_cska12_csa8_csa_component_fa18_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa18_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa18_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa18_and1 = s_CSAwallace_cska12_csa9_csa_component_fa18_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa18_or0 = s_CSAwallace_cska12_csa9_csa_component_fa18_and0 | s_CSAwallace_cska12_csa9_csa_component_fa18_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa19_xor0 = s_CSAwallace_cska12_csa8_csa_component_fa19_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa19_and0 = s_CSAwallace_cska12_csa8_csa_component_fa19_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa19_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa19_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa19_and1 = s_CSAwallace_cska12_csa9_csa_component_fa19_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa19_or0 = s_CSAwallace_cska12_csa9_csa_component_fa19_and0 | s_CSAwallace_cska12_csa9_csa_component_fa19_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa20_xor0 = s_CSAwallace_cska12_csa7_csa_component_fa20_xor1 ^ s_CSAwallace_cska12_csa8_csa_component_fa19_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa20_and0 = s_CSAwallace_cska12_csa7_csa_component_fa20_xor1 & s_CSAwallace_cska12_csa8_csa_component_fa19_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa20_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa20_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa19_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa20_and1 = s_CSAwallace_cska12_csa9_csa_component_fa20_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa19_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa20_or0 = s_CSAwallace_cska12_csa9_csa_component_fa20_and0 | s_CSAwallace_cska12_csa9_csa_component_fa20_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa21_xor0 = ~s_CSAwallace_cska12_csa7_csa_component_fa21_xor1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa21_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa21_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa20_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa21_and1 = s_CSAwallace_cska12_csa9_csa_component_fa21_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa20_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa21_or0 = s_CSAwallace_cska12_csa7_csa_component_fa21_xor1 | s_CSAwallace_cska12_csa9_csa_component_fa21_and1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa22_xor0 = ~s_CSAwallace_cska12_csa7_csa_component_fa22_xor1;
  assign s_CSAwallace_cska12_csa9_csa_component_fa22_xor1 = s_CSAwallace_cska12_csa9_csa_component_fa22_xor0 ^ s_CSAwallace_cska12_csa7_csa_component_fa21_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa22_and1 = s_CSAwallace_cska12_csa9_csa_component_fa22_xor0 & s_CSAwallace_cska12_csa7_csa_component_fa21_or0;
  assign s_CSAwallace_cska12_csa9_csa_component_fa22_or0 = s_CSAwallace_cska12_csa7_csa_component_fa22_xor1 | s_CSAwallace_cska12_csa9_csa_component_fa22_and1;
  assign s_CSAwallace_cska12_u_cska24_and_propagate00 = s_CSAwallace_cska12_and_0_0 & s_CSAwallace_cska12_csa4_csa_component_fa2_xor0;
  assign s_CSAwallace_cska12_u_cska24_and_propagate01 = s_CSAwallace_cska12_csa0_csa_component_fa1_xor0 & s_CSAwallace_cska12_csa6_csa_component_fa3_xor0;
  assign s_CSAwallace_cska12_u_cska24_and_propagate02 = s_CSAwallace_cska12_u_cska24_and_propagate00 & s_CSAwallace_cska12_u_cska24_and_propagate01;
  assign s_CSAwallace_cska12_u_cska24_mux2to10_not0 = ~s_CSAwallace_cska12_u_cska24_and_propagate02;
  assign s_CSAwallace_cska12_u_cska24_xor6 = s_CSAwallace_cska12_csa9_csa_component_fa6_xor0 ^ s_CSAwallace_cska12_csa9_csa_component_fa5_and0;
  assign s_CSAwallace_cska12_u_cska24_fa5_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa6_xor0 ^ s_CSAwallace_cska12_csa9_csa_component_fa5_and0;
  assign s_CSAwallace_cska12_u_cska24_fa5_and0 = s_CSAwallace_cska12_csa9_csa_component_fa6_xor0 & s_CSAwallace_cska12_csa9_csa_component_fa5_and0;
  assign s_CSAwallace_cska12_u_cska24_xor7 = s_CSAwallace_cska12_csa9_csa_component_fa7_xor0 ^ s_CSAwallace_cska12_csa9_csa_component_fa6_and0;
  assign s_CSAwallace_cska12_u_cska24_fa6_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa7_xor0 ^ s_CSAwallace_cska12_csa9_csa_component_fa6_and0;
  assign s_CSAwallace_cska12_u_cska24_fa6_and0 = s_CSAwallace_cska12_csa9_csa_component_fa7_xor0 & s_CSAwallace_cska12_csa9_csa_component_fa6_and0;
  assign s_CSAwallace_cska12_u_cska24_fa6_xor1 = s_CSAwallace_cska12_u_cska24_fa6_xor0 ^ s_CSAwallace_cska12_u_cska24_fa5_and0;
  assign s_CSAwallace_cska12_u_cska24_fa6_and1 = s_CSAwallace_cska12_u_cska24_fa6_xor0 & s_CSAwallace_cska12_u_cska24_fa5_and0;
  assign s_CSAwallace_cska12_u_cska24_fa6_or0 = s_CSAwallace_cska12_u_cska24_fa6_and0 | s_CSAwallace_cska12_u_cska24_fa6_and1;
  assign s_CSAwallace_cska12_u_cska24_and_propagate13 = s_CSAwallace_cska12_csa8_csa_component_fa4_xor0 & s_CSAwallace_cska12_u_cska24_xor6;
  assign s_CSAwallace_cska12_u_cska24_and_propagate14 = s_CSAwallace_cska12_csa9_csa_component_fa5_xor0 & s_CSAwallace_cska12_u_cska24_xor7;
  assign s_CSAwallace_cska12_u_cska24_and_propagate15 = s_CSAwallace_cska12_u_cska24_and_propagate13 & s_CSAwallace_cska12_u_cska24_and_propagate14;
  assign s_CSAwallace_cska12_u_cska24_mux2to11_not0 = ~s_CSAwallace_cska12_u_cska24_and_propagate15;
  assign s_CSAwallace_cska12_u_cska24_mux2to11_and1 = s_CSAwallace_cska12_u_cska24_fa6_or0 & s_CSAwallace_cska12_u_cska24_mux2to11_not0;
  assign s_CSAwallace_cska12_u_cska24_xor8 = s_CSAwallace_cska12_csa9_csa_component_fa8_xor0 ^ s_CSAwallace_cska12_csa9_csa_component_fa7_and0;
  assign s_CSAwallace_cska12_u_cska24_fa7_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa8_xor0 ^ s_CSAwallace_cska12_csa9_csa_component_fa7_and0;
  assign s_CSAwallace_cska12_u_cska24_fa7_and0 = s_CSAwallace_cska12_csa9_csa_component_fa8_xor0 & s_CSAwallace_cska12_csa9_csa_component_fa7_and0;
  assign s_CSAwallace_cska12_u_cska24_fa7_xor1 = s_CSAwallace_cska12_u_cska24_fa7_xor0 ^ s_CSAwallace_cska12_u_cska24_mux2to11_and1;
  assign s_CSAwallace_cska12_u_cska24_fa7_and1 = s_CSAwallace_cska12_u_cska24_fa7_xor0 & s_CSAwallace_cska12_u_cska24_mux2to11_and1;
  assign s_CSAwallace_cska12_u_cska24_fa7_or0 = s_CSAwallace_cska12_u_cska24_fa7_and0 | s_CSAwallace_cska12_u_cska24_fa7_and1;
  assign s_CSAwallace_cska12_u_cska24_xor9 = s_CSAwallace_cska12_csa9_csa_component_fa9_xor0 ^ s_CSAwallace_cska12_csa9_csa_component_fa8_and0;
  assign s_CSAwallace_cska12_u_cska24_fa8_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa9_xor0 ^ s_CSAwallace_cska12_csa9_csa_component_fa8_and0;
  assign s_CSAwallace_cska12_u_cska24_fa8_and0 = s_CSAwallace_cska12_csa9_csa_component_fa9_xor0 & s_CSAwallace_cska12_csa9_csa_component_fa8_and0;
  assign s_CSAwallace_cska12_u_cska24_fa8_xor1 = s_CSAwallace_cska12_u_cska24_fa8_xor0 ^ s_CSAwallace_cska12_u_cska24_fa7_or0;
  assign s_CSAwallace_cska12_u_cska24_fa8_and1 = s_CSAwallace_cska12_u_cska24_fa8_xor0 & s_CSAwallace_cska12_u_cska24_fa7_or0;
  assign s_CSAwallace_cska12_u_cska24_fa8_or0 = s_CSAwallace_cska12_u_cska24_fa8_and0 | s_CSAwallace_cska12_u_cska24_fa8_and1;
  assign s_CSAwallace_cska12_u_cska24_xor10 = s_CSAwallace_cska12_csa9_csa_component_fa10_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa9_and0;
  assign s_CSAwallace_cska12_u_cska24_fa9_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa10_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa9_and0;
  assign s_CSAwallace_cska12_u_cska24_fa9_and0 = s_CSAwallace_cska12_csa9_csa_component_fa10_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa9_and0;
  assign s_CSAwallace_cska12_u_cska24_fa9_xor1 = s_CSAwallace_cska12_u_cska24_fa9_xor0 ^ s_CSAwallace_cska12_u_cska24_fa8_or0;
  assign s_CSAwallace_cska12_u_cska24_fa9_and1 = s_CSAwallace_cska12_u_cska24_fa9_xor0 & s_CSAwallace_cska12_u_cska24_fa8_or0;
  assign s_CSAwallace_cska12_u_cska24_fa9_or0 = s_CSAwallace_cska12_u_cska24_fa9_and0 | s_CSAwallace_cska12_u_cska24_fa9_and1;
  assign s_CSAwallace_cska12_u_cska24_xor11 = s_CSAwallace_cska12_csa9_csa_component_fa11_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_u_cska24_fa10_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa11_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_u_cska24_fa10_and0 = s_CSAwallace_cska12_csa9_csa_component_fa11_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa10_or0;
  assign s_CSAwallace_cska12_u_cska24_fa10_xor1 = s_CSAwallace_cska12_u_cska24_fa10_xor0 ^ s_CSAwallace_cska12_u_cska24_fa9_or0;
  assign s_CSAwallace_cska12_u_cska24_fa10_and1 = s_CSAwallace_cska12_u_cska24_fa10_xor0 & s_CSAwallace_cska12_u_cska24_fa9_or0;
  assign s_CSAwallace_cska12_u_cska24_fa10_or0 = s_CSAwallace_cska12_u_cska24_fa10_and0 | s_CSAwallace_cska12_u_cska24_fa10_and1;
  assign s_CSAwallace_cska12_u_cska24_and_propagate26 = s_CSAwallace_cska12_u_cska24_xor8 & s_CSAwallace_cska12_u_cska24_xor10;
  assign s_CSAwallace_cska12_u_cska24_and_propagate27 = s_CSAwallace_cska12_u_cska24_xor9 & s_CSAwallace_cska12_u_cska24_xor11;
  assign s_CSAwallace_cska12_u_cska24_and_propagate28 = s_CSAwallace_cska12_u_cska24_and_propagate26 & s_CSAwallace_cska12_u_cska24_and_propagate27;
  assign s_CSAwallace_cska12_u_cska24_mux2to12_and0 = s_CSAwallace_cska12_u_cska24_mux2to11_and1 & s_CSAwallace_cska12_u_cska24_and_propagate28;
  assign s_CSAwallace_cska12_u_cska24_mux2to12_not0 = ~s_CSAwallace_cska12_u_cska24_and_propagate28;
  assign s_CSAwallace_cska12_u_cska24_mux2to12_and1 = s_CSAwallace_cska12_u_cska24_fa10_or0 & s_CSAwallace_cska12_u_cska24_mux2to12_not0;
  assign s_CSAwallace_cska12_u_cska24_mux2to12_xor0 = s_CSAwallace_cska12_u_cska24_mux2to12_and0 ^ s_CSAwallace_cska12_u_cska24_mux2to12_and1;
  assign s_CSAwallace_cska12_u_cska24_xor12 = s_CSAwallace_cska12_csa9_csa_component_fa12_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_u_cska24_fa11_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa12_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_u_cska24_fa11_and0 = s_CSAwallace_cska12_csa9_csa_component_fa12_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa11_or0;
  assign s_CSAwallace_cska12_u_cska24_fa11_xor1 = s_CSAwallace_cska12_u_cska24_fa11_xor0 ^ s_CSAwallace_cska12_u_cska24_mux2to12_xor0;
  assign s_CSAwallace_cska12_u_cska24_fa11_and1 = s_CSAwallace_cska12_u_cska24_fa11_xor0 & s_CSAwallace_cska12_u_cska24_mux2to12_xor0;
  assign s_CSAwallace_cska12_u_cska24_fa11_or0 = s_CSAwallace_cska12_u_cska24_fa11_and0 | s_CSAwallace_cska12_u_cska24_fa11_and1;
  assign s_CSAwallace_cska12_u_cska24_xor13 = s_CSAwallace_cska12_csa9_csa_component_fa13_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_u_cska24_fa12_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa13_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_u_cska24_fa12_and0 = s_CSAwallace_cska12_csa9_csa_component_fa13_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa12_or0;
  assign s_CSAwallace_cska12_u_cska24_fa12_xor1 = s_CSAwallace_cska12_u_cska24_fa12_xor0 ^ s_CSAwallace_cska12_u_cska24_fa11_or0;
  assign s_CSAwallace_cska12_u_cska24_fa12_and1 = s_CSAwallace_cska12_u_cska24_fa12_xor0 & s_CSAwallace_cska12_u_cska24_fa11_or0;
  assign s_CSAwallace_cska12_u_cska24_fa12_or0 = s_CSAwallace_cska12_u_cska24_fa12_and0 | s_CSAwallace_cska12_u_cska24_fa12_and1;
  assign s_CSAwallace_cska12_u_cska24_xor14 = s_CSAwallace_cska12_csa9_csa_component_fa14_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_u_cska24_fa13_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa14_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_u_cska24_fa13_and0 = s_CSAwallace_cska12_csa9_csa_component_fa14_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa13_or0;
  assign s_CSAwallace_cska12_u_cska24_fa13_xor1 = s_CSAwallace_cska12_u_cska24_fa13_xor0 ^ s_CSAwallace_cska12_u_cska24_fa12_or0;
  assign s_CSAwallace_cska12_u_cska24_fa13_and1 = s_CSAwallace_cska12_u_cska24_fa13_xor0 & s_CSAwallace_cska12_u_cska24_fa12_or0;
  assign s_CSAwallace_cska12_u_cska24_fa13_or0 = s_CSAwallace_cska12_u_cska24_fa13_and0 | s_CSAwallace_cska12_u_cska24_fa13_and1;
  assign s_CSAwallace_cska12_u_cska24_xor15 = s_CSAwallace_cska12_csa9_csa_component_fa15_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_u_cska24_fa14_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa15_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_u_cska24_fa14_and0 = s_CSAwallace_cska12_csa9_csa_component_fa15_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa14_or0;
  assign s_CSAwallace_cska12_u_cska24_fa14_xor1 = s_CSAwallace_cska12_u_cska24_fa14_xor0 ^ s_CSAwallace_cska12_u_cska24_fa13_or0;
  assign s_CSAwallace_cska12_u_cska24_fa14_and1 = s_CSAwallace_cska12_u_cska24_fa14_xor0 & s_CSAwallace_cska12_u_cska24_fa13_or0;
  assign s_CSAwallace_cska12_u_cska24_fa14_or0 = s_CSAwallace_cska12_u_cska24_fa14_and0 | s_CSAwallace_cska12_u_cska24_fa14_and1;
  assign s_CSAwallace_cska12_u_cska24_and_propagate39 = s_CSAwallace_cska12_u_cska24_xor12 & s_CSAwallace_cska12_u_cska24_xor14;
  assign s_CSAwallace_cska12_u_cska24_and_propagate310 = s_CSAwallace_cska12_u_cska24_xor13 & s_CSAwallace_cska12_u_cska24_xor15;
  assign s_CSAwallace_cska12_u_cska24_and_propagate311 = s_CSAwallace_cska12_u_cska24_and_propagate39 & s_CSAwallace_cska12_u_cska24_and_propagate310;
  assign s_CSAwallace_cska12_u_cska24_mux2to13_and0 = s_CSAwallace_cska12_u_cska24_mux2to12_xor0 & s_CSAwallace_cska12_u_cska24_and_propagate311;
  assign s_CSAwallace_cska12_u_cska24_mux2to13_not0 = ~s_CSAwallace_cska12_u_cska24_and_propagate311;
  assign s_CSAwallace_cska12_u_cska24_mux2to13_and1 = s_CSAwallace_cska12_u_cska24_fa14_or0 & s_CSAwallace_cska12_u_cska24_mux2to13_not0;
  assign s_CSAwallace_cska12_u_cska24_mux2to13_xor0 = s_CSAwallace_cska12_u_cska24_mux2to13_and0 ^ s_CSAwallace_cska12_u_cska24_mux2to13_and1;
  assign s_CSAwallace_cska12_u_cska24_xor16 = s_CSAwallace_cska12_csa9_csa_component_fa16_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_u_cska24_fa15_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa16_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_u_cska24_fa15_and0 = s_CSAwallace_cska12_csa9_csa_component_fa16_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa15_or0;
  assign s_CSAwallace_cska12_u_cska24_fa15_xor1 = s_CSAwallace_cska12_u_cska24_fa15_xor0 ^ s_CSAwallace_cska12_u_cska24_mux2to13_xor0;
  assign s_CSAwallace_cska12_u_cska24_fa15_and1 = s_CSAwallace_cska12_u_cska24_fa15_xor0 & s_CSAwallace_cska12_u_cska24_mux2to13_xor0;
  assign s_CSAwallace_cska12_u_cska24_fa15_or0 = s_CSAwallace_cska12_u_cska24_fa15_and0 | s_CSAwallace_cska12_u_cska24_fa15_and1;
  assign s_CSAwallace_cska12_u_cska24_xor17 = s_CSAwallace_cska12_csa9_csa_component_fa17_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_u_cska24_fa16_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa17_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_u_cska24_fa16_and0 = s_CSAwallace_cska12_csa9_csa_component_fa17_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa16_or0;
  assign s_CSAwallace_cska12_u_cska24_fa16_xor1 = s_CSAwallace_cska12_u_cska24_fa16_xor0 ^ s_CSAwallace_cska12_u_cska24_fa15_or0;
  assign s_CSAwallace_cska12_u_cska24_fa16_and1 = s_CSAwallace_cska12_u_cska24_fa16_xor0 & s_CSAwallace_cska12_u_cska24_fa15_or0;
  assign s_CSAwallace_cska12_u_cska24_fa16_or0 = s_CSAwallace_cska12_u_cska24_fa16_and0 | s_CSAwallace_cska12_u_cska24_fa16_and1;
  assign s_CSAwallace_cska12_u_cska24_xor18 = s_CSAwallace_cska12_csa9_csa_component_fa18_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_u_cska24_fa17_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa18_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_u_cska24_fa17_and0 = s_CSAwallace_cska12_csa9_csa_component_fa18_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa17_or0;
  assign s_CSAwallace_cska12_u_cska24_fa17_xor1 = s_CSAwallace_cska12_u_cska24_fa17_xor0 ^ s_CSAwallace_cska12_u_cska24_fa16_or0;
  assign s_CSAwallace_cska12_u_cska24_fa17_and1 = s_CSAwallace_cska12_u_cska24_fa17_xor0 & s_CSAwallace_cska12_u_cska24_fa16_or0;
  assign s_CSAwallace_cska12_u_cska24_fa17_or0 = s_CSAwallace_cska12_u_cska24_fa17_and0 | s_CSAwallace_cska12_u_cska24_fa17_and1;
  assign s_CSAwallace_cska12_u_cska24_xor19 = s_CSAwallace_cska12_csa9_csa_component_fa19_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_u_cska24_fa18_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa19_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_u_cska24_fa18_and0 = s_CSAwallace_cska12_csa9_csa_component_fa19_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa18_or0;
  assign s_CSAwallace_cska12_u_cska24_fa18_xor1 = s_CSAwallace_cska12_u_cska24_fa18_xor0 ^ s_CSAwallace_cska12_u_cska24_fa17_or0;
  assign s_CSAwallace_cska12_u_cska24_fa18_and1 = s_CSAwallace_cska12_u_cska24_fa18_xor0 & s_CSAwallace_cska12_u_cska24_fa17_or0;
  assign s_CSAwallace_cska12_u_cska24_fa18_or0 = s_CSAwallace_cska12_u_cska24_fa18_and0 | s_CSAwallace_cska12_u_cska24_fa18_and1;
  assign s_CSAwallace_cska12_u_cska24_and_propagate412 = s_CSAwallace_cska12_u_cska24_xor16 & s_CSAwallace_cska12_u_cska24_xor18;
  assign s_CSAwallace_cska12_u_cska24_and_propagate413 = s_CSAwallace_cska12_u_cska24_xor17 & s_CSAwallace_cska12_u_cska24_xor19;
  assign s_CSAwallace_cska12_u_cska24_and_propagate414 = s_CSAwallace_cska12_u_cska24_and_propagate412 & s_CSAwallace_cska12_u_cska24_and_propagate413;
  assign s_CSAwallace_cska12_u_cska24_mux2to14_and0 = s_CSAwallace_cska12_u_cska24_mux2to13_xor0 & s_CSAwallace_cska12_u_cska24_and_propagate414;
  assign s_CSAwallace_cska12_u_cska24_mux2to14_not0 = ~s_CSAwallace_cska12_u_cska24_and_propagate414;
  assign s_CSAwallace_cska12_u_cska24_mux2to14_and1 = s_CSAwallace_cska12_u_cska24_fa18_or0 & s_CSAwallace_cska12_u_cska24_mux2to14_not0;
  assign s_CSAwallace_cska12_u_cska24_mux2to14_xor0 = s_CSAwallace_cska12_u_cska24_mux2to14_and0 ^ s_CSAwallace_cska12_u_cska24_mux2to14_and1;
  assign s_CSAwallace_cska12_u_cska24_xor20 = s_CSAwallace_cska12_csa9_csa_component_fa20_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa19_or0;
  assign s_CSAwallace_cska12_u_cska24_fa19_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa20_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa19_or0;
  assign s_CSAwallace_cska12_u_cska24_fa19_and0 = s_CSAwallace_cska12_csa9_csa_component_fa20_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa19_or0;
  assign s_CSAwallace_cska12_u_cska24_fa19_xor1 = s_CSAwallace_cska12_u_cska24_fa19_xor0 ^ s_CSAwallace_cska12_u_cska24_mux2to14_xor0;
  assign s_CSAwallace_cska12_u_cska24_fa19_and1 = s_CSAwallace_cska12_u_cska24_fa19_xor0 & s_CSAwallace_cska12_u_cska24_mux2to14_xor0;
  assign s_CSAwallace_cska12_u_cska24_fa19_or0 = s_CSAwallace_cska12_u_cska24_fa19_and0 | s_CSAwallace_cska12_u_cska24_fa19_and1;
  assign s_CSAwallace_cska12_u_cska24_xor21 = s_CSAwallace_cska12_csa9_csa_component_fa21_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa20_or0;
  assign s_CSAwallace_cska12_u_cska24_fa20_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa21_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa20_or0;
  assign s_CSAwallace_cska12_u_cska24_fa20_and0 = s_CSAwallace_cska12_csa9_csa_component_fa21_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa20_or0;
  assign s_CSAwallace_cska12_u_cska24_fa20_xor1 = s_CSAwallace_cska12_u_cska24_fa20_xor0 ^ s_CSAwallace_cska12_u_cska24_fa19_or0;
  assign s_CSAwallace_cska12_u_cska24_fa20_and1 = s_CSAwallace_cska12_u_cska24_fa20_xor0 & s_CSAwallace_cska12_u_cska24_fa19_or0;
  assign s_CSAwallace_cska12_u_cska24_fa20_or0 = s_CSAwallace_cska12_u_cska24_fa20_and0 | s_CSAwallace_cska12_u_cska24_fa20_and1;
  assign s_CSAwallace_cska12_u_cska24_xor22 = s_CSAwallace_cska12_csa9_csa_component_fa22_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa21_or0;
  assign s_CSAwallace_cska12_u_cska24_fa21_xor0 = s_CSAwallace_cska12_csa9_csa_component_fa22_xor1 ^ s_CSAwallace_cska12_csa9_csa_component_fa21_or0;
  assign s_CSAwallace_cska12_u_cska24_fa21_and0 = s_CSAwallace_cska12_csa9_csa_component_fa22_xor1 & s_CSAwallace_cska12_csa9_csa_component_fa21_or0;
  assign s_CSAwallace_cska12_u_cska24_fa21_xor1 = s_CSAwallace_cska12_u_cska24_fa21_xor0 ^ s_CSAwallace_cska12_u_cska24_fa20_or0;
  assign s_CSAwallace_cska12_u_cska24_fa21_and1 = s_CSAwallace_cska12_u_cska24_fa21_xor0 & s_CSAwallace_cska12_u_cska24_fa20_or0;
  assign s_CSAwallace_cska12_u_cska24_fa21_or0 = s_CSAwallace_cska12_u_cska24_fa21_and0 | s_CSAwallace_cska12_u_cska24_fa21_and1;
  assign s_CSAwallace_cska12_u_cska24_xor23 = s_CSAwallace_cska12_csa7_csa_component_fa22_or0 ^ s_CSAwallace_cska12_csa9_csa_component_fa22_or0;
  assign s_CSAwallace_cska12_u_cska24_fa22_xor0 = s_CSAwallace_cska12_csa7_csa_component_fa22_or0 ^ s_CSAwallace_cska12_csa9_csa_component_fa22_or0;
  assign s_CSAwallace_cska12_u_cska24_fa22_and0 = s_CSAwallace_cska12_csa7_csa_component_fa22_or0 & s_CSAwallace_cska12_csa9_csa_component_fa22_or0;
  assign s_CSAwallace_cska12_u_cska24_fa22_xor1 = s_CSAwallace_cska12_u_cska24_fa22_xor0 ^ s_CSAwallace_cska12_u_cska24_fa21_or0;
  assign s_CSAwallace_cska12_u_cska24_fa22_and1 = s_CSAwallace_cska12_u_cska24_fa22_xor0 & s_CSAwallace_cska12_u_cska24_fa21_or0;
  assign s_CSAwallace_cska12_u_cska24_fa22_or0 = s_CSAwallace_cska12_u_cska24_fa22_and0 | s_CSAwallace_cska12_u_cska24_fa22_and1;
  assign s_CSAwallace_cska12_u_cska24_and_propagate515 = s_CSAwallace_cska12_u_cska24_xor20 & s_CSAwallace_cska12_u_cska24_xor22;
  assign s_CSAwallace_cska12_u_cska24_and_propagate516 = s_CSAwallace_cska12_u_cska24_xor21 & s_CSAwallace_cska12_u_cska24_xor23;
  assign s_CSAwallace_cska12_u_cska24_and_propagate517 = s_CSAwallace_cska12_u_cska24_and_propagate515 & s_CSAwallace_cska12_u_cska24_and_propagate516;
  assign s_CSAwallace_cska12_u_cska24_mux2to15_and0 = s_CSAwallace_cska12_u_cska24_mux2to14_xor0 & s_CSAwallace_cska12_u_cska24_and_propagate517;
  assign s_CSAwallace_cska12_u_cska24_mux2to15_not0 = ~s_CSAwallace_cska12_u_cska24_and_propagate517;
  assign s_CSAwallace_cska12_u_cska24_mux2to15_and1 = s_CSAwallace_cska12_u_cska24_fa22_or0 & s_CSAwallace_cska12_u_cska24_mux2to15_not0;
  assign s_CSAwallace_cska12_u_cska24_mux2to15_xor0 = s_CSAwallace_cska12_u_cska24_mux2to15_and0 ^ s_CSAwallace_cska12_u_cska24_mux2to15_and1;
  assign s_CSAwallace_cska12_xor0 = ~s_CSAwallace_cska12_u_cska24_fa22_xor1;

  assign s_CSAwallace_cska12_out[0] = s_CSAwallace_cska12_and_0_0;
  assign s_CSAwallace_cska12_out[1] = s_CSAwallace_cska12_csa0_csa_component_fa1_xor0;
  assign s_CSAwallace_cska12_out[2] = s_CSAwallace_cska12_csa4_csa_component_fa2_xor0;
  assign s_CSAwallace_cska12_out[3] = s_CSAwallace_cska12_csa6_csa_component_fa3_xor0;
  assign s_CSAwallace_cska12_out[4] = s_CSAwallace_cska12_csa8_csa_component_fa4_xor0;
  assign s_CSAwallace_cska12_out[5] = s_CSAwallace_cska12_csa9_csa_component_fa5_xor0;
  assign s_CSAwallace_cska12_out[6] = s_CSAwallace_cska12_u_cska24_fa5_xor0;
  assign s_CSAwallace_cska12_out[7] = s_CSAwallace_cska12_u_cska24_fa6_xor1;
  assign s_CSAwallace_cska12_out[8] = s_CSAwallace_cska12_u_cska24_fa7_xor1;
  assign s_CSAwallace_cska12_out[9] = s_CSAwallace_cska12_u_cska24_fa8_xor1;
  assign s_CSAwallace_cska12_out[10] = s_CSAwallace_cska12_u_cska24_fa9_xor1;
  assign s_CSAwallace_cska12_out[11] = s_CSAwallace_cska12_u_cska24_fa10_xor1;
  assign s_CSAwallace_cska12_out[12] = s_CSAwallace_cska12_u_cska24_fa11_xor1;
  assign s_CSAwallace_cska12_out[13] = s_CSAwallace_cska12_u_cska24_fa12_xor1;
  assign s_CSAwallace_cska12_out[14] = s_CSAwallace_cska12_u_cska24_fa13_xor1;
  assign s_CSAwallace_cska12_out[15] = s_CSAwallace_cska12_u_cska24_fa14_xor1;
  assign s_CSAwallace_cska12_out[16] = s_CSAwallace_cska12_u_cska24_fa15_xor1;
  assign s_CSAwallace_cska12_out[17] = s_CSAwallace_cska12_u_cska24_fa16_xor1;
  assign s_CSAwallace_cska12_out[18] = s_CSAwallace_cska12_u_cska24_fa17_xor1;
  assign s_CSAwallace_cska12_out[19] = s_CSAwallace_cska12_u_cska24_fa18_xor1;
  assign s_CSAwallace_cska12_out[20] = s_CSAwallace_cska12_u_cska24_fa19_xor1;
  assign s_CSAwallace_cska12_out[21] = s_CSAwallace_cska12_u_cska24_fa20_xor1;
  assign s_CSAwallace_cska12_out[22] = s_CSAwallace_cska12_u_cska24_fa21_xor1;
  assign s_CSAwallace_cska12_out[23] = s_CSAwallace_cska12_xor0;
endmodule