module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(a[0], b[0], pg_logic_or0);
  and_gate and_gate_pg_logic_and0(a[0], b[0], pg_logic_and0);
  xor_gate xor_gate_pg_logic_xor0(a[0], b[0], pg_logic_xor0);
endmodule

module h_s_cla8(input [7:0] a, input [7:0] b, output [8:0] h_s_cla8_out);
  wire [0:0] h_s_cla8_pg_logic0_or0;
  wire [0:0] h_s_cla8_pg_logic0_and0;
  wire [0:0] h_s_cla8_pg_logic0_xor0;
  wire [0:0] h_s_cla8_pg_logic1_or0;
  wire [0:0] h_s_cla8_pg_logic1_and0;
  wire [0:0] h_s_cla8_pg_logic1_xor0;
  wire [0:0] h_s_cla8_xor1;
  wire [0:0] h_s_cla8_and0;
  wire [0:0] h_s_cla8_or0;
  wire [0:0] h_s_cla8_pg_logic2_or0;
  wire [0:0] h_s_cla8_pg_logic2_and0;
  wire [0:0] h_s_cla8_pg_logic2_xor0;
  wire [0:0] h_s_cla8_xor2;
  wire [0:0] h_s_cla8_and1;
  wire [0:0] h_s_cla8_and2;
  wire [0:0] h_s_cla8_and3;
  wire [0:0] h_s_cla8_and4;
  wire [0:0] h_s_cla8_or1;
  wire [0:0] h_s_cla8_or2;
  wire [0:0] h_s_cla8_pg_logic3_or0;
  wire [0:0] h_s_cla8_pg_logic3_and0;
  wire [0:0] h_s_cla8_pg_logic3_xor0;
  wire [0:0] h_s_cla8_xor3;
  wire [0:0] h_s_cla8_and5;
  wire [0:0] h_s_cla8_and6;
  wire [0:0] h_s_cla8_and7;
  wire [0:0] h_s_cla8_and8;
  wire [0:0] h_s_cla8_and9;
  wire [0:0] h_s_cla8_and10;
  wire [0:0] h_s_cla8_and11;
  wire [0:0] h_s_cla8_or3;
  wire [0:0] h_s_cla8_or4;
  wire [0:0] h_s_cla8_or5;
  wire [0:0] h_s_cla8_pg_logic4_or0;
  wire [0:0] h_s_cla8_pg_logic4_and0;
  wire [0:0] h_s_cla8_pg_logic4_xor0;
  wire [0:0] h_s_cla8_xor4;
  wire [0:0] h_s_cla8_and12;
  wire [0:0] h_s_cla8_or6;
  wire [0:0] h_s_cla8_pg_logic5_or0;
  wire [0:0] h_s_cla8_pg_logic5_and0;
  wire [0:0] h_s_cla8_pg_logic5_xor0;
  wire [0:0] h_s_cla8_xor5;
  wire [0:0] h_s_cla8_and13;
  wire [0:0] h_s_cla8_and14;
  wire [0:0] h_s_cla8_and15;
  wire [0:0] h_s_cla8_or7;
  wire [0:0] h_s_cla8_or8;
  wire [0:0] h_s_cla8_pg_logic6_or0;
  wire [0:0] h_s_cla8_pg_logic6_and0;
  wire [0:0] h_s_cla8_pg_logic6_xor0;
  wire [0:0] h_s_cla8_xor6;
  wire [0:0] h_s_cla8_and16;
  wire [0:0] h_s_cla8_and17;
  wire [0:0] h_s_cla8_and18;
  wire [0:0] h_s_cla8_and19;
  wire [0:0] h_s_cla8_and20;
  wire [0:0] h_s_cla8_and21;
  wire [0:0] h_s_cla8_or9;
  wire [0:0] h_s_cla8_or10;
  wire [0:0] h_s_cla8_or11;
  wire [0:0] h_s_cla8_pg_logic7_or0;
  wire [0:0] h_s_cla8_pg_logic7_and0;
  wire [0:0] h_s_cla8_pg_logic7_xor0;
  wire [0:0] h_s_cla8_xor7;
  wire [0:0] h_s_cla8_and22;
  wire [0:0] h_s_cla8_and23;
  wire [0:0] h_s_cla8_and24;
  wire [0:0] h_s_cla8_and25;
  wire [0:0] h_s_cla8_and26;
  wire [0:0] h_s_cla8_and27;
  wire [0:0] h_s_cla8_and28;
  wire [0:0] h_s_cla8_and29;
  wire [0:0] h_s_cla8_and30;
  wire [0:0] h_s_cla8_and31;
  wire [0:0] h_s_cla8_or12;
  wire [0:0] h_s_cla8_or13;
  wire [0:0] h_s_cla8_or14;
  wire [0:0] h_s_cla8_or15;
  wire [0:0] h_s_cla8_xor8;
  wire [0:0] h_s_cla8_xor9;

  pg_logic pg_logic_h_s_cla8_pg_logic0_out(a[0], b[0], h_s_cla8_pg_logic0_or0, h_s_cla8_pg_logic0_and0, h_s_cla8_pg_logic0_xor0);
  pg_logic pg_logic_h_s_cla8_pg_logic1_out(a[1], b[1], h_s_cla8_pg_logic1_or0, h_s_cla8_pg_logic1_and0, h_s_cla8_pg_logic1_xor0);
  xor_gate xor_gate_h_s_cla8_xor1(h_s_cla8_pg_logic1_xor0[0], h_s_cla8_pg_logic0_and0[0], h_s_cla8_xor1);
  and_gate and_gate_h_s_cla8_and0(h_s_cla8_pg_logic0_and0[0], h_s_cla8_pg_logic1_or0[0], h_s_cla8_and0);
  or_gate or_gate_h_s_cla8_or0(h_s_cla8_pg_logic1_and0[0], h_s_cla8_and0[0], h_s_cla8_or0);
  pg_logic pg_logic_h_s_cla8_pg_logic2_out(a[2], b[2], h_s_cla8_pg_logic2_or0, h_s_cla8_pg_logic2_and0, h_s_cla8_pg_logic2_xor0);
  xor_gate xor_gate_h_s_cla8_xor2(h_s_cla8_pg_logic2_xor0[0], h_s_cla8_or0[0], h_s_cla8_xor2);
  and_gate and_gate_h_s_cla8_and1(h_s_cla8_pg_logic2_or0[0], h_s_cla8_pg_logic0_or0[0], h_s_cla8_and1);
  and_gate and_gate_h_s_cla8_and2(h_s_cla8_pg_logic0_and0[0], h_s_cla8_pg_logic2_or0[0], h_s_cla8_and2);
  and_gate and_gate_h_s_cla8_and3(h_s_cla8_and2[0], h_s_cla8_pg_logic1_or0[0], h_s_cla8_and3);
  and_gate and_gate_h_s_cla8_and4(h_s_cla8_pg_logic1_and0[0], h_s_cla8_pg_logic2_or0[0], h_s_cla8_and4);
  or_gate or_gate_h_s_cla8_or1(h_s_cla8_and3[0], h_s_cla8_and4[0], h_s_cla8_or1);
  or_gate or_gate_h_s_cla8_or2(h_s_cla8_pg_logic2_and0[0], h_s_cla8_or1[0], h_s_cla8_or2);
  pg_logic pg_logic_h_s_cla8_pg_logic3_out(a[3], b[3], h_s_cla8_pg_logic3_or0, h_s_cla8_pg_logic3_and0, h_s_cla8_pg_logic3_xor0);
  xor_gate xor_gate_h_s_cla8_xor3(h_s_cla8_pg_logic3_xor0[0], h_s_cla8_or2[0], h_s_cla8_xor3);
  and_gate and_gate_h_s_cla8_and5(h_s_cla8_pg_logic3_or0[0], h_s_cla8_pg_logic1_or0[0], h_s_cla8_and5);
  and_gate and_gate_h_s_cla8_and6(h_s_cla8_pg_logic0_and0[0], h_s_cla8_pg_logic2_or0[0], h_s_cla8_and6);
  and_gate and_gate_h_s_cla8_and7(h_s_cla8_pg_logic3_or0[0], h_s_cla8_pg_logic1_or0[0], h_s_cla8_and7);
  and_gate and_gate_h_s_cla8_and8(h_s_cla8_and6[0], h_s_cla8_and7[0], h_s_cla8_and8);
  and_gate and_gate_h_s_cla8_and9(h_s_cla8_pg_logic1_and0[0], h_s_cla8_pg_logic3_or0[0], h_s_cla8_and9);
  and_gate and_gate_h_s_cla8_and10(h_s_cla8_and9[0], h_s_cla8_pg_logic2_or0[0], h_s_cla8_and10);
  and_gate and_gate_h_s_cla8_and11(h_s_cla8_pg_logic2_and0[0], h_s_cla8_pg_logic3_or0[0], h_s_cla8_and11);
  or_gate or_gate_h_s_cla8_or3(h_s_cla8_and8[0], h_s_cla8_and11[0], h_s_cla8_or3);
  or_gate or_gate_h_s_cla8_or4(h_s_cla8_and10[0], h_s_cla8_or3[0], h_s_cla8_or4);
  or_gate or_gate_h_s_cla8_or5(h_s_cla8_pg_logic3_and0[0], h_s_cla8_or4[0], h_s_cla8_or5);
  pg_logic pg_logic_h_s_cla8_pg_logic4_out(a[4], b[4], h_s_cla8_pg_logic4_or0, h_s_cla8_pg_logic4_and0, h_s_cla8_pg_logic4_xor0);
  xor_gate xor_gate_h_s_cla8_xor4(h_s_cla8_pg_logic4_xor0[0], h_s_cla8_or5[0], h_s_cla8_xor4);
  and_gate and_gate_h_s_cla8_and12(h_s_cla8_or5[0], h_s_cla8_pg_logic4_or0[0], h_s_cla8_and12);
  or_gate or_gate_h_s_cla8_or6(h_s_cla8_pg_logic4_and0[0], h_s_cla8_and12[0], h_s_cla8_or6);
  pg_logic pg_logic_h_s_cla8_pg_logic5_out(a[5], b[5], h_s_cla8_pg_logic5_or0, h_s_cla8_pg_logic5_and0, h_s_cla8_pg_logic5_xor0);
  xor_gate xor_gate_h_s_cla8_xor5(h_s_cla8_pg_logic5_xor0[0], h_s_cla8_or6[0], h_s_cla8_xor5);
  and_gate and_gate_h_s_cla8_and13(h_s_cla8_or5[0], h_s_cla8_pg_logic5_or0[0], h_s_cla8_and13);
  and_gate and_gate_h_s_cla8_and14(h_s_cla8_and13[0], h_s_cla8_pg_logic4_or0[0], h_s_cla8_and14);
  and_gate and_gate_h_s_cla8_and15(h_s_cla8_pg_logic4_and0[0], h_s_cla8_pg_logic5_or0[0], h_s_cla8_and15);
  or_gate or_gate_h_s_cla8_or7(h_s_cla8_and14[0], h_s_cla8_and15[0], h_s_cla8_or7);
  or_gate or_gate_h_s_cla8_or8(h_s_cla8_pg_logic5_and0[0], h_s_cla8_or7[0], h_s_cla8_or8);
  pg_logic pg_logic_h_s_cla8_pg_logic6_out(a[6], b[6], h_s_cla8_pg_logic6_or0, h_s_cla8_pg_logic6_and0, h_s_cla8_pg_logic6_xor0);
  xor_gate xor_gate_h_s_cla8_xor6(h_s_cla8_pg_logic6_xor0[0], h_s_cla8_or8[0], h_s_cla8_xor6);
  and_gate and_gate_h_s_cla8_and16(h_s_cla8_or5[0], h_s_cla8_pg_logic5_or0[0], h_s_cla8_and16);
  and_gate and_gate_h_s_cla8_and17(h_s_cla8_pg_logic6_or0[0], h_s_cla8_pg_logic4_or0[0], h_s_cla8_and17);
  and_gate and_gate_h_s_cla8_and18(h_s_cla8_and16[0], h_s_cla8_and17[0], h_s_cla8_and18);
  and_gate and_gate_h_s_cla8_and19(h_s_cla8_pg_logic4_and0[0], h_s_cla8_pg_logic6_or0[0], h_s_cla8_and19);
  and_gate and_gate_h_s_cla8_and20(h_s_cla8_and19[0], h_s_cla8_pg_logic5_or0[0], h_s_cla8_and20);
  and_gate and_gate_h_s_cla8_and21(h_s_cla8_pg_logic5_and0[0], h_s_cla8_pg_logic6_or0[0], h_s_cla8_and21);
  or_gate or_gate_h_s_cla8_or9(h_s_cla8_and18[0], h_s_cla8_and20[0], h_s_cla8_or9);
  or_gate or_gate_h_s_cla8_or10(h_s_cla8_or9[0], h_s_cla8_and21[0], h_s_cla8_or10);
  or_gate or_gate_h_s_cla8_or11(h_s_cla8_pg_logic6_and0[0], h_s_cla8_or10[0], h_s_cla8_or11);
  pg_logic pg_logic_h_s_cla8_pg_logic7_out(a[7], b[7], h_s_cla8_pg_logic7_or0, h_s_cla8_pg_logic7_and0, h_s_cla8_pg_logic7_xor0);
  xor_gate xor_gate_h_s_cla8_xor7(h_s_cla8_pg_logic7_xor0[0], h_s_cla8_or11[0], h_s_cla8_xor7);
  and_gate and_gate_h_s_cla8_and22(h_s_cla8_or5[0], h_s_cla8_pg_logic6_or0[0], h_s_cla8_and22);
  and_gate and_gate_h_s_cla8_and23(h_s_cla8_pg_logic7_or0[0], h_s_cla8_pg_logic5_or0[0], h_s_cla8_and23);
  and_gate and_gate_h_s_cla8_and24(h_s_cla8_and22[0], h_s_cla8_and23[0], h_s_cla8_and24);
  and_gate and_gate_h_s_cla8_and25(h_s_cla8_and24[0], h_s_cla8_pg_logic4_or0[0], h_s_cla8_and25);
  and_gate and_gate_h_s_cla8_and26(h_s_cla8_pg_logic4_and0[0], h_s_cla8_pg_logic6_or0[0], h_s_cla8_and26);
  and_gate and_gate_h_s_cla8_and27(h_s_cla8_pg_logic7_or0[0], h_s_cla8_pg_logic5_or0[0], h_s_cla8_and27);
  and_gate and_gate_h_s_cla8_and28(h_s_cla8_and26[0], h_s_cla8_and27[0], h_s_cla8_and28);
  and_gate and_gate_h_s_cla8_and29(h_s_cla8_pg_logic5_and0[0], h_s_cla8_pg_logic7_or0[0], h_s_cla8_and29);
  and_gate and_gate_h_s_cla8_and30(h_s_cla8_and29[0], h_s_cla8_pg_logic6_or0[0], h_s_cla8_and30);
  and_gate and_gate_h_s_cla8_and31(h_s_cla8_pg_logic6_and0[0], h_s_cla8_pg_logic7_or0[0], h_s_cla8_and31);
  or_gate or_gate_h_s_cla8_or12(h_s_cla8_and25[0], h_s_cla8_and30[0], h_s_cla8_or12);
  or_gate or_gate_h_s_cla8_or13(h_s_cla8_and28[0], h_s_cla8_and31[0], h_s_cla8_or13);
  or_gate or_gate_h_s_cla8_or14(h_s_cla8_or12[0], h_s_cla8_or13[0], h_s_cla8_or14);
  or_gate or_gate_h_s_cla8_or15(h_s_cla8_pg_logic7_and0[0], h_s_cla8_or14[0], h_s_cla8_or15);
  xor_gate xor_gate_h_s_cla8_xor8(a[7], b[7], h_s_cla8_xor8);
  xor_gate xor_gate_h_s_cla8_xor9(h_s_cla8_xor8[0], h_s_cla8_or15[0], h_s_cla8_xor9);

  assign h_s_cla8_out[0] = h_s_cla8_pg_logic0_xor0[0];
  assign h_s_cla8_out[1] = h_s_cla8_xor1[0];
  assign h_s_cla8_out[2] = h_s_cla8_xor2[0];
  assign h_s_cla8_out[3] = h_s_cla8_xor3[0];
  assign h_s_cla8_out[4] = h_s_cla8_xor4[0];
  assign h_s_cla8_out[5] = h_s_cla8_xor5[0];
  assign h_s_cla8_out[6] = h_s_cla8_xor6[0];
  assign h_s_cla8_out[7] = h_s_cla8_xor7[0];
  assign h_s_cla8_out[8] = h_s_cla8_xor9[0];
endmodule