module f_u_wallace_rca12(input [11:0] a, input [11:0] b, output [23:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire f_u_wallace_rca12_and_2_0_a_2;
  wire f_u_wallace_rca12_and_2_0_b_0;
  wire f_u_wallace_rca12_and_2_0_y0;
  wire f_u_wallace_rca12_and_1_1_a_1;
  wire f_u_wallace_rca12_and_1_1_b_1;
  wire f_u_wallace_rca12_and_1_1_y0;
  wire f_u_wallace_rca12_ha0_f_u_wallace_rca12_and_2_0_y0;
  wire f_u_wallace_rca12_ha0_f_u_wallace_rca12_and_1_1_y0;
  wire f_u_wallace_rca12_ha0_y0;
  wire f_u_wallace_rca12_ha0_y1;
  wire f_u_wallace_rca12_and_3_0_a_3;
  wire f_u_wallace_rca12_and_3_0_b_0;
  wire f_u_wallace_rca12_and_3_0_y0;
  wire f_u_wallace_rca12_and_2_1_a_2;
  wire f_u_wallace_rca12_and_2_1_b_1;
  wire f_u_wallace_rca12_and_2_1_y0;
  wire f_u_wallace_rca12_fa0_f_u_wallace_rca12_ha0_y1;
  wire f_u_wallace_rca12_fa0_f_u_wallace_rca12_and_3_0_y0;
  wire f_u_wallace_rca12_fa0_y0;
  wire f_u_wallace_rca12_fa0_y1;
  wire f_u_wallace_rca12_fa0_f_u_wallace_rca12_and_2_1_y0;
  wire f_u_wallace_rca12_fa0_y2;
  wire f_u_wallace_rca12_fa0_y3;
  wire f_u_wallace_rca12_fa0_y4;
  wire f_u_wallace_rca12_and_4_0_a_4;
  wire f_u_wallace_rca12_and_4_0_b_0;
  wire f_u_wallace_rca12_and_4_0_y0;
  wire f_u_wallace_rca12_and_3_1_a_3;
  wire f_u_wallace_rca12_and_3_1_b_1;
  wire f_u_wallace_rca12_and_3_1_y0;
  wire f_u_wallace_rca12_fa1_f_u_wallace_rca12_fa0_y4;
  wire f_u_wallace_rca12_fa1_f_u_wallace_rca12_and_4_0_y0;
  wire f_u_wallace_rca12_fa1_y0;
  wire f_u_wallace_rca12_fa1_y1;
  wire f_u_wallace_rca12_fa1_f_u_wallace_rca12_and_3_1_y0;
  wire f_u_wallace_rca12_fa1_y2;
  wire f_u_wallace_rca12_fa1_y3;
  wire f_u_wallace_rca12_fa1_y4;
  wire f_u_wallace_rca12_and_5_0_a_5;
  wire f_u_wallace_rca12_and_5_0_b_0;
  wire f_u_wallace_rca12_and_5_0_y0;
  wire f_u_wallace_rca12_and_4_1_a_4;
  wire f_u_wallace_rca12_and_4_1_b_1;
  wire f_u_wallace_rca12_and_4_1_y0;
  wire f_u_wallace_rca12_fa2_f_u_wallace_rca12_fa1_y4;
  wire f_u_wallace_rca12_fa2_f_u_wallace_rca12_and_5_0_y0;
  wire f_u_wallace_rca12_fa2_y0;
  wire f_u_wallace_rca12_fa2_y1;
  wire f_u_wallace_rca12_fa2_f_u_wallace_rca12_and_4_1_y0;
  wire f_u_wallace_rca12_fa2_y2;
  wire f_u_wallace_rca12_fa2_y3;
  wire f_u_wallace_rca12_fa2_y4;
  wire f_u_wallace_rca12_and_6_0_a_6;
  wire f_u_wallace_rca12_and_6_0_b_0;
  wire f_u_wallace_rca12_and_6_0_y0;
  wire f_u_wallace_rca12_and_5_1_a_5;
  wire f_u_wallace_rca12_and_5_1_b_1;
  wire f_u_wallace_rca12_and_5_1_y0;
  wire f_u_wallace_rca12_fa3_f_u_wallace_rca12_fa2_y4;
  wire f_u_wallace_rca12_fa3_f_u_wallace_rca12_and_6_0_y0;
  wire f_u_wallace_rca12_fa3_y0;
  wire f_u_wallace_rca12_fa3_y1;
  wire f_u_wallace_rca12_fa3_f_u_wallace_rca12_and_5_1_y0;
  wire f_u_wallace_rca12_fa3_y2;
  wire f_u_wallace_rca12_fa3_y3;
  wire f_u_wallace_rca12_fa3_y4;
  wire f_u_wallace_rca12_and_7_0_a_7;
  wire f_u_wallace_rca12_and_7_0_b_0;
  wire f_u_wallace_rca12_and_7_0_y0;
  wire f_u_wallace_rca12_and_6_1_a_6;
  wire f_u_wallace_rca12_and_6_1_b_1;
  wire f_u_wallace_rca12_and_6_1_y0;
  wire f_u_wallace_rca12_fa4_f_u_wallace_rca12_fa3_y4;
  wire f_u_wallace_rca12_fa4_f_u_wallace_rca12_and_7_0_y0;
  wire f_u_wallace_rca12_fa4_y0;
  wire f_u_wallace_rca12_fa4_y1;
  wire f_u_wallace_rca12_fa4_f_u_wallace_rca12_and_6_1_y0;
  wire f_u_wallace_rca12_fa4_y2;
  wire f_u_wallace_rca12_fa4_y3;
  wire f_u_wallace_rca12_fa4_y4;
  wire f_u_wallace_rca12_and_8_0_a_8;
  wire f_u_wallace_rca12_and_8_0_b_0;
  wire f_u_wallace_rca12_and_8_0_y0;
  wire f_u_wallace_rca12_and_7_1_a_7;
  wire f_u_wallace_rca12_and_7_1_b_1;
  wire f_u_wallace_rca12_and_7_1_y0;
  wire f_u_wallace_rca12_fa5_f_u_wallace_rca12_fa4_y4;
  wire f_u_wallace_rca12_fa5_f_u_wallace_rca12_and_8_0_y0;
  wire f_u_wallace_rca12_fa5_y0;
  wire f_u_wallace_rca12_fa5_y1;
  wire f_u_wallace_rca12_fa5_f_u_wallace_rca12_and_7_1_y0;
  wire f_u_wallace_rca12_fa5_y2;
  wire f_u_wallace_rca12_fa5_y3;
  wire f_u_wallace_rca12_fa5_y4;
  wire f_u_wallace_rca12_and_9_0_a_9;
  wire f_u_wallace_rca12_and_9_0_b_0;
  wire f_u_wallace_rca12_and_9_0_y0;
  wire f_u_wallace_rca12_and_8_1_a_8;
  wire f_u_wallace_rca12_and_8_1_b_1;
  wire f_u_wallace_rca12_and_8_1_y0;
  wire f_u_wallace_rca12_fa6_f_u_wallace_rca12_fa5_y4;
  wire f_u_wallace_rca12_fa6_f_u_wallace_rca12_and_9_0_y0;
  wire f_u_wallace_rca12_fa6_y0;
  wire f_u_wallace_rca12_fa6_y1;
  wire f_u_wallace_rca12_fa6_f_u_wallace_rca12_and_8_1_y0;
  wire f_u_wallace_rca12_fa6_y2;
  wire f_u_wallace_rca12_fa6_y3;
  wire f_u_wallace_rca12_fa6_y4;
  wire f_u_wallace_rca12_and_10_0_a_10;
  wire f_u_wallace_rca12_and_10_0_b_0;
  wire f_u_wallace_rca12_and_10_0_y0;
  wire f_u_wallace_rca12_and_9_1_a_9;
  wire f_u_wallace_rca12_and_9_1_b_1;
  wire f_u_wallace_rca12_and_9_1_y0;
  wire f_u_wallace_rca12_fa7_f_u_wallace_rca12_fa6_y4;
  wire f_u_wallace_rca12_fa7_f_u_wallace_rca12_and_10_0_y0;
  wire f_u_wallace_rca12_fa7_y0;
  wire f_u_wallace_rca12_fa7_y1;
  wire f_u_wallace_rca12_fa7_f_u_wallace_rca12_and_9_1_y0;
  wire f_u_wallace_rca12_fa7_y2;
  wire f_u_wallace_rca12_fa7_y3;
  wire f_u_wallace_rca12_fa7_y4;
  wire f_u_wallace_rca12_and_11_0_a_11;
  wire f_u_wallace_rca12_and_11_0_b_0;
  wire f_u_wallace_rca12_and_11_0_y0;
  wire f_u_wallace_rca12_and_10_1_a_10;
  wire f_u_wallace_rca12_and_10_1_b_1;
  wire f_u_wallace_rca12_and_10_1_y0;
  wire f_u_wallace_rca12_fa8_f_u_wallace_rca12_fa7_y4;
  wire f_u_wallace_rca12_fa8_f_u_wallace_rca12_and_11_0_y0;
  wire f_u_wallace_rca12_fa8_y0;
  wire f_u_wallace_rca12_fa8_y1;
  wire f_u_wallace_rca12_fa8_f_u_wallace_rca12_and_10_1_y0;
  wire f_u_wallace_rca12_fa8_y2;
  wire f_u_wallace_rca12_fa8_y3;
  wire f_u_wallace_rca12_fa8_y4;
  wire f_u_wallace_rca12_and_11_1_a_11;
  wire f_u_wallace_rca12_and_11_1_b_1;
  wire f_u_wallace_rca12_and_11_1_y0;
  wire f_u_wallace_rca12_and_10_2_a_10;
  wire f_u_wallace_rca12_and_10_2_b_2;
  wire f_u_wallace_rca12_and_10_2_y0;
  wire f_u_wallace_rca12_fa9_f_u_wallace_rca12_fa8_y4;
  wire f_u_wallace_rca12_fa9_f_u_wallace_rca12_and_11_1_y0;
  wire f_u_wallace_rca12_fa9_y0;
  wire f_u_wallace_rca12_fa9_y1;
  wire f_u_wallace_rca12_fa9_f_u_wallace_rca12_and_10_2_y0;
  wire f_u_wallace_rca12_fa9_y2;
  wire f_u_wallace_rca12_fa9_y3;
  wire f_u_wallace_rca12_fa9_y4;
  wire f_u_wallace_rca12_and_11_2_a_11;
  wire f_u_wallace_rca12_and_11_2_b_2;
  wire f_u_wallace_rca12_and_11_2_y0;
  wire f_u_wallace_rca12_and_10_3_a_10;
  wire f_u_wallace_rca12_and_10_3_b_3;
  wire f_u_wallace_rca12_and_10_3_y0;
  wire f_u_wallace_rca12_fa10_f_u_wallace_rca12_fa9_y4;
  wire f_u_wallace_rca12_fa10_f_u_wallace_rca12_and_11_2_y0;
  wire f_u_wallace_rca12_fa10_y0;
  wire f_u_wallace_rca12_fa10_y1;
  wire f_u_wallace_rca12_fa10_f_u_wallace_rca12_and_10_3_y0;
  wire f_u_wallace_rca12_fa10_y2;
  wire f_u_wallace_rca12_fa10_y3;
  wire f_u_wallace_rca12_fa10_y4;
  wire f_u_wallace_rca12_and_11_3_a_11;
  wire f_u_wallace_rca12_and_11_3_b_3;
  wire f_u_wallace_rca12_and_11_3_y0;
  wire f_u_wallace_rca12_and_10_4_a_10;
  wire f_u_wallace_rca12_and_10_4_b_4;
  wire f_u_wallace_rca12_and_10_4_y0;
  wire f_u_wallace_rca12_fa11_f_u_wallace_rca12_fa10_y4;
  wire f_u_wallace_rca12_fa11_f_u_wallace_rca12_and_11_3_y0;
  wire f_u_wallace_rca12_fa11_y0;
  wire f_u_wallace_rca12_fa11_y1;
  wire f_u_wallace_rca12_fa11_f_u_wallace_rca12_and_10_4_y0;
  wire f_u_wallace_rca12_fa11_y2;
  wire f_u_wallace_rca12_fa11_y3;
  wire f_u_wallace_rca12_fa11_y4;
  wire f_u_wallace_rca12_and_11_4_a_11;
  wire f_u_wallace_rca12_and_11_4_b_4;
  wire f_u_wallace_rca12_and_11_4_y0;
  wire f_u_wallace_rca12_and_10_5_a_10;
  wire f_u_wallace_rca12_and_10_5_b_5;
  wire f_u_wallace_rca12_and_10_5_y0;
  wire f_u_wallace_rca12_fa12_f_u_wallace_rca12_fa11_y4;
  wire f_u_wallace_rca12_fa12_f_u_wallace_rca12_and_11_4_y0;
  wire f_u_wallace_rca12_fa12_y0;
  wire f_u_wallace_rca12_fa12_y1;
  wire f_u_wallace_rca12_fa12_f_u_wallace_rca12_and_10_5_y0;
  wire f_u_wallace_rca12_fa12_y2;
  wire f_u_wallace_rca12_fa12_y3;
  wire f_u_wallace_rca12_fa12_y4;
  wire f_u_wallace_rca12_and_11_5_a_11;
  wire f_u_wallace_rca12_and_11_5_b_5;
  wire f_u_wallace_rca12_and_11_5_y0;
  wire f_u_wallace_rca12_and_10_6_a_10;
  wire f_u_wallace_rca12_and_10_6_b_6;
  wire f_u_wallace_rca12_and_10_6_y0;
  wire f_u_wallace_rca12_fa13_f_u_wallace_rca12_fa12_y4;
  wire f_u_wallace_rca12_fa13_f_u_wallace_rca12_and_11_5_y0;
  wire f_u_wallace_rca12_fa13_y0;
  wire f_u_wallace_rca12_fa13_y1;
  wire f_u_wallace_rca12_fa13_f_u_wallace_rca12_and_10_6_y0;
  wire f_u_wallace_rca12_fa13_y2;
  wire f_u_wallace_rca12_fa13_y3;
  wire f_u_wallace_rca12_fa13_y4;
  wire f_u_wallace_rca12_and_11_6_a_11;
  wire f_u_wallace_rca12_and_11_6_b_6;
  wire f_u_wallace_rca12_and_11_6_y0;
  wire f_u_wallace_rca12_and_10_7_a_10;
  wire f_u_wallace_rca12_and_10_7_b_7;
  wire f_u_wallace_rca12_and_10_7_y0;
  wire f_u_wallace_rca12_fa14_f_u_wallace_rca12_fa13_y4;
  wire f_u_wallace_rca12_fa14_f_u_wallace_rca12_and_11_6_y0;
  wire f_u_wallace_rca12_fa14_y0;
  wire f_u_wallace_rca12_fa14_y1;
  wire f_u_wallace_rca12_fa14_f_u_wallace_rca12_and_10_7_y0;
  wire f_u_wallace_rca12_fa14_y2;
  wire f_u_wallace_rca12_fa14_y3;
  wire f_u_wallace_rca12_fa14_y4;
  wire f_u_wallace_rca12_and_11_7_a_11;
  wire f_u_wallace_rca12_and_11_7_b_7;
  wire f_u_wallace_rca12_and_11_7_y0;
  wire f_u_wallace_rca12_and_10_8_a_10;
  wire f_u_wallace_rca12_and_10_8_b_8;
  wire f_u_wallace_rca12_and_10_8_y0;
  wire f_u_wallace_rca12_fa15_f_u_wallace_rca12_fa14_y4;
  wire f_u_wallace_rca12_fa15_f_u_wallace_rca12_and_11_7_y0;
  wire f_u_wallace_rca12_fa15_y0;
  wire f_u_wallace_rca12_fa15_y1;
  wire f_u_wallace_rca12_fa15_f_u_wallace_rca12_and_10_8_y0;
  wire f_u_wallace_rca12_fa15_y2;
  wire f_u_wallace_rca12_fa15_y3;
  wire f_u_wallace_rca12_fa15_y4;
  wire f_u_wallace_rca12_and_11_8_a_11;
  wire f_u_wallace_rca12_and_11_8_b_8;
  wire f_u_wallace_rca12_and_11_8_y0;
  wire f_u_wallace_rca12_and_10_9_a_10;
  wire f_u_wallace_rca12_and_10_9_b_9;
  wire f_u_wallace_rca12_and_10_9_y0;
  wire f_u_wallace_rca12_fa16_f_u_wallace_rca12_fa15_y4;
  wire f_u_wallace_rca12_fa16_f_u_wallace_rca12_and_11_8_y0;
  wire f_u_wallace_rca12_fa16_y0;
  wire f_u_wallace_rca12_fa16_y1;
  wire f_u_wallace_rca12_fa16_f_u_wallace_rca12_and_10_9_y0;
  wire f_u_wallace_rca12_fa16_y2;
  wire f_u_wallace_rca12_fa16_y3;
  wire f_u_wallace_rca12_fa16_y4;
  wire f_u_wallace_rca12_and_11_9_a_11;
  wire f_u_wallace_rca12_and_11_9_b_9;
  wire f_u_wallace_rca12_and_11_9_y0;
  wire f_u_wallace_rca12_and_10_10_a_10;
  wire f_u_wallace_rca12_and_10_10_b_10;
  wire f_u_wallace_rca12_and_10_10_y0;
  wire f_u_wallace_rca12_fa17_f_u_wallace_rca12_fa16_y4;
  wire f_u_wallace_rca12_fa17_f_u_wallace_rca12_and_11_9_y0;
  wire f_u_wallace_rca12_fa17_y0;
  wire f_u_wallace_rca12_fa17_y1;
  wire f_u_wallace_rca12_fa17_f_u_wallace_rca12_and_10_10_y0;
  wire f_u_wallace_rca12_fa17_y2;
  wire f_u_wallace_rca12_fa17_y3;
  wire f_u_wallace_rca12_fa17_y4;
  wire f_u_wallace_rca12_and_1_2_a_1;
  wire f_u_wallace_rca12_and_1_2_b_2;
  wire f_u_wallace_rca12_and_1_2_y0;
  wire f_u_wallace_rca12_and_0_3_a_0;
  wire f_u_wallace_rca12_and_0_3_b_3;
  wire f_u_wallace_rca12_and_0_3_y0;
  wire f_u_wallace_rca12_ha1_f_u_wallace_rca12_and_1_2_y0;
  wire f_u_wallace_rca12_ha1_f_u_wallace_rca12_and_0_3_y0;
  wire f_u_wallace_rca12_ha1_y0;
  wire f_u_wallace_rca12_ha1_y1;
  wire f_u_wallace_rca12_and_2_2_a_2;
  wire f_u_wallace_rca12_and_2_2_b_2;
  wire f_u_wallace_rca12_and_2_2_y0;
  wire f_u_wallace_rca12_and_1_3_a_1;
  wire f_u_wallace_rca12_and_1_3_b_3;
  wire f_u_wallace_rca12_and_1_3_y0;
  wire f_u_wallace_rca12_fa18_f_u_wallace_rca12_ha1_y1;
  wire f_u_wallace_rca12_fa18_f_u_wallace_rca12_and_2_2_y0;
  wire f_u_wallace_rca12_fa18_y0;
  wire f_u_wallace_rca12_fa18_y1;
  wire f_u_wallace_rca12_fa18_f_u_wallace_rca12_and_1_3_y0;
  wire f_u_wallace_rca12_fa18_y2;
  wire f_u_wallace_rca12_fa18_y3;
  wire f_u_wallace_rca12_fa18_y4;
  wire f_u_wallace_rca12_and_3_2_a_3;
  wire f_u_wallace_rca12_and_3_2_b_2;
  wire f_u_wallace_rca12_and_3_2_y0;
  wire f_u_wallace_rca12_and_2_3_a_2;
  wire f_u_wallace_rca12_and_2_3_b_3;
  wire f_u_wallace_rca12_and_2_3_y0;
  wire f_u_wallace_rca12_fa19_f_u_wallace_rca12_fa18_y4;
  wire f_u_wallace_rca12_fa19_f_u_wallace_rca12_and_3_2_y0;
  wire f_u_wallace_rca12_fa19_y0;
  wire f_u_wallace_rca12_fa19_y1;
  wire f_u_wallace_rca12_fa19_f_u_wallace_rca12_and_2_3_y0;
  wire f_u_wallace_rca12_fa19_y2;
  wire f_u_wallace_rca12_fa19_y3;
  wire f_u_wallace_rca12_fa19_y4;
  wire f_u_wallace_rca12_and_4_2_a_4;
  wire f_u_wallace_rca12_and_4_2_b_2;
  wire f_u_wallace_rca12_and_4_2_y0;
  wire f_u_wallace_rca12_and_3_3_a_3;
  wire f_u_wallace_rca12_and_3_3_b_3;
  wire f_u_wallace_rca12_and_3_3_y0;
  wire f_u_wallace_rca12_fa20_f_u_wallace_rca12_fa19_y4;
  wire f_u_wallace_rca12_fa20_f_u_wallace_rca12_and_4_2_y0;
  wire f_u_wallace_rca12_fa20_y0;
  wire f_u_wallace_rca12_fa20_y1;
  wire f_u_wallace_rca12_fa20_f_u_wallace_rca12_and_3_3_y0;
  wire f_u_wallace_rca12_fa20_y2;
  wire f_u_wallace_rca12_fa20_y3;
  wire f_u_wallace_rca12_fa20_y4;
  wire f_u_wallace_rca12_and_5_2_a_5;
  wire f_u_wallace_rca12_and_5_2_b_2;
  wire f_u_wallace_rca12_and_5_2_y0;
  wire f_u_wallace_rca12_and_4_3_a_4;
  wire f_u_wallace_rca12_and_4_3_b_3;
  wire f_u_wallace_rca12_and_4_3_y0;
  wire f_u_wallace_rca12_fa21_f_u_wallace_rca12_fa20_y4;
  wire f_u_wallace_rca12_fa21_f_u_wallace_rca12_and_5_2_y0;
  wire f_u_wallace_rca12_fa21_y0;
  wire f_u_wallace_rca12_fa21_y1;
  wire f_u_wallace_rca12_fa21_f_u_wallace_rca12_and_4_3_y0;
  wire f_u_wallace_rca12_fa21_y2;
  wire f_u_wallace_rca12_fa21_y3;
  wire f_u_wallace_rca12_fa21_y4;
  wire f_u_wallace_rca12_and_6_2_a_6;
  wire f_u_wallace_rca12_and_6_2_b_2;
  wire f_u_wallace_rca12_and_6_2_y0;
  wire f_u_wallace_rca12_and_5_3_a_5;
  wire f_u_wallace_rca12_and_5_3_b_3;
  wire f_u_wallace_rca12_and_5_3_y0;
  wire f_u_wallace_rca12_fa22_f_u_wallace_rca12_fa21_y4;
  wire f_u_wallace_rca12_fa22_f_u_wallace_rca12_and_6_2_y0;
  wire f_u_wallace_rca12_fa22_y0;
  wire f_u_wallace_rca12_fa22_y1;
  wire f_u_wallace_rca12_fa22_f_u_wallace_rca12_and_5_3_y0;
  wire f_u_wallace_rca12_fa22_y2;
  wire f_u_wallace_rca12_fa22_y3;
  wire f_u_wallace_rca12_fa22_y4;
  wire f_u_wallace_rca12_and_7_2_a_7;
  wire f_u_wallace_rca12_and_7_2_b_2;
  wire f_u_wallace_rca12_and_7_2_y0;
  wire f_u_wallace_rca12_and_6_3_a_6;
  wire f_u_wallace_rca12_and_6_3_b_3;
  wire f_u_wallace_rca12_and_6_3_y0;
  wire f_u_wallace_rca12_fa23_f_u_wallace_rca12_fa22_y4;
  wire f_u_wallace_rca12_fa23_f_u_wallace_rca12_and_7_2_y0;
  wire f_u_wallace_rca12_fa23_y0;
  wire f_u_wallace_rca12_fa23_y1;
  wire f_u_wallace_rca12_fa23_f_u_wallace_rca12_and_6_3_y0;
  wire f_u_wallace_rca12_fa23_y2;
  wire f_u_wallace_rca12_fa23_y3;
  wire f_u_wallace_rca12_fa23_y4;
  wire f_u_wallace_rca12_and_8_2_a_8;
  wire f_u_wallace_rca12_and_8_2_b_2;
  wire f_u_wallace_rca12_and_8_2_y0;
  wire f_u_wallace_rca12_and_7_3_a_7;
  wire f_u_wallace_rca12_and_7_3_b_3;
  wire f_u_wallace_rca12_and_7_3_y0;
  wire f_u_wallace_rca12_fa24_f_u_wallace_rca12_fa23_y4;
  wire f_u_wallace_rca12_fa24_f_u_wallace_rca12_and_8_2_y0;
  wire f_u_wallace_rca12_fa24_y0;
  wire f_u_wallace_rca12_fa24_y1;
  wire f_u_wallace_rca12_fa24_f_u_wallace_rca12_and_7_3_y0;
  wire f_u_wallace_rca12_fa24_y2;
  wire f_u_wallace_rca12_fa24_y3;
  wire f_u_wallace_rca12_fa24_y4;
  wire f_u_wallace_rca12_and_9_2_a_9;
  wire f_u_wallace_rca12_and_9_2_b_2;
  wire f_u_wallace_rca12_and_9_2_y0;
  wire f_u_wallace_rca12_and_8_3_a_8;
  wire f_u_wallace_rca12_and_8_3_b_3;
  wire f_u_wallace_rca12_and_8_3_y0;
  wire f_u_wallace_rca12_fa25_f_u_wallace_rca12_fa24_y4;
  wire f_u_wallace_rca12_fa25_f_u_wallace_rca12_and_9_2_y0;
  wire f_u_wallace_rca12_fa25_y0;
  wire f_u_wallace_rca12_fa25_y1;
  wire f_u_wallace_rca12_fa25_f_u_wallace_rca12_and_8_3_y0;
  wire f_u_wallace_rca12_fa25_y2;
  wire f_u_wallace_rca12_fa25_y3;
  wire f_u_wallace_rca12_fa25_y4;
  wire f_u_wallace_rca12_and_9_3_a_9;
  wire f_u_wallace_rca12_and_9_3_b_3;
  wire f_u_wallace_rca12_and_9_3_y0;
  wire f_u_wallace_rca12_and_8_4_a_8;
  wire f_u_wallace_rca12_and_8_4_b_4;
  wire f_u_wallace_rca12_and_8_4_y0;
  wire f_u_wallace_rca12_fa26_f_u_wallace_rca12_fa25_y4;
  wire f_u_wallace_rca12_fa26_f_u_wallace_rca12_and_9_3_y0;
  wire f_u_wallace_rca12_fa26_y0;
  wire f_u_wallace_rca12_fa26_y1;
  wire f_u_wallace_rca12_fa26_f_u_wallace_rca12_and_8_4_y0;
  wire f_u_wallace_rca12_fa26_y2;
  wire f_u_wallace_rca12_fa26_y3;
  wire f_u_wallace_rca12_fa26_y4;
  wire f_u_wallace_rca12_and_9_4_a_9;
  wire f_u_wallace_rca12_and_9_4_b_4;
  wire f_u_wallace_rca12_and_9_4_y0;
  wire f_u_wallace_rca12_and_8_5_a_8;
  wire f_u_wallace_rca12_and_8_5_b_5;
  wire f_u_wallace_rca12_and_8_5_y0;
  wire f_u_wallace_rca12_fa27_f_u_wallace_rca12_fa26_y4;
  wire f_u_wallace_rca12_fa27_f_u_wallace_rca12_and_9_4_y0;
  wire f_u_wallace_rca12_fa27_y0;
  wire f_u_wallace_rca12_fa27_y1;
  wire f_u_wallace_rca12_fa27_f_u_wallace_rca12_and_8_5_y0;
  wire f_u_wallace_rca12_fa27_y2;
  wire f_u_wallace_rca12_fa27_y3;
  wire f_u_wallace_rca12_fa27_y4;
  wire f_u_wallace_rca12_and_9_5_a_9;
  wire f_u_wallace_rca12_and_9_5_b_5;
  wire f_u_wallace_rca12_and_9_5_y0;
  wire f_u_wallace_rca12_and_8_6_a_8;
  wire f_u_wallace_rca12_and_8_6_b_6;
  wire f_u_wallace_rca12_and_8_6_y0;
  wire f_u_wallace_rca12_fa28_f_u_wallace_rca12_fa27_y4;
  wire f_u_wallace_rca12_fa28_f_u_wallace_rca12_and_9_5_y0;
  wire f_u_wallace_rca12_fa28_y0;
  wire f_u_wallace_rca12_fa28_y1;
  wire f_u_wallace_rca12_fa28_f_u_wallace_rca12_and_8_6_y0;
  wire f_u_wallace_rca12_fa28_y2;
  wire f_u_wallace_rca12_fa28_y3;
  wire f_u_wallace_rca12_fa28_y4;
  wire f_u_wallace_rca12_and_9_6_a_9;
  wire f_u_wallace_rca12_and_9_6_b_6;
  wire f_u_wallace_rca12_and_9_6_y0;
  wire f_u_wallace_rca12_and_8_7_a_8;
  wire f_u_wallace_rca12_and_8_7_b_7;
  wire f_u_wallace_rca12_and_8_7_y0;
  wire f_u_wallace_rca12_fa29_f_u_wallace_rca12_fa28_y4;
  wire f_u_wallace_rca12_fa29_f_u_wallace_rca12_and_9_6_y0;
  wire f_u_wallace_rca12_fa29_y0;
  wire f_u_wallace_rca12_fa29_y1;
  wire f_u_wallace_rca12_fa29_f_u_wallace_rca12_and_8_7_y0;
  wire f_u_wallace_rca12_fa29_y2;
  wire f_u_wallace_rca12_fa29_y3;
  wire f_u_wallace_rca12_fa29_y4;
  wire f_u_wallace_rca12_and_9_7_a_9;
  wire f_u_wallace_rca12_and_9_7_b_7;
  wire f_u_wallace_rca12_and_9_7_y0;
  wire f_u_wallace_rca12_and_8_8_a_8;
  wire f_u_wallace_rca12_and_8_8_b_8;
  wire f_u_wallace_rca12_and_8_8_y0;
  wire f_u_wallace_rca12_fa30_f_u_wallace_rca12_fa29_y4;
  wire f_u_wallace_rca12_fa30_f_u_wallace_rca12_and_9_7_y0;
  wire f_u_wallace_rca12_fa30_y0;
  wire f_u_wallace_rca12_fa30_y1;
  wire f_u_wallace_rca12_fa30_f_u_wallace_rca12_and_8_8_y0;
  wire f_u_wallace_rca12_fa30_y2;
  wire f_u_wallace_rca12_fa30_y3;
  wire f_u_wallace_rca12_fa30_y4;
  wire f_u_wallace_rca12_and_9_8_a_9;
  wire f_u_wallace_rca12_and_9_8_b_8;
  wire f_u_wallace_rca12_and_9_8_y0;
  wire f_u_wallace_rca12_and_8_9_a_8;
  wire f_u_wallace_rca12_and_8_9_b_9;
  wire f_u_wallace_rca12_and_8_9_y0;
  wire f_u_wallace_rca12_fa31_f_u_wallace_rca12_fa30_y4;
  wire f_u_wallace_rca12_fa31_f_u_wallace_rca12_and_9_8_y0;
  wire f_u_wallace_rca12_fa31_y0;
  wire f_u_wallace_rca12_fa31_y1;
  wire f_u_wallace_rca12_fa31_f_u_wallace_rca12_and_8_9_y0;
  wire f_u_wallace_rca12_fa31_y2;
  wire f_u_wallace_rca12_fa31_y3;
  wire f_u_wallace_rca12_fa31_y4;
  wire f_u_wallace_rca12_and_9_9_a_9;
  wire f_u_wallace_rca12_and_9_9_b_9;
  wire f_u_wallace_rca12_and_9_9_y0;
  wire f_u_wallace_rca12_and_8_10_a_8;
  wire f_u_wallace_rca12_and_8_10_b_10;
  wire f_u_wallace_rca12_and_8_10_y0;
  wire f_u_wallace_rca12_fa32_f_u_wallace_rca12_fa31_y4;
  wire f_u_wallace_rca12_fa32_f_u_wallace_rca12_and_9_9_y0;
  wire f_u_wallace_rca12_fa32_y0;
  wire f_u_wallace_rca12_fa32_y1;
  wire f_u_wallace_rca12_fa32_f_u_wallace_rca12_and_8_10_y0;
  wire f_u_wallace_rca12_fa32_y2;
  wire f_u_wallace_rca12_fa32_y3;
  wire f_u_wallace_rca12_fa32_y4;
  wire f_u_wallace_rca12_and_9_10_a_9;
  wire f_u_wallace_rca12_and_9_10_b_10;
  wire f_u_wallace_rca12_and_9_10_y0;
  wire f_u_wallace_rca12_and_8_11_a_8;
  wire f_u_wallace_rca12_and_8_11_b_11;
  wire f_u_wallace_rca12_and_8_11_y0;
  wire f_u_wallace_rca12_fa33_f_u_wallace_rca12_fa32_y4;
  wire f_u_wallace_rca12_fa33_f_u_wallace_rca12_and_9_10_y0;
  wire f_u_wallace_rca12_fa33_y0;
  wire f_u_wallace_rca12_fa33_y1;
  wire f_u_wallace_rca12_fa33_f_u_wallace_rca12_and_8_11_y0;
  wire f_u_wallace_rca12_fa33_y2;
  wire f_u_wallace_rca12_fa33_y3;
  wire f_u_wallace_rca12_fa33_y4;
  wire f_u_wallace_rca12_and_0_4_a_0;
  wire f_u_wallace_rca12_and_0_4_b_4;
  wire f_u_wallace_rca12_and_0_4_y0;
  wire f_u_wallace_rca12_ha2_f_u_wallace_rca12_and_0_4_y0;
  wire f_u_wallace_rca12_ha2_f_u_wallace_rca12_fa1_y2;
  wire f_u_wallace_rca12_ha2_y0;
  wire f_u_wallace_rca12_ha2_y1;
  wire f_u_wallace_rca12_and_1_4_a_1;
  wire f_u_wallace_rca12_and_1_4_b_4;
  wire f_u_wallace_rca12_and_1_4_y0;
  wire f_u_wallace_rca12_and_0_5_a_0;
  wire f_u_wallace_rca12_and_0_5_b_5;
  wire f_u_wallace_rca12_and_0_5_y0;
  wire f_u_wallace_rca12_fa34_f_u_wallace_rca12_ha2_y1;
  wire f_u_wallace_rca12_fa34_f_u_wallace_rca12_and_1_4_y0;
  wire f_u_wallace_rca12_fa34_y0;
  wire f_u_wallace_rca12_fa34_y1;
  wire f_u_wallace_rca12_fa34_f_u_wallace_rca12_and_0_5_y0;
  wire f_u_wallace_rca12_fa34_y2;
  wire f_u_wallace_rca12_fa34_y3;
  wire f_u_wallace_rca12_fa34_y4;
  wire f_u_wallace_rca12_and_2_4_a_2;
  wire f_u_wallace_rca12_and_2_4_b_4;
  wire f_u_wallace_rca12_and_2_4_y0;
  wire f_u_wallace_rca12_and_1_5_a_1;
  wire f_u_wallace_rca12_and_1_5_b_5;
  wire f_u_wallace_rca12_and_1_5_y0;
  wire f_u_wallace_rca12_fa35_f_u_wallace_rca12_fa34_y4;
  wire f_u_wallace_rca12_fa35_f_u_wallace_rca12_and_2_4_y0;
  wire f_u_wallace_rca12_fa35_y0;
  wire f_u_wallace_rca12_fa35_y1;
  wire f_u_wallace_rca12_fa35_f_u_wallace_rca12_and_1_5_y0;
  wire f_u_wallace_rca12_fa35_y2;
  wire f_u_wallace_rca12_fa35_y3;
  wire f_u_wallace_rca12_fa35_y4;
  wire f_u_wallace_rca12_and_3_4_a_3;
  wire f_u_wallace_rca12_and_3_4_b_4;
  wire f_u_wallace_rca12_and_3_4_y0;
  wire f_u_wallace_rca12_and_2_5_a_2;
  wire f_u_wallace_rca12_and_2_5_b_5;
  wire f_u_wallace_rca12_and_2_5_y0;
  wire f_u_wallace_rca12_fa36_f_u_wallace_rca12_fa35_y4;
  wire f_u_wallace_rca12_fa36_f_u_wallace_rca12_and_3_4_y0;
  wire f_u_wallace_rca12_fa36_y0;
  wire f_u_wallace_rca12_fa36_y1;
  wire f_u_wallace_rca12_fa36_f_u_wallace_rca12_and_2_5_y0;
  wire f_u_wallace_rca12_fa36_y2;
  wire f_u_wallace_rca12_fa36_y3;
  wire f_u_wallace_rca12_fa36_y4;
  wire f_u_wallace_rca12_and_4_4_a_4;
  wire f_u_wallace_rca12_and_4_4_b_4;
  wire f_u_wallace_rca12_and_4_4_y0;
  wire f_u_wallace_rca12_and_3_5_a_3;
  wire f_u_wallace_rca12_and_3_5_b_5;
  wire f_u_wallace_rca12_and_3_5_y0;
  wire f_u_wallace_rca12_fa37_f_u_wallace_rca12_fa36_y4;
  wire f_u_wallace_rca12_fa37_f_u_wallace_rca12_and_4_4_y0;
  wire f_u_wallace_rca12_fa37_y0;
  wire f_u_wallace_rca12_fa37_y1;
  wire f_u_wallace_rca12_fa37_f_u_wallace_rca12_and_3_5_y0;
  wire f_u_wallace_rca12_fa37_y2;
  wire f_u_wallace_rca12_fa37_y3;
  wire f_u_wallace_rca12_fa37_y4;
  wire f_u_wallace_rca12_and_5_4_a_5;
  wire f_u_wallace_rca12_and_5_4_b_4;
  wire f_u_wallace_rca12_and_5_4_y0;
  wire f_u_wallace_rca12_and_4_5_a_4;
  wire f_u_wallace_rca12_and_4_5_b_5;
  wire f_u_wallace_rca12_and_4_5_y0;
  wire f_u_wallace_rca12_fa38_f_u_wallace_rca12_fa37_y4;
  wire f_u_wallace_rca12_fa38_f_u_wallace_rca12_and_5_4_y0;
  wire f_u_wallace_rca12_fa38_y0;
  wire f_u_wallace_rca12_fa38_y1;
  wire f_u_wallace_rca12_fa38_f_u_wallace_rca12_and_4_5_y0;
  wire f_u_wallace_rca12_fa38_y2;
  wire f_u_wallace_rca12_fa38_y3;
  wire f_u_wallace_rca12_fa38_y4;
  wire f_u_wallace_rca12_and_6_4_a_6;
  wire f_u_wallace_rca12_and_6_4_b_4;
  wire f_u_wallace_rca12_and_6_4_y0;
  wire f_u_wallace_rca12_and_5_5_a_5;
  wire f_u_wallace_rca12_and_5_5_b_5;
  wire f_u_wallace_rca12_and_5_5_y0;
  wire f_u_wallace_rca12_fa39_f_u_wallace_rca12_fa38_y4;
  wire f_u_wallace_rca12_fa39_f_u_wallace_rca12_and_6_4_y0;
  wire f_u_wallace_rca12_fa39_y0;
  wire f_u_wallace_rca12_fa39_y1;
  wire f_u_wallace_rca12_fa39_f_u_wallace_rca12_and_5_5_y0;
  wire f_u_wallace_rca12_fa39_y2;
  wire f_u_wallace_rca12_fa39_y3;
  wire f_u_wallace_rca12_fa39_y4;
  wire f_u_wallace_rca12_and_7_4_a_7;
  wire f_u_wallace_rca12_and_7_4_b_4;
  wire f_u_wallace_rca12_and_7_4_y0;
  wire f_u_wallace_rca12_and_6_5_a_6;
  wire f_u_wallace_rca12_and_6_5_b_5;
  wire f_u_wallace_rca12_and_6_5_y0;
  wire f_u_wallace_rca12_fa40_f_u_wallace_rca12_fa39_y4;
  wire f_u_wallace_rca12_fa40_f_u_wallace_rca12_and_7_4_y0;
  wire f_u_wallace_rca12_fa40_y0;
  wire f_u_wallace_rca12_fa40_y1;
  wire f_u_wallace_rca12_fa40_f_u_wallace_rca12_and_6_5_y0;
  wire f_u_wallace_rca12_fa40_y2;
  wire f_u_wallace_rca12_fa40_y3;
  wire f_u_wallace_rca12_fa40_y4;
  wire f_u_wallace_rca12_and_7_5_a_7;
  wire f_u_wallace_rca12_and_7_5_b_5;
  wire f_u_wallace_rca12_and_7_5_y0;
  wire f_u_wallace_rca12_and_6_6_a_6;
  wire f_u_wallace_rca12_and_6_6_b_6;
  wire f_u_wallace_rca12_and_6_6_y0;
  wire f_u_wallace_rca12_fa41_f_u_wallace_rca12_fa40_y4;
  wire f_u_wallace_rca12_fa41_f_u_wallace_rca12_and_7_5_y0;
  wire f_u_wallace_rca12_fa41_y0;
  wire f_u_wallace_rca12_fa41_y1;
  wire f_u_wallace_rca12_fa41_f_u_wallace_rca12_and_6_6_y0;
  wire f_u_wallace_rca12_fa41_y2;
  wire f_u_wallace_rca12_fa41_y3;
  wire f_u_wallace_rca12_fa41_y4;
  wire f_u_wallace_rca12_and_7_6_a_7;
  wire f_u_wallace_rca12_and_7_6_b_6;
  wire f_u_wallace_rca12_and_7_6_y0;
  wire f_u_wallace_rca12_and_6_7_a_6;
  wire f_u_wallace_rca12_and_6_7_b_7;
  wire f_u_wallace_rca12_and_6_7_y0;
  wire f_u_wallace_rca12_fa42_f_u_wallace_rca12_fa41_y4;
  wire f_u_wallace_rca12_fa42_f_u_wallace_rca12_and_7_6_y0;
  wire f_u_wallace_rca12_fa42_y0;
  wire f_u_wallace_rca12_fa42_y1;
  wire f_u_wallace_rca12_fa42_f_u_wallace_rca12_and_6_7_y0;
  wire f_u_wallace_rca12_fa42_y2;
  wire f_u_wallace_rca12_fa42_y3;
  wire f_u_wallace_rca12_fa42_y4;
  wire f_u_wallace_rca12_and_7_7_a_7;
  wire f_u_wallace_rca12_and_7_7_b_7;
  wire f_u_wallace_rca12_and_7_7_y0;
  wire f_u_wallace_rca12_and_6_8_a_6;
  wire f_u_wallace_rca12_and_6_8_b_8;
  wire f_u_wallace_rca12_and_6_8_y0;
  wire f_u_wallace_rca12_fa43_f_u_wallace_rca12_fa42_y4;
  wire f_u_wallace_rca12_fa43_f_u_wallace_rca12_and_7_7_y0;
  wire f_u_wallace_rca12_fa43_y0;
  wire f_u_wallace_rca12_fa43_y1;
  wire f_u_wallace_rca12_fa43_f_u_wallace_rca12_and_6_8_y0;
  wire f_u_wallace_rca12_fa43_y2;
  wire f_u_wallace_rca12_fa43_y3;
  wire f_u_wallace_rca12_fa43_y4;
  wire f_u_wallace_rca12_and_7_8_a_7;
  wire f_u_wallace_rca12_and_7_8_b_8;
  wire f_u_wallace_rca12_and_7_8_y0;
  wire f_u_wallace_rca12_and_6_9_a_6;
  wire f_u_wallace_rca12_and_6_9_b_9;
  wire f_u_wallace_rca12_and_6_9_y0;
  wire f_u_wallace_rca12_fa44_f_u_wallace_rca12_fa43_y4;
  wire f_u_wallace_rca12_fa44_f_u_wallace_rca12_and_7_8_y0;
  wire f_u_wallace_rca12_fa44_y0;
  wire f_u_wallace_rca12_fa44_y1;
  wire f_u_wallace_rca12_fa44_f_u_wallace_rca12_and_6_9_y0;
  wire f_u_wallace_rca12_fa44_y2;
  wire f_u_wallace_rca12_fa44_y3;
  wire f_u_wallace_rca12_fa44_y4;
  wire f_u_wallace_rca12_and_7_9_a_7;
  wire f_u_wallace_rca12_and_7_9_b_9;
  wire f_u_wallace_rca12_and_7_9_y0;
  wire f_u_wallace_rca12_and_6_10_a_6;
  wire f_u_wallace_rca12_and_6_10_b_10;
  wire f_u_wallace_rca12_and_6_10_y0;
  wire f_u_wallace_rca12_fa45_f_u_wallace_rca12_fa44_y4;
  wire f_u_wallace_rca12_fa45_f_u_wallace_rca12_and_7_9_y0;
  wire f_u_wallace_rca12_fa45_y0;
  wire f_u_wallace_rca12_fa45_y1;
  wire f_u_wallace_rca12_fa45_f_u_wallace_rca12_and_6_10_y0;
  wire f_u_wallace_rca12_fa45_y2;
  wire f_u_wallace_rca12_fa45_y3;
  wire f_u_wallace_rca12_fa45_y4;
  wire f_u_wallace_rca12_and_7_10_a_7;
  wire f_u_wallace_rca12_and_7_10_b_10;
  wire f_u_wallace_rca12_and_7_10_y0;
  wire f_u_wallace_rca12_and_6_11_a_6;
  wire f_u_wallace_rca12_and_6_11_b_11;
  wire f_u_wallace_rca12_and_6_11_y0;
  wire f_u_wallace_rca12_fa46_f_u_wallace_rca12_fa45_y4;
  wire f_u_wallace_rca12_fa46_f_u_wallace_rca12_and_7_10_y0;
  wire f_u_wallace_rca12_fa46_y0;
  wire f_u_wallace_rca12_fa46_y1;
  wire f_u_wallace_rca12_fa46_f_u_wallace_rca12_and_6_11_y0;
  wire f_u_wallace_rca12_fa46_y2;
  wire f_u_wallace_rca12_fa46_y3;
  wire f_u_wallace_rca12_fa46_y4;
  wire f_u_wallace_rca12_and_7_11_a_7;
  wire f_u_wallace_rca12_and_7_11_b_11;
  wire f_u_wallace_rca12_and_7_11_y0;
  wire f_u_wallace_rca12_fa47_f_u_wallace_rca12_fa46_y4;
  wire f_u_wallace_rca12_fa47_f_u_wallace_rca12_and_7_11_y0;
  wire f_u_wallace_rca12_fa47_y0;
  wire f_u_wallace_rca12_fa47_y1;
  wire f_u_wallace_rca12_fa47_f_u_wallace_rca12_fa15_y2;
  wire f_u_wallace_rca12_fa47_y2;
  wire f_u_wallace_rca12_fa47_y3;
  wire f_u_wallace_rca12_fa47_y4;
  wire f_u_wallace_rca12_ha3_f_u_wallace_rca12_fa2_y2;
  wire f_u_wallace_rca12_ha3_f_u_wallace_rca12_fa19_y2;
  wire f_u_wallace_rca12_ha3_y0;
  wire f_u_wallace_rca12_ha3_y1;
  wire f_u_wallace_rca12_and_0_6_a_0;
  wire f_u_wallace_rca12_and_0_6_b_6;
  wire f_u_wallace_rca12_and_0_6_y0;
  wire f_u_wallace_rca12_fa48_f_u_wallace_rca12_ha3_y1;
  wire f_u_wallace_rca12_fa48_f_u_wallace_rca12_and_0_6_y0;
  wire f_u_wallace_rca12_fa48_y0;
  wire f_u_wallace_rca12_fa48_y1;
  wire f_u_wallace_rca12_fa48_f_u_wallace_rca12_fa3_y2;
  wire f_u_wallace_rca12_fa48_y2;
  wire f_u_wallace_rca12_fa48_y3;
  wire f_u_wallace_rca12_fa48_y4;
  wire f_u_wallace_rca12_and_1_6_a_1;
  wire f_u_wallace_rca12_and_1_6_b_6;
  wire f_u_wallace_rca12_and_1_6_y0;
  wire f_u_wallace_rca12_and_0_7_a_0;
  wire f_u_wallace_rca12_and_0_7_b_7;
  wire f_u_wallace_rca12_and_0_7_y0;
  wire f_u_wallace_rca12_fa49_f_u_wallace_rca12_fa48_y4;
  wire f_u_wallace_rca12_fa49_f_u_wallace_rca12_and_1_6_y0;
  wire f_u_wallace_rca12_fa49_y0;
  wire f_u_wallace_rca12_fa49_y1;
  wire f_u_wallace_rca12_fa49_f_u_wallace_rca12_and_0_7_y0;
  wire f_u_wallace_rca12_fa49_y2;
  wire f_u_wallace_rca12_fa49_y3;
  wire f_u_wallace_rca12_fa49_y4;
  wire f_u_wallace_rca12_and_2_6_a_2;
  wire f_u_wallace_rca12_and_2_6_b_6;
  wire f_u_wallace_rca12_and_2_6_y0;
  wire f_u_wallace_rca12_and_1_7_a_1;
  wire f_u_wallace_rca12_and_1_7_b_7;
  wire f_u_wallace_rca12_and_1_7_y0;
  wire f_u_wallace_rca12_fa50_f_u_wallace_rca12_fa49_y4;
  wire f_u_wallace_rca12_fa50_f_u_wallace_rca12_and_2_6_y0;
  wire f_u_wallace_rca12_fa50_y0;
  wire f_u_wallace_rca12_fa50_y1;
  wire f_u_wallace_rca12_fa50_f_u_wallace_rca12_and_1_7_y0;
  wire f_u_wallace_rca12_fa50_y2;
  wire f_u_wallace_rca12_fa50_y3;
  wire f_u_wallace_rca12_fa50_y4;
  wire f_u_wallace_rca12_and_3_6_a_3;
  wire f_u_wallace_rca12_and_3_6_b_6;
  wire f_u_wallace_rca12_and_3_6_y0;
  wire f_u_wallace_rca12_and_2_7_a_2;
  wire f_u_wallace_rca12_and_2_7_b_7;
  wire f_u_wallace_rca12_and_2_7_y0;
  wire f_u_wallace_rca12_fa51_f_u_wallace_rca12_fa50_y4;
  wire f_u_wallace_rca12_fa51_f_u_wallace_rca12_and_3_6_y0;
  wire f_u_wallace_rca12_fa51_y0;
  wire f_u_wallace_rca12_fa51_y1;
  wire f_u_wallace_rca12_fa51_f_u_wallace_rca12_and_2_7_y0;
  wire f_u_wallace_rca12_fa51_y2;
  wire f_u_wallace_rca12_fa51_y3;
  wire f_u_wallace_rca12_fa51_y4;
  wire f_u_wallace_rca12_and_4_6_a_4;
  wire f_u_wallace_rca12_and_4_6_b_6;
  wire f_u_wallace_rca12_and_4_6_y0;
  wire f_u_wallace_rca12_and_3_7_a_3;
  wire f_u_wallace_rca12_and_3_7_b_7;
  wire f_u_wallace_rca12_and_3_7_y0;
  wire f_u_wallace_rca12_fa52_f_u_wallace_rca12_fa51_y4;
  wire f_u_wallace_rca12_fa52_f_u_wallace_rca12_and_4_6_y0;
  wire f_u_wallace_rca12_fa52_y0;
  wire f_u_wallace_rca12_fa52_y1;
  wire f_u_wallace_rca12_fa52_f_u_wallace_rca12_and_3_7_y0;
  wire f_u_wallace_rca12_fa52_y2;
  wire f_u_wallace_rca12_fa52_y3;
  wire f_u_wallace_rca12_fa52_y4;
  wire f_u_wallace_rca12_and_5_6_a_5;
  wire f_u_wallace_rca12_and_5_6_b_6;
  wire f_u_wallace_rca12_and_5_6_y0;
  wire f_u_wallace_rca12_and_4_7_a_4;
  wire f_u_wallace_rca12_and_4_7_b_7;
  wire f_u_wallace_rca12_and_4_7_y0;
  wire f_u_wallace_rca12_fa53_f_u_wallace_rca12_fa52_y4;
  wire f_u_wallace_rca12_fa53_f_u_wallace_rca12_and_5_6_y0;
  wire f_u_wallace_rca12_fa53_y0;
  wire f_u_wallace_rca12_fa53_y1;
  wire f_u_wallace_rca12_fa53_f_u_wallace_rca12_and_4_7_y0;
  wire f_u_wallace_rca12_fa53_y2;
  wire f_u_wallace_rca12_fa53_y3;
  wire f_u_wallace_rca12_fa53_y4;
  wire f_u_wallace_rca12_and_5_7_a_5;
  wire f_u_wallace_rca12_and_5_7_b_7;
  wire f_u_wallace_rca12_and_5_7_y0;
  wire f_u_wallace_rca12_and_4_8_a_4;
  wire f_u_wallace_rca12_and_4_8_b_8;
  wire f_u_wallace_rca12_and_4_8_y0;
  wire f_u_wallace_rca12_fa54_f_u_wallace_rca12_fa53_y4;
  wire f_u_wallace_rca12_fa54_f_u_wallace_rca12_and_5_7_y0;
  wire f_u_wallace_rca12_fa54_y0;
  wire f_u_wallace_rca12_fa54_y1;
  wire f_u_wallace_rca12_fa54_f_u_wallace_rca12_and_4_8_y0;
  wire f_u_wallace_rca12_fa54_y2;
  wire f_u_wallace_rca12_fa54_y3;
  wire f_u_wallace_rca12_fa54_y4;
  wire f_u_wallace_rca12_and_5_8_a_5;
  wire f_u_wallace_rca12_and_5_8_b_8;
  wire f_u_wallace_rca12_and_5_8_y0;
  wire f_u_wallace_rca12_and_4_9_a_4;
  wire f_u_wallace_rca12_and_4_9_b_9;
  wire f_u_wallace_rca12_and_4_9_y0;
  wire f_u_wallace_rca12_fa55_f_u_wallace_rca12_fa54_y4;
  wire f_u_wallace_rca12_fa55_f_u_wallace_rca12_and_5_8_y0;
  wire f_u_wallace_rca12_fa55_y0;
  wire f_u_wallace_rca12_fa55_y1;
  wire f_u_wallace_rca12_fa55_f_u_wallace_rca12_and_4_9_y0;
  wire f_u_wallace_rca12_fa55_y2;
  wire f_u_wallace_rca12_fa55_y3;
  wire f_u_wallace_rca12_fa55_y4;
  wire f_u_wallace_rca12_and_5_9_a_5;
  wire f_u_wallace_rca12_and_5_9_b_9;
  wire f_u_wallace_rca12_and_5_9_y0;
  wire f_u_wallace_rca12_and_4_10_a_4;
  wire f_u_wallace_rca12_and_4_10_b_10;
  wire f_u_wallace_rca12_and_4_10_y0;
  wire f_u_wallace_rca12_fa56_f_u_wallace_rca12_fa55_y4;
  wire f_u_wallace_rca12_fa56_f_u_wallace_rca12_and_5_9_y0;
  wire f_u_wallace_rca12_fa56_y0;
  wire f_u_wallace_rca12_fa56_y1;
  wire f_u_wallace_rca12_fa56_f_u_wallace_rca12_and_4_10_y0;
  wire f_u_wallace_rca12_fa56_y2;
  wire f_u_wallace_rca12_fa56_y3;
  wire f_u_wallace_rca12_fa56_y4;
  wire f_u_wallace_rca12_and_5_10_a_5;
  wire f_u_wallace_rca12_and_5_10_b_10;
  wire f_u_wallace_rca12_and_5_10_y0;
  wire f_u_wallace_rca12_and_4_11_a_4;
  wire f_u_wallace_rca12_and_4_11_b_11;
  wire f_u_wallace_rca12_and_4_11_y0;
  wire f_u_wallace_rca12_fa57_f_u_wallace_rca12_fa56_y4;
  wire f_u_wallace_rca12_fa57_f_u_wallace_rca12_and_5_10_y0;
  wire f_u_wallace_rca12_fa57_y0;
  wire f_u_wallace_rca12_fa57_y1;
  wire f_u_wallace_rca12_fa57_f_u_wallace_rca12_and_4_11_y0;
  wire f_u_wallace_rca12_fa57_y2;
  wire f_u_wallace_rca12_fa57_y3;
  wire f_u_wallace_rca12_fa57_y4;
  wire f_u_wallace_rca12_and_5_11_a_5;
  wire f_u_wallace_rca12_and_5_11_b_11;
  wire f_u_wallace_rca12_and_5_11_y0;
  wire f_u_wallace_rca12_fa58_f_u_wallace_rca12_fa57_y4;
  wire f_u_wallace_rca12_fa58_f_u_wallace_rca12_and_5_11_y0;
  wire f_u_wallace_rca12_fa58_y0;
  wire f_u_wallace_rca12_fa58_y1;
  wire f_u_wallace_rca12_fa58_f_u_wallace_rca12_fa13_y2;
  wire f_u_wallace_rca12_fa58_y2;
  wire f_u_wallace_rca12_fa58_y3;
  wire f_u_wallace_rca12_fa58_y4;
  wire f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa58_y4;
  wire f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa14_y2;
  wire f_u_wallace_rca12_fa59_y0;
  wire f_u_wallace_rca12_fa59_y1;
  wire f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa31_y2;
  wire f_u_wallace_rca12_fa59_y2;
  wire f_u_wallace_rca12_fa59_y3;
  wire f_u_wallace_rca12_fa59_y4;
  wire f_u_wallace_rca12_ha4_f_u_wallace_rca12_fa20_y2;
  wire f_u_wallace_rca12_ha4_f_u_wallace_rca12_fa35_y2;
  wire f_u_wallace_rca12_ha4_y0;
  wire f_u_wallace_rca12_ha4_y1;
  wire f_u_wallace_rca12_fa60_f_u_wallace_rca12_ha4_y1;
  wire f_u_wallace_rca12_fa60_f_u_wallace_rca12_fa4_y2;
  wire f_u_wallace_rca12_fa60_y0;
  wire f_u_wallace_rca12_fa60_y1;
  wire f_u_wallace_rca12_fa60_f_u_wallace_rca12_fa21_y2;
  wire f_u_wallace_rca12_fa60_y2;
  wire f_u_wallace_rca12_fa60_y3;
  wire f_u_wallace_rca12_fa60_y4;
  wire f_u_wallace_rca12_and_0_8_a_0;
  wire f_u_wallace_rca12_and_0_8_b_8;
  wire f_u_wallace_rca12_and_0_8_y0;
  wire f_u_wallace_rca12_fa61_f_u_wallace_rca12_fa60_y4;
  wire f_u_wallace_rca12_fa61_f_u_wallace_rca12_and_0_8_y0;
  wire f_u_wallace_rca12_fa61_y0;
  wire f_u_wallace_rca12_fa61_y1;
  wire f_u_wallace_rca12_fa61_f_u_wallace_rca12_fa5_y2;
  wire f_u_wallace_rca12_fa61_y2;
  wire f_u_wallace_rca12_fa61_y3;
  wire f_u_wallace_rca12_fa61_y4;
  wire f_u_wallace_rca12_and_1_8_a_1;
  wire f_u_wallace_rca12_and_1_8_b_8;
  wire f_u_wallace_rca12_and_1_8_y0;
  wire f_u_wallace_rca12_and_0_9_a_0;
  wire f_u_wallace_rca12_and_0_9_b_9;
  wire f_u_wallace_rca12_and_0_9_y0;
  wire f_u_wallace_rca12_fa62_f_u_wallace_rca12_fa61_y4;
  wire f_u_wallace_rca12_fa62_f_u_wallace_rca12_and_1_8_y0;
  wire f_u_wallace_rca12_fa62_y0;
  wire f_u_wallace_rca12_fa62_y1;
  wire f_u_wallace_rca12_fa62_f_u_wallace_rca12_and_0_9_y0;
  wire f_u_wallace_rca12_fa62_y2;
  wire f_u_wallace_rca12_fa62_y3;
  wire f_u_wallace_rca12_fa62_y4;
  wire f_u_wallace_rca12_and_2_8_a_2;
  wire f_u_wallace_rca12_and_2_8_b_8;
  wire f_u_wallace_rca12_and_2_8_y0;
  wire f_u_wallace_rca12_and_1_9_a_1;
  wire f_u_wallace_rca12_and_1_9_b_9;
  wire f_u_wallace_rca12_and_1_9_y0;
  wire f_u_wallace_rca12_fa63_f_u_wallace_rca12_fa62_y4;
  wire f_u_wallace_rca12_fa63_f_u_wallace_rca12_and_2_8_y0;
  wire f_u_wallace_rca12_fa63_y0;
  wire f_u_wallace_rca12_fa63_y1;
  wire f_u_wallace_rca12_fa63_f_u_wallace_rca12_and_1_9_y0;
  wire f_u_wallace_rca12_fa63_y2;
  wire f_u_wallace_rca12_fa63_y3;
  wire f_u_wallace_rca12_fa63_y4;
  wire f_u_wallace_rca12_and_3_8_a_3;
  wire f_u_wallace_rca12_and_3_8_b_8;
  wire f_u_wallace_rca12_and_3_8_y0;
  wire f_u_wallace_rca12_and_2_9_a_2;
  wire f_u_wallace_rca12_and_2_9_b_9;
  wire f_u_wallace_rca12_and_2_9_y0;
  wire f_u_wallace_rca12_fa64_f_u_wallace_rca12_fa63_y4;
  wire f_u_wallace_rca12_fa64_f_u_wallace_rca12_and_3_8_y0;
  wire f_u_wallace_rca12_fa64_y0;
  wire f_u_wallace_rca12_fa64_y1;
  wire f_u_wallace_rca12_fa64_f_u_wallace_rca12_and_2_9_y0;
  wire f_u_wallace_rca12_fa64_y2;
  wire f_u_wallace_rca12_fa64_y3;
  wire f_u_wallace_rca12_fa64_y4;
  wire f_u_wallace_rca12_and_3_9_a_3;
  wire f_u_wallace_rca12_and_3_9_b_9;
  wire f_u_wallace_rca12_and_3_9_y0;
  wire f_u_wallace_rca12_and_2_10_a_2;
  wire f_u_wallace_rca12_and_2_10_b_10;
  wire f_u_wallace_rca12_and_2_10_y0;
  wire f_u_wallace_rca12_fa65_f_u_wallace_rca12_fa64_y4;
  wire f_u_wallace_rca12_fa65_f_u_wallace_rca12_and_3_9_y0;
  wire f_u_wallace_rca12_fa65_y0;
  wire f_u_wallace_rca12_fa65_y1;
  wire f_u_wallace_rca12_fa65_f_u_wallace_rca12_and_2_10_y0;
  wire f_u_wallace_rca12_fa65_y2;
  wire f_u_wallace_rca12_fa65_y3;
  wire f_u_wallace_rca12_fa65_y4;
  wire f_u_wallace_rca12_and_3_10_a_3;
  wire f_u_wallace_rca12_and_3_10_b_10;
  wire f_u_wallace_rca12_and_3_10_y0;
  wire f_u_wallace_rca12_and_2_11_a_2;
  wire f_u_wallace_rca12_and_2_11_b_11;
  wire f_u_wallace_rca12_and_2_11_y0;
  wire f_u_wallace_rca12_fa66_f_u_wallace_rca12_fa65_y4;
  wire f_u_wallace_rca12_fa66_f_u_wallace_rca12_and_3_10_y0;
  wire f_u_wallace_rca12_fa66_y0;
  wire f_u_wallace_rca12_fa66_y1;
  wire f_u_wallace_rca12_fa66_f_u_wallace_rca12_and_2_11_y0;
  wire f_u_wallace_rca12_fa66_y2;
  wire f_u_wallace_rca12_fa66_y3;
  wire f_u_wallace_rca12_fa66_y4;
  wire f_u_wallace_rca12_and_3_11_a_3;
  wire f_u_wallace_rca12_and_3_11_b_11;
  wire f_u_wallace_rca12_and_3_11_y0;
  wire f_u_wallace_rca12_fa67_f_u_wallace_rca12_fa66_y4;
  wire f_u_wallace_rca12_fa67_f_u_wallace_rca12_and_3_11_y0;
  wire f_u_wallace_rca12_fa67_y0;
  wire f_u_wallace_rca12_fa67_y1;
  wire f_u_wallace_rca12_fa67_f_u_wallace_rca12_fa11_y2;
  wire f_u_wallace_rca12_fa67_y2;
  wire f_u_wallace_rca12_fa67_y3;
  wire f_u_wallace_rca12_fa67_y4;
  wire f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa67_y4;
  wire f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa12_y2;
  wire f_u_wallace_rca12_fa68_y0;
  wire f_u_wallace_rca12_fa68_y1;
  wire f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa29_y2;
  wire f_u_wallace_rca12_fa68_y2;
  wire f_u_wallace_rca12_fa68_y3;
  wire f_u_wallace_rca12_fa68_y4;
  wire f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa68_y4;
  wire f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa30_y2;
  wire f_u_wallace_rca12_fa69_y0;
  wire f_u_wallace_rca12_fa69_y1;
  wire f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa45_y2;
  wire f_u_wallace_rca12_fa69_y2;
  wire f_u_wallace_rca12_fa69_y3;
  wire f_u_wallace_rca12_fa69_y4;
  wire f_u_wallace_rca12_ha5_f_u_wallace_rca12_fa36_y2;
  wire f_u_wallace_rca12_ha5_f_u_wallace_rca12_fa49_y2;
  wire f_u_wallace_rca12_ha5_y0;
  wire f_u_wallace_rca12_ha5_y1;
  wire f_u_wallace_rca12_fa70_f_u_wallace_rca12_ha5_y1;
  wire f_u_wallace_rca12_fa70_f_u_wallace_rca12_fa22_y2;
  wire f_u_wallace_rca12_fa70_y0;
  wire f_u_wallace_rca12_fa70_y1;
  wire f_u_wallace_rca12_fa70_f_u_wallace_rca12_fa37_y2;
  wire f_u_wallace_rca12_fa70_y2;
  wire f_u_wallace_rca12_fa70_y3;
  wire f_u_wallace_rca12_fa70_y4;
  wire f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa70_y4;
  wire f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa6_y2;
  wire f_u_wallace_rca12_fa71_y0;
  wire f_u_wallace_rca12_fa71_y1;
  wire f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa23_y2;
  wire f_u_wallace_rca12_fa71_y2;
  wire f_u_wallace_rca12_fa71_y3;
  wire f_u_wallace_rca12_fa71_y4;
  wire f_u_wallace_rca12_and_0_10_a_0;
  wire f_u_wallace_rca12_and_0_10_b_10;
  wire f_u_wallace_rca12_and_0_10_y0;
  wire f_u_wallace_rca12_fa72_f_u_wallace_rca12_fa71_y4;
  wire f_u_wallace_rca12_fa72_f_u_wallace_rca12_and_0_10_y0;
  wire f_u_wallace_rca12_fa72_y0;
  wire f_u_wallace_rca12_fa72_y1;
  wire f_u_wallace_rca12_fa72_f_u_wallace_rca12_fa7_y2;
  wire f_u_wallace_rca12_fa72_y2;
  wire f_u_wallace_rca12_fa72_y3;
  wire f_u_wallace_rca12_fa72_y4;
  wire f_u_wallace_rca12_and_1_10_a_1;
  wire f_u_wallace_rca12_and_1_10_b_10;
  wire f_u_wallace_rca12_and_1_10_y0;
  wire f_u_wallace_rca12_and_0_11_a_0;
  wire f_u_wallace_rca12_and_0_11_b_11;
  wire f_u_wallace_rca12_and_0_11_y0;
  wire f_u_wallace_rca12_fa73_f_u_wallace_rca12_fa72_y4;
  wire f_u_wallace_rca12_fa73_f_u_wallace_rca12_and_1_10_y0;
  wire f_u_wallace_rca12_fa73_y0;
  wire f_u_wallace_rca12_fa73_y1;
  wire f_u_wallace_rca12_fa73_f_u_wallace_rca12_and_0_11_y0;
  wire f_u_wallace_rca12_fa73_y2;
  wire f_u_wallace_rca12_fa73_y3;
  wire f_u_wallace_rca12_fa73_y4;
  wire f_u_wallace_rca12_and_1_11_a_1;
  wire f_u_wallace_rca12_and_1_11_b_11;
  wire f_u_wallace_rca12_and_1_11_y0;
  wire f_u_wallace_rca12_fa74_f_u_wallace_rca12_fa73_y4;
  wire f_u_wallace_rca12_fa74_f_u_wallace_rca12_and_1_11_y0;
  wire f_u_wallace_rca12_fa74_y0;
  wire f_u_wallace_rca12_fa74_y1;
  wire f_u_wallace_rca12_fa74_f_u_wallace_rca12_fa9_y2;
  wire f_u_wallace_rca12_fa74_y2;
  wire f_u_wallace_rca12_fa74_y3;
  wire f_u_wallace_rca12_fa74_y4;
  wire f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa74_y4;
  wire f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa10_y2;
  wire f_u_wallace_rca12_fa75_y0;
  wire f_u_wallace_rca12_fa75_y1;
  wire f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa27_y2;
  wire f_u_wallace_rca12_fa75_y2;
  wire f_u_wallace_rca12_fa75_y3;
  wire f_u_wallace_rca12_fa75_y4;
  wire f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa75_y4;
  wire f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa28_y2;
  wire f_u_wallace_rca12_fa76_y0;
  wire f_u_wallace_rca12_fa76_y1;
  wire f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa43_y2;
  wire f_u_wallace_rca12_fa76_y2;
  wire f_u_wallace_rca12_fa76_y3;
  wire f_u_wallace_rca12_fa76_y4;
  wire f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa76_y4;
  wire f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa44_y2;
  wire f_u_wallace_rca12_fa77_y0;
  wire f_u_wallace_rca12_fa77_y1;
  wire f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa57_y2;
  wire f_u_wallace_rca12_fa77_y2;
  wire f_u_wallace_rca12_fa77_y3;
  wire f_u_wallace_rca12_fa77_y4;
  wire f_u_wallace_rca12_ha6_f_u_wallace_rca12_fa50_y2;
  wire f_u_wallace_rca12_ha6_f_u_wallace_rca12_fa61_y2;
  wire f_u_wallace_rca12_ha6_y0;
  wire f_u_wallace_rca12_ha6_y1;
  wire f_u_wallace_rca12_fa78_f_u_wallace_rca12_ha6_y1;
  wire f_u_wallace_rca12_fa78_f_u_wallace_rca12_fa38_y2;
  wire f_u_wallace_rca12_fa78_y0;
  wire f_u_wallace_rca12_fa78_y1;
  wire f_u_wallace_rca12_fa78_f_u_wallace_rca12_fa51_y2;
  wire f_u_wallace_rca12_fa78_y2;
  wire f_u_wallace_rca12_fa78_y3;
  wire f_u_wallace_rca12_fa78_y4;
  wire f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa78_y4;
  wire f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa24_y2;
  wire f_u_wallace_rca12_fa79_y0;
  wire f_u_wallace_rca12_fa79_y1;
  wire f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa39_y2;
  wire f_u_wallace_rca12_fa79_y2;
  wire f_u_wallace_rca12_fa79_y3;
  wire f_u_wallace_rca12_fa79_y4;
  wire f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa79_y4;
  wire f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa8_y2;
  wire f_u_wallace_rca12_fa80_y0;
  wire f_u_wallace_rca12_fa80_y1;
  wire f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa25_y2;
  wire f_u_wallace_rca12_fa80_y2;
  wire f_u_wallace_rca12_fa80_y3;
  wire f_u_wallace_rca12_fa80_y4;
  wire f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa80_y4;
  wire f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa26_y2;
  wire f_u_wallace_rca12_fa81_y0;
  wire f_u_wallace_rca12_fa81_y1;
  wire f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa41_y2;
  wire f_u_wallace_rca12_fa81_y2;
  wire f_u_wallace_rca12_fa81_y3;
  wire f_u_wallace_rca12_fa81_y4;
  wire f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa81_y4;
  wire f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa42_y2;
  wire f_u_wallace_rca12_fa82_y0;
  wire f_u_wallace_rca12_fa82_y1;
  wire f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa55_y2;
  wire f_u_wallace_rca12_fa82_y2;
  wire f_u_wallace_rca12_fa82_y3;
  wire f_u_wallace_rca12_fa82_y4;
  wire f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa82_y4;
  wire f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa56_y2;
  wire f_u_wallace_rca12_fa83_y0;
  wire f_u_wallace_rca12_fa83_y1;
  wire f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa67_y2;
  wire f_u_wallace_rca12_fa83_y2;
  wire f_u_wallace_rca12_fa83_y3;
  wire f_u_wallace_rca12_fa83_y4;
  wire f_u_wallace_rca12_ha7_f_u_wallace_rca12_fa62_y2;
  wire f_u_wallace_rca12_ha7_f_u_wallace_rca12_fa71_y2;
  wire f_u_wallace_rca12_ha7_y0;
  wire f_u_wallace_rca12_ha7_y1;
  wire f_u_wallace_rca12_fa84_f_u_wallace_rca12_ha7_y1;
  wire f_u_wallace_rca12_fa84_f_u_wallace_rca12_fa52_y2;
  wire f_u_wallace_rca12_fa84_y0;
  wire f_u_wallace_rca12_fa84_y1;
  wire f_u_wallace_rca12_fa84_f_u_wallace_rca12_fa63_y2;
  wire f_u_wallace_rca12_fa84_y2;
  wire f_u_wallace_rca12_fa84_y3;
  wire f_u_wallace_rca12_fa84_y4;
  wire f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa84_y4;
  wire f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa40_y2;
  wire f_u_wallace_rca12_fa85_y0;
  wire f_u_wallace_rca12_fa85_y1;
  wire f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa53_y2;
  wire f_u_wallace_rca12_fa85_y2;
  wire f_u_wallace_rca12_fa85_y3;
  wire f_u_wallace_rca12_fa85_y4;
  wire f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa85_y4;
  wire f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa54_y2;
  wire f_u_wallace_rca12_fa86_y0;
  wire f_u_wallace_rca12_fa86_y1;
  wire f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa65_y2;
  wire f_u_wallace_rca12_fa86_y2;
  wire f_u_wallace_rca12_fa86_y3;
  wire f_u_wallace_rca12_fa86_y4;
  wire f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa86_y4;
  wire f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa66_y2;
  wire f_u_wallace_rca12_fa87_y0;
  wire f_u_wallace_rca12_fa87_y1;
  wire f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa75_y2;
  wire f_u_wallace_rca12_fa87_y2;
  wire f_u_wallace_rca12_fa87_y3;
  wire f_u_wallace_rca12_fa87_y4;
  wire f_u_wallace_rca12_ha8_f_u_wallace_rca12_fa72_y2;
  wire f_u_wallace_rca12_ha8_f_u_wallace_rca12_fa79_y2;
  wire f_u_wallace_rca12_ha8_y0;
  wire f_u_wallace_rca12_ha8_y1;
  wire f_u_wallace_rca12_fa88_f_u_wallace_rca12_ha8_y1;
  wire f_u_wallace_rca12_fa88_f_u_wallace_rca12_fa64_y2;
  wire f_u_wallace_rca12_fa88_y0;
  wire f_u_wallace_rca12_fa88_y1;
  wire f_u_wallace_rca12_fa88_f_u_wallace_rca12_fa73_y2;
  wire f_u_wallace_rca12_fa88_y2;
  wire f_u_wallace_rca12_fa88_y3;
  wire f_u_wallace_rca12_fa88_y4;
  wire f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa88_y4;
  wire f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa74_y2;
  wire f_u_wallace_rca12_fa89_y0;
  wire f_u_wallace_rca12_fa89_y1;
  wire f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa81_y2;
  wire f_u_wallace_rca12_fa89_y2;
  wire f_u_wallace_rca12_fa89_y3;
  wire f_u_wallace_rca12_fa89_y4;
  wire f_u_wallace_rca12_ha9_f_u_wallace_rca12_fa80_y2;
  wire f_u_wallace_rca12_ha9_f_u_wallace_rca12_fa85_y2;
  wire f_u_wallace_rca12_ha9_y0;
  wire f_u_wallace_rca12_ha9_y1;
  wire f_u_wallace_rca12_ha10_f_u_wallace_rca12_ha9_y1;
  wire f_u_wallace_rca12_ha10_f_u_wallace_rca12_fa86_y2;
  wire f_u_wallace_rca12_ha10_y0;
  wire f_u_wallace_rca12_ha10_y1;
  wire f_u_wallace_rca12_fa90_f_u_wallace_rca12_ha10_y1;
  wire f_u_wallace_rca12_fa90_f_u_wallace_rca12_fa89_y4;
  wire f_u_wallace_rca12_fa90_y0;
  wire f_u_wallace_rca12_fa90_y1;
  wire f_u_wallace_rca12_fa90_f_u_wallace_rca12_fa82_y2;
  wire f_u_wallace_rca12_fa90_y2;
  wire f_u_wallace_rca12_fa90_y3;
  wire f_u_wallace_rca12_fa90_y4;
  wire f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa90_y4;
  wire f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa87_y4;
  wire f_u_wallace_rca12_fa91_y0;
  wire f_u_wallace_rca12_fa91_y1;
  wire f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa76_y2;
  wire f_u_wallace_rca12_fa91_y2;
  wire f_u_wallace_rca12_fa91_y3;
  wire f_u_wallace_rca12_fa91_y4;
  wire f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa91_y4;
  wire f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa83_y4;
  wire f_u_wallace_rca12_fa92_y0;
  wire f_u_wallace_rca12_fa92_y1;
  wire f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa68_y2;
  wire f_u_wallace_rca12_fa92_y2;
  wire f_u_wallace_rca12_fa92_y3;
  wire f_u_wallace_rca12_fa92_y4;
  wire f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa92_y4;
  wire f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa77_y4;
  wire f_u_wallace_rca12_fa93_y0;
  wire f_u_wallace_rca12_fa93_y1;
  wire f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa58_y2;
  wire f_u_wallace_rca12_fa93_y2;
  wire f_u_wallace_rca12_fa93_y3;
  wire f_u_wallace_rca12_fa93_y4;
  wire f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa93_y4;
  wire f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa69_y4;
  wire f_u_wallace_rca12_fa94_y0;
  wire f_u_wallace_rca12_fa94_y1;
  wire f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa46_y2;
  wire f_u_wallace_rca12_fa94_y2;
  wire f_u_wallace_rca12_fa94_y3;
  wire f_u_wallace_rca12_fa94_y4;
  wire f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa94_y4;
  wire f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa59_y4;
  wire f_u_wallace_rca12_fa95_y0;
  wire f_u_wallace_rca12_fa95_y1;
  wire f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa32_y2;
  wire f_u_wallace_rca12_fa95_y2;
  wire f_u_wallace_rca12_fa95_y3;
  wire f_u_wallace_rca12_fa95_y4;
  wire f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa95_y4;
  wire f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa47_y4;
  wire f_u_wallace_rca12_fa96_y0;
  wire f_u_wallace_rca12_fa96_y1;
  wire f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa16_y2;
  wire f_u_wallace_rca12_fa96_y2;
  wire f_u_wallace_rca12_fa96_y3;
  wire f_u_wallace_rca12_fa96_y4;
  wire f_u_wallace_rca12_and_9_11_a_9;
  wire f_u_wallace_rca12_and_9_11_b_11;
  wire f_u_wallace_rca12_and_9_11_y0;
  wire f_u_wallace_rca12_fa97_f_u_wallace_rca12_fa96_y4;
  wire f_u_wallace_rca12_fa97_f_u_wallace_rca12_fa33_y4;
  wire f_u_wallace_rca12_fa97_y0;
  wire f_u_wallace_rca12_fa97_y1;
  wire f_u_wallace_rca12_fa97_f_u_wallace_rca12_and_9_11_y0;
  wire f_u_wallace_rca12_fa97_y2;
  wire f_u_wallace_rca12_fa97_y3;
  wire f_u_wallace_rca12_fa97_y4;
  wire f_u_wallace_rca12_and_11_10_a_11;
  wire f_u_wallace_rca12_and_11_10_b_10;
  wire f_u_wallace_rca12_and_11_10_y0;
  wire f_u_wallace_rca12_fa98_f_u_wallace_rca12_fa97_y4;
  wire f_u_wallace_rca12_fa98_f_u_wallace_rca12_fa17_y4;
  wire f_u_wallace_rca12_fa98_y0;
  wire f_u_wallace_rca12_fa98_y1;
  wire f_u_wallace_rca12_fa98_f_u_wallace_rca12_and_11_10_y0;
  wire f_u_wallace_rca12_fa98_y2;
  wire f_u_wallace_rca12_fa98_y3;
  wire f_u_wallace_rca12_fa98_y4;
  wire f_u_wallace_rca12_and_0_0_a_0;
  wire f_u_wallace_rca12_and_0_0_b_0;
  wire f_u_wallace_rca12_and_0_0_y0;
  wire f_u_wallace_rca12_and_1_0_a_1;
  wire f_u_wallace_rca12_and_1_0_b_0;
  wire f_u_wallace_rca12_and_1_0_y0;
  wire f_u_wallace_rca12_and_0_2_a_0;
  wire f_u_wallace_rca12_and_0_2_b_2;
  wire f_u_wallace_rca12_and_0_2_y0;
  wire f_u_wallace_rca12_and_10_11_a_10;
  wire f_u_wallace_rca12_and_10_11_b_11;
  wire f_u_wallace_rca12_and_10_11_y0;
  wire f_u_wallace_rca12_and_0_1_a_0;
  wire f_u_wallace_rca12_and_0_1_b_1;
  wire f_u_wallace_rca12_and_0_1_y0;
  wire f_u_wallace_rca12_and_11_11_a_11;
  wire f_u_wallace_rca12_and_11_11_b_11;
  wire f_u_wallace_rca12_and_11_11_y0;
  wire f_u_wallace_rca12_u_rca22_ha_f_u_wallace_rca12_and_1_0_y0;
  wire f_u_wallace_rca12_u_rca22_ha_f_u_wallace_rca12_and_0_1_y0;
  wire f_u_wallace_rca12_u_rca22_ha_y0;
  wire f_u_wallace_rca12_u_rca22_ha_y1;
  wire f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_and_0_2_y0;
  wire f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_ha0_y0;
  wire f_u_wallace_rca12_u_rca22_fa1_y0;
  wire f_u_wallace_rca12_u_rca22_fa1_y1;
  wire f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_u_rca22_ha_y1;
  wire f_u_wallace_rca12_u_rca22_fa1_y2;
  wire f_u_wallace_rca12_u_rca22_fa1_y3;
  wire f_u_wallace_rca12_u_rca22_fa1_y4;
  wire f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_fa0_y2;
  wire f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_ha1_y0;
  wire f_u_wallace_rca12_u_rca22_fa2_y0;
  wire f_u_wallace_rca12_u_rca22_fa2_y1;
  wire f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_u_rca22_fa1_y4;
  wire f_u_wallace_rca12_u_rca22_fa2_y2;
  wire f_u_wallace_rca12_u_rca22_fa2_y3;
  wire f_u_wallace_rca12_u_rca22_fa2_y4;
  wire f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_fa18_y2;
  wire f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_ha2_y0;
  wire f_u_wallace_rca12_u_rca22_fa3_y0;
  wire f_u_wallace_rca12_u_rca22_fa3_y1;
  wire f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_u_rca22_fa2_y4;
  wire f_u_wallace_rca12_u_rca22_fa3_y2;
  wire f_u_wallace_rca12_u_rca22_fa3_y3;
  wire f_u_wallace_rca12_u_rca22_fa3_y4;
  wire f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_fa34_y2;
  wire f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_ha3_y0;
  wire f_u_wallace_rca12_u_rca22_fa4_y0;
  wire f_u_wallace_rca12_u_rca22_fa4_y1;
  wire f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_u_rca22_fa3_y4;
  wire f_u_wallace_rca12_u_rca22_fa4_y2;
  wire f_u_wallace_rca12_u_rca22_fa4_y3;
  wire f_u_wallace_rca12_u_rca22_fa4_y4;
  wire f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_fa48_y2;
  wire f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_ha4_y0;
  wire f_u_wallace_rca12_u_rca22_fa5_y0;
  wire f_u_wallace_rca12_u_rca22_fa5_y1;
  wire f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_u_rca22_fa4_y4;
  wire f_u_wallace_rca12_u_rca22_fa5_y2;
  wire f_u_wallace_rca12_u_rca22_fa5_y3;
  wire f_u_wallace_rca12_u_rca22_fa5_y4;
  wire f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_fa60_y2;
  wire f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_ha5_y0;
  wire f_u_wallace_rca12_u_rca22_fa6_y0;
  wire f_u_wallace_rca12_u_rca22_fa6_y1;
  wire f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_u_rca22_fa5_y4;
  wire f_u_wallace_rca12_u_rca22_fa6_y2;
  wire f_u_wallace_rca12_u_rca22_fa6_y3;
  wire f_u_wallace_rca12_u_rca22_fa6_y4;
  wire f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_fa70_y2;
  wire f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_ha6_y0;
  wire f_u_wallace_rca12_u_rca22_fa7_y0;
  wire f_u_wallace_rca12_u_rca22_fa7_y1;
  wire f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_u_rca22_fa6_y4;
  wire f_u_wallace_rca12_u_rca22_fa7_y2;
  wire f_u_wallace_rca12_u_rca22_fa7_y3;
  wire f_u_wallace_rca12_u_rca22_fa7_y4;
  wire f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_fa78_y2;
  wire f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_ha7_y0;
  wire f_u_wallace_rca12_u_rca22_fa8_y0;
  wire f_u_wallace_rca12_u_rca22_fa8_y1;
  wire f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_u_rca22_fa7_y4;
  wire f_u_wallace_rca12_u_rca22_fa8_y2;
  wire f_u_wallace_rca12_u_rca22_fa8_y3;
  wire f_u_wallace_rca12_u_rca22_fa8_y4;
  wire f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_fa84_y2;
  wire f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_ha8_y0;
  wire f_u_wallace_rca12_u_rca22_fa9_y0;
  wire f_u_wallace_rca12_u_rca22_fa9_y1;
  wire f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_u_rca22_fa8_y4;
  wire f_u_wallace_rca12_u_rca22_fa9_y2;
  wire f_u_wallace_rca12_u_rca22_fa9_y3;
  wire f_u_wallace_rca12_u_rca22_fa9_y4;
  wire f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_fa88_y2;
  wire f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_ha9_y0;
  wire f_u_wallace_rca12_u_rca22_fa10_y0;
  wire f_u_wallace_rca12_u_rca22_fa10_y1;
  wire f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_u_rca22_fa9_y4;
  wire f_u_wallace_rca12_u_rca22_fa10_y2;
  wire f_u_wallace_rca12_u_rca22_fa10_y3;
  wire f_u_wallace_rca12_u_rca22_fa10_y4;
  wire f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_fa89_y2;
  wire f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_ha10_y0;
  wire f_u_wallace_rca12_u_rca22_fa11_y0;
  wire f_u_wallace_rca12_u_rca22_fa11_y1;
  wire f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_u_rca22_fa10_y4;
  wire f_u_wallace_rca12_u_rca22_fa11_y2;
  wire f_u_wallace_rca12_u_rca22_fa11_y3;
  wire f_u_wallace_rca12_u_rca22_fa11_y4;
  wire f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_fa87_y2;
  wire f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_fa90_y2;
  wire f_u_wallace_rca12_u_rca22_fa12_y0;
  wire f_u_wallace_rca12_u_rca22_fa12_y1;
  wire f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_u_rca22_fa11_y4;
  wire f_u_wallace_rca12_u_rca22_fa12_y2;
  wire f_u_wallace_rca12_u_rca22_fa12_y3;
  wire f_u_wallace_rca12_u_rca22_fa12_y4;
  wire f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_fa83_y2;
  wire f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_fa91_y2;
  wire f_u_wallace_rca12_u_rca22_fa13_y0;
  wire f_u_wallace_rca12_u_rca22_fa13_y1;
  wire f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_u_rca22_fa12_y4;
  wire f_u_wallace_rca12_u_rca22_fa13_y2;
  wire f_u_wallace_rca12_u_rca22_fa13_y3;
  wire f_u_wallace_rca12_u_rca22_fa13_y4;
  wire f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_fa77_y2;
  wire f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_fa92_y2;
  wire f_u_wallace_rca12_u_rca22_fa14_y0;
  wire f_u_wallace_rca12_u_rca22_fa14_y1;
  wire f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_u_rca22_fa13_y4;
  wire f_u_wallace_rca12_u_rca22_fa14_y2;
  wire f_u_wallace_rca12_u_rca22_fa14_y3;
  wire f_u_wallace_rca12_u_rca22_fa14_y4;
  wire f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_fa69_y2;
  wire f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_fa93_y2;
  wire f_u_wallace_rca12_u_rca22_fa15_y0;
  wire f_u_wallace_rca12_u_rca22_fa15_y1;
  wire f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_u_rca22_fa14_y4;
  wire f_u_wallace_rca12_u_rca22_fa15_y2;
  wire f_u_wallace_rca12_u_rca22_fa15_y3;
  wire f_u_wallace_rca12_u_rca22_fa15_y4;
  wire f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_fa59_y2;
  wire f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_fa94_y2;
  wire f_u_wallace_rca12_u_rca22_fa16_y0;
  wire f_u_wallace_rca12_u_rca22_fa16_y1;
  wire f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_u_rca22_fa15_y4;
  wire f_u_wallace_rca12_u_rca22_fa16_y2;
  wire f_u_wallace_rca12_u_rca22_fa16_y3;
  wire f_u_wallace_rca12_u_rca22_fa16_y4;
  wire f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_fa47_y2;
  wire f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_fa95_y2;
  wire f_u_wallace_rca12_u_rca22_fa17_y0;
  wire f_u_wallace_rca12_u_rca22_fa17_y1;
  wire f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_u_rca22_fa16_y4;
  wire f_u_wallace_rca12_u_rca22_fa17_y2;
  wire f_u_wallace_rca12_u_rca22_fa17_y3;
  wire f_u_wallace_rca12_u_rca22_fa17_y4;
  wire f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_fa33_y2;
  wire f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_fa96_y2;
  wire f_u_wallace_rca12_u_rca22_fa18_y0;
  wire f_u_wallace_rca12_u_rca22_fa18_y1;
  wire f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_u_rca22_fa17_y4;
  wire f_u_wallace_rca12_u_rca22_fa18_y2;
  wire f_u_wallace_rca12_u_rca22_fa18_y3;
  wire f_u_wallace_rca12_u_rca22_fa18_y4;
  wire f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_fa17_y2;
  wire f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_fa97_y2;
  wire f_u_wallace_rca12_u_rca22_fa19_y0;
  wire f_u_wallace_rca12_u_rca22_fa19_y1;
  wire f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_u_rca22_fa18_y4;
  wire f_u_wallace_rca12_u_rca22_fa19_y2;
  wire f_u_wallace_rca12_u_rca22_fa19_y3;
  wire f_u_wallace_rca12_u_rca22_fa19_y4;
  wire f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_and_10_11_y0;
  wire f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_fa98_y2;
  wire f_u_wallace_rca12_u_rca22_fa20_y0;
  wire f_u_wallace_rca12_u_rca22_fa20_y1;
  wire f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_u_rca22_fa19_y4;
  wire f_u_wallace_rca12_u_rca22_fa20_y2;
  wire f_u_wallace_rca12_u_rca22_fa20_y3;
  wire f_u_wallace_rca12_u_rca22_fa20_y4;
  wire f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_fa98_y4;
  wire f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_and_11_11_y0;
  wire f_u_wallace_rca12_u_rca22_fa21_y0;
  wire f_u_wallace_rca12_u_rca22_fa21_y1;
  wire f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_u_rca22_fa20_y4;
  wire f_u_wallace_rca12_u_rca22_fa21_y2;
  wire f_u_wallace_rca12_u_rca22_fa21_y3;
  wire f_u_wallace_rca12_u_rca22_fa21_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign f_u_wallace_rca12_and_2_0_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_2_0_y0 = f_u_wallace_rca12_and_2_0_a_2 & f_u_wallace_rca12_and_2_0_b_0;
  assign f_u_wallace_rca12_and_1_1_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_1_1_y0 = f_u_wallace_rca12_and_1_1_a_1 & f_u_wallace_rca12_and_1_1_b_1;
  assign f_u_wallace_rca12_ha0_f_u_wallace_rca12_and_2_0_y0 = f_u_wallace_rca12_and_2_0_y0;
  assign f_u_wallace_rca12_ha0_f_u_wallace_rca12_and_1_1_y0 = f_u_wallace_rca12_and_1_1_y0;
  assign f_u_wallace_rca12_ha0_y0 = f_u_wallace_rca12_ha0_f_u_wallace_rca12_and_2_0_y0 ^ f_u_wallace_rca12_ha0_f_u_wallace_rca12_and_1_1_y0;
  assign f_u_wallace_rca12_ha0_y1 = f_u_wallace_rca12_ha0_f_u_wallace_rca12_and_2_0_y0 & f_u_wallace_rca12_ha0_f_u_wallace_rca12_and_1_1_y0;
  assign f_u_wallace_rca12_and_3_0_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_3_0_y0 = f_u_wallace_rca12_and_3_0_a_3 & f_u_wallace_rca12_and_3_0_b_0;
  assign f_u_wallace_rca12_and_2_1_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_2_1_y0 = f_u_wallace_rca12_and_2_1_a_2 & f_u_wallace_rca12_and_2_1_b_1;
  assign f_u_wallace_rca12_fa0_f_u_wallace_rca12_ha0_y1 = f_u_wallace_rca12_ha0_y1;
  assign f_u_wallace_rca12_fa0_f_u_wallace_rca12_and_3_0_y0 = f_u_wallace_rca12_and_3_0_y0;
  assign f_u_wallace_rca12_fa0_f_u_wallace_rca12_and_2_1_y0 = f_u_wallace_rca12_and_2_1_y0;
  assign f_u_wallace_rca12_fa0_y0 = f_u_wallace_rca12_fa0_f_u_wallace_rca12_ha0_y1 ^ f_u_wallace_rca12_fa0_f_u_wallace_rca12_and_3_0_y0;
  assign f_u_wallace_rca12_fa0_y1 = f_u_wallace_rca12_fa0_f_u_wallace_rca12_ha0_y1 & f_u_wallace_rca12_fa0_f_u_wallace_rca12_and_3_0_y0;
  assign f_u_wallace_rca12_fa0_y2 = f_u_wallace_rca12_fa0_y0 ^ f_u_wallace_rca12_fa0_f_u_wallace_rca12_and_2_1_y0;
  assign f_u_wallace_rca12_fa0_y3 = f_u_wallace_rca12_fa0_y0 & f_u_wallace_rca12_fa0_f_u_wallace_rca12_and_2_1_y0;
  assign f_u_wallace_rca12_fa0_y4 = f_u_wallace_rca12_fa0_y1 | f_u_wallace_rca12_fa0_y3;
  assign f_u_wallace_rca12_and_4_0_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_4_0_y0 = f_u_wallace_rca12_and_4_0_a_4 & f_u_wallace_rca12_and_4_0_b_0;
  assign f_u_wallace_rca12_and_3_1_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_3_1_y0 = f_u_wallace_rca12_and_3_1_a_3 & f_u_wallace_rca12_and_3_1_b_1;
  assign f_u_wallace_rca12_fa1_f_u_wallace_rca12_fa0_y4 = f_u_wallace_rca12_fa0_y4;
  assign f_u_wallace_rca12_fa1_f_u_wallace_rca12_and_4_0_y0 = f_u_wallace_rca12_and_4_0_y0;
  assign f_u_wallace_rca12_fa1_f_u_wallace_rca12_and_3_1_y0 = f_u_wallace_rca12_and_3_1_y0;
  assign f_u_wallace_rca12_fa1_y0 = f_u_wallace_rca12_fa1_f_u_wallace_rca12_fa0_y4 ^ f_u_wallace_rca12_fa1_f_u_wallace_rca12_and_4_0_y0;
  assign f_u_wallace_rca12_fa1_y1 = f_u_wallace_rca12_fa1_f_u_wallace_rca12_fa0_y4 & f_u_wallace_rca12_fa1_f_u_wallace_rca12_and_4_0_y0;
  assign f_u_wallace_rca12_fa1_y2 = f_u_wallace_rca12_fa1_y0 ^ f_u_wallace_rca12_fa1_f_u_wallace_rca12_and_3_1_y0;
  assign f_u_wallace_rca12_fa1_y3 = f_u_wallace_rca12_fa1_y0 & f_u_wallace_rca12_fa1_f_u_wallace_rca12_and_3_1_y0;
  assign f_u_wallace_rca12_fa1_y4 = f_u_wallace_rca12_fa1_y1 | f_u_wallace_rca12_fa1_y3;
  assign f_u_wallace_rca12_and_5_0_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_5_0_y0 = f_u_wallace_rca12_and_5_0_a_5 & f_u_wallace_rca12_and_5_0_b_0;
  assign f_u_wallace_rca12_and_4_1_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_4_1_y0 = f_u_wallace_rca12_and_4_1_a_4 & f_u_wallace_rca12_and_4_1_b_1;
  assign f_u_wallace_rca12_fa2_f_u_wallace_rca12_fa1_y4 = f_u_wallace_rca12_fa1_y4;
  assign f_u_wallace_rca12_fa2_f_u_wallace_rca12_and_5_0_y0 = f_u_wallace_rca12_and_5_0_y0;
  assign f_u_wallace_rca12_fa2_f_u_wallace_rca12_and_4_1_y0 = f_u_wallace_rca12_and_4_1_y0;
  assign f_u_wallace_rca12_fa2_y0 = f_u_wallace_rca12_fa2_f_u_wallace_rca12_fa1_y4 ^ f_u_wallace_rca12_fa2_f_u_wallace_rca12_and_5_0_y0;
  assign f_u_wallace_rca12_fa2_y1 = f_u_wallace_rca12_fa2_f_u_wallace_rca12_fa1_y4 & f_u_wallace_rca12_fa2_f_u_wallace_rca12_and_5_0_y0;
  assign f_u_wallace_rca12_fa2_y2 = f_u_wallace_rca12_fa2_y0 ^ f_u_wallace_rca12_fa2_f_u_wallace_rca12_and_4_1_y0;
  assign f_u_wallace_rca12_fa2_y3 = f_u_wallace_rca12_fa2_y0 & f_u_wallace_rca12_fa2_f_u_wallace_rca12_and_4_1_y0;
  assign f_u_wallace_rca12_fa2_y4 = f_u_wallace_rca12_fa2_y1 | f_u_wallace_rca12_fa2_y3;
  assign f_u_wallace_rca12_and_6_0_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_6_0_y0 = f_u_wallace_rca12_and_6_0_a_6 & f_u_wallace_rca12_and_6_0_b_0;
  assign f_u_wallace_rca12_and_5_1_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_5_1_y0 = f_u_wallace_rca12_and_5_1_a_5 & f_u_wallace_rca12_and_5_1_b_1;
  assign f_u_wallace_rca12_fa3_f_u_wallace_rca12_fa2_y4 = f_u_wallace_rca12_fa2_y4;
  assign f_u_wallace_rca12_fa3_f_u_wallace_rca12_and_6_0_y0 = f_u_wallace_rca12_and_6_0_y0;
  assign f_u_wallace_rca12_fa3_f_u_wallace_rca12_and_5_1_y0 = f_u_wallace_rca12_and_5_1_y0;
  assign f_u_wallace_rca12_fa3_y0 = f_u_wallace_rca12_fa3_f_u_wallace_rca12_fa2_y4 ^ f_u_wallace_rca12_fa3_f_u_wallace_rca12_and_6_0_y0;
  assign f_u_wallace_rca12_fa3_y1 = f_u_wallace_rca12_fa3_f_u_wallace_rca12_fa2_y4 & f_u_wallace_rca12_fa3_f_u_wallace_rca12_and_6_0_y0;
  assign f_u_wallace_rca12_fa3_y2 = f_u_wallace_rca12_fa3_y0 ^ f_u_wallace_rca12_fa3_f_u_wallace_rca12_and_5_1_y0;
  assign f_u_wallace_rca12_fa3_y3 = f_u_wallace_rca12_fa3_y0 & f_u_wallace_rca12_fa3_f_u_wallace_rca12_and_5_1_y0;
  assign f_u_wallace_rca12_fa3_y4 = f_u_wallace_rca12_fa3_y1 | f_u_wallace_rca12_fa3_y3;
  assign f_u_wallace_rca12_and_7_0_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_7_0_y0 = f_u_wallace_rca12_and_7_0_a_7 & f_u_wallace_rca12_and_7_0_b_0;
  assign f_u_wallace_rca12_and_6_1_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_6_1_y0 = f_u_wallace_rca12_and_6_1_a_6 & f_u_wallace_rca12_and_6_1_b_1;
  assign f_u_wallace_rca12_fa4_f_u_wallace_rca12_fa3_y4 = f_u_wallace_rca12_fa3_y4;
  assign f_u_wallace_rca12_fa4_f_u_wallace_rca12_and_7_0_y0 = f_u_wallace_rca12_and_7_0_y0;
  assign f_u_wallace_rca12_fa4_f_u_wallace_rca12_and_6_1_y0 = f_u_wallace_rca12_and_6_1_y0;
  assign f_u_wallace_rca12_fa4_y0 = f_u_wallace_rca12_fa4_f_u_wallace_rca12_fa3_y4 ^ f_u_wallace_rca12_fa4_f_u_wallace_rca12_and_7_0_y0;
  assign f_u_wallace_rca12_fa4_y1 = f_u_wallace_rca12_fa4_f_u_wallace_rca12_fa3_y4 & f_u_wallace_rca12_fa4_f_u_wallace_rca12_and_7_0_y0;
  assign f_u_wallace_rca12_fa4_y2 = f_u_wallace_rca12_fa4_y0 ^ f_u_wallace_rca12_fa4_f_u_wallace_rca12_and_6_1_y0;
  assign f_u_wallace_rca12_fa4_y3 = f_u_wallace_rca12_fa4_y0 & f_u_wallace_rca12_fa4_f_u_wallace_rca12_and_6_1_y0;
  assign f_u_wallace_rca12_fa4_y4 = f_u_wallace_rca12_fa4_y1 | f_u_wallace_rca12_fa4_y3;
  assign f_u_wallace_rca12_and_8_0_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_8_0_y0 = f_u_wallace_rca12_and_8_0_a_8 & f_u_wallace_rca12_and_8_0_b_0;
  assign f_u_wallace_rca12_and_7_1_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_7_1_y0 = f_u_wallace_rca12_and_7_1_a_7 & f_u_wallace_rca12_and_7_1_b_1;
  assign f_u_wallace_rca12_fa5_f_u_wallace_rca12_fa4_y4 = f_u_wallace_rca12_fa4_y4;
  assign f_u_wallace_rca12_fa5_f_u_wallace_rca12_and_8_0_y0 = f_u_wallace_rca12_and_8_0_y0;
  assign f_u_wallace_rca12_fa5_f_u_wallace_rca12_and_7_1_y0 = f_u_wallace_rca12_and_7_1_y0;
  assign f_u_wallace_rca12_fa5_y0 = f_u_wallace_rca12_fa5_f_u_wallace_rca12_fa4_y4 ^ f_u_wallace_rca12_fa5_f_u_wallace_rca12_and_8_0_y0;
  assign f_u_wallace_rca12_fa5_y1 = f_u_wallace_rca12_fa5_f_u_wallace_rca12_fa4_y4 & f_u_wallace_rca12_fa5_f_u_wallace_rca12_and_8_0_y0;
  assign f_u_wallace_rca12_fa5_y2 = f_u_wallace_rca12_fa5_y0 ^ f_u_wallace_rca12_fa5_f_u_wallace_rca12_and_7_1_y0;
  assign f_u_wallace_rca12_fa5_y3 = f_u_wallace_rca12_fa5_y0 & f_u_wallace_rca12_fa5_f_u_wallace_rca12_and_7_1_y0;
  assign f_u_wallace_rca12_fa5_y4 = f_u_wallace_rca12_fa5_y1 | f_u_wallace_rca12_fa5_y3;
  assign f_u_wallace_rca12_and_9_0_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_9_0_y0 = f_u_wallace_rca12_and_9_0_a_9 & f_u_wallace_rca12_and_9_0_b_0;
  assign f_u_wallace_rca12_and_8_1_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_8_1_y0 = f_u_wallace_rca12_and_8_1_a_8 & f_u_wallace_rca12_and_8_1_b_1;
  assign f_u_wallace_rca12_fa6_f_u_wallace_rca12_fa5_y4 = f_u_wallace_rca12_fa5_y4;
  assign f_u_wallace_rca12_fa6_f_u_wallace_rca12_and_9_0_y0 = f_u_wallace_rca12_and_9_0_y0;
  assign f_u_wallace_rca12_fa6_f_u_wallace_rca12_and_8_1_y0 = f_u_wallace_rca12_and_8_1_y0;
  assign f_u_wallace_rca12_fa6_y0 = f_u_wallace_rca12_fa6_f_u_wallace_rca12_fa5_y4 ^ f_u_wallace_rca12_fa6_f_u_wallace_rca12_and_9_0_y0;
  assign f_u_wallace_rca12_fa6_y1 = f_u_wallace_rca12_fa6_f_u_wallace_rca12_fa5_y4 & f_u_wallace_rca12_fa6_f_u_wallace_rca12_and_9_0_y0;
  assign f_u_wallace_rca12_fa6_y2 = f_u_wallace_rca12_fa6_y0 ^ f_u_wallace_rca12_fa6_f_u_wallace_rca12_and_8_1_y0;
  assign f_u_wallace_rca12_fa6_y3 = f_u_wallace_rca12_fa6_y0 & f_u_wallace_rca12_fa6_f_u_wallace_rca12_and_8_1_y0;
  assign f_u_wallace_rca12_fa6_y4 = f_u_wallace_rca12_fa6_y1 | f_u_wallace_rca12_fa6_y3;
  assign f_u_wallace_rca12_and_10_0_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_10_0_y0 = f_u_wallace_rca12_and_10_0_a_10 & f_u_wallace_rca12_and_10_0_b_0;
  assign f_u_wallace_rca12_and_9_1_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_9_1_y0 = f_u_wallace_rca12_and_9_1_a_9 & f_u_wallace_rca12_and_9_1_b_1;
  assign f_u_wallace_rca12_fa7_f_u_wallace_rca12_fa6_y4 = f_u_wallace_rca12_fa6_y4;
  assign f_u_wallace_rca12_fa7_f_u_wallace_rca12_and_10_0_y0 = f_u_wallace_rca12_and_10_0_y0;
  assign f_u_wallace_rca12_fa7_f_u_wallace_rca12_and_9_1_y0 = f_u_wallace_rca12_and_9_1_y0;
  assign f_u_wallace_rca12_fa7_y0 = f_u_wallace_rca12_fa7_f_u_wallace_rca12_fa6_y4 ^ f_u_wallace_rca12_fa7_f_u_wallace_rca12_and_10_0_y0;
  assign f_u_wallace_rca12_fa7_y1 = f_u_wallace_rca12_fa7_f_u_wallace_rca12_fa6_y4 & f_u_wallace_rca12_fa7_f_u_wallace_rca12_and_10_0_y0;
  assign f_u_wallace_rca12_fa7_y2 = f_u_wallace_rca12_fa7_y0 ^ f_u_wallace_rca12_fa7_f_u_wallace_rca12_and_9_1_y0;
  assign f_u_wallace_rca12_fa7_y3 = f_u_wallace_rca12_fa7_y0 & f_u_wallace_rca12_fa7_f_u_wallace_rca12_and_9_1_y0;
  assign f_u_wallace_rca12_fa7_y4 = f_u_wallace_rca12_fa7_y1 | f_u_wallace_rca12_fa7_y3;
  assign f_u_wallace_rca12_and_11_0_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_11_0_y0 = f_u_wallace_rca12_and_11_0_a_11 & f_u_wallace_rca12_and_11_0_b_0;
  assign f_u_wallace_rca12_and_10_1_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_10_1_y0 = f_u_wallace_rca12_and_10_1_a_10 & f_u_wallace_rca12_and_10_1_b_1;
  assign f_u_wallace_rca12_fa8_f_u_wallace_rca12_fa7_y4 = f_u_wallace_rca12_fa7_y4;
  assign f_u_wallace_rca12_fa8_f_u_wallace_rca12_and_11_0_y0 = f_u_wallace_rca12_and_11_0_y0;
  assign f_u_wallace_rca12_fa8_f_u_wallace_rca12_and_10_1_y0 = f_u_wallace_rca12_and_10_1_y0;
  assign f_u_wallace_rca12_fa8_y0 = f_u_wallace_rca12_fa8_f_u_wallace_rca12_fa7_y4 ^ f_u_wallace_rca12_fa8_f_u_wallace_rca12_and_11_0_y0;
  assign f_u_wallace_rca12_fa8_y1 = f_u_wallace_rca12_fa8_f_u_wallace_rca12_fa7_y4 & f_u_wallace_rca12_fa8_f_u_wallace_rca12_and_11_0_y0;
  assign f_u_wallace_rca12_fa8_y2 = f_u_wallace_rca12_fa8_y0 ^ f_u_wallace_rca12_fa8_f_u_wallace_rca12_and_10_1_y0;
  assign f_u_wallace_rca12_fa8_y3 = f_u_wallace_rca12_fa8_y0 & f_u_wallace_rca12_fa8_f_u_wallace_rca12_and_10_1_y0;
  assign f_u_wallace_rca12_fa8_y4 = f_u_wallace_rca12_fa8_y1 | f_u_wallace_rca12_fa8_y3;
  assign f_u_wallace_rca12_and_11_1_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_11_1_y0 = f_u_wallace_rca12_and_11_1_a_11 & f_u_wallace_rca12_and_11_1_b_1;
  assign f_u_wallace_rca12_and_10_2_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_10_2_y0 = f_u_wallace_rca12_and_10_2_a_10 & f_u_wallace_rca12_and_10_2_b_2;
  assign f_u_wallace_rca12_fa9_f_u_wallace_rca12_fa8_y4 = f_u_wallace_rca12_fa8_y4;
  assign f_u_wallace_rca12_fa9_f_u_wallace_rca12_and_11_1_y0 = f_u_wallace_rca12_and_11_1_y0;
  assign f_u_wallace_rca12_fa9_f_u_wallace_rca12_and_10_2_y0 = f_u_wallace_rca12_and_10_2_y0;
  assign f_u_wallace_rca12_fa9_y0 = f_u_wallace_rca12_fa9_f_u_wallace_rca12_fa8_y4 ^ f_u_wallace_rca12_fa9_f_u_wallace_rca12_and_11_1_y0;
  assign f_u_wallace_rca12_fa9_y1 = f_u_wallace_rca12_fa9_f_u_wallace_rca12_fa8_y4 & f_u_wallace_rca12_fa9_f_u_wallace_rca12_and_11_1_y0;
  assign f_u_wallace_rca12_fa9_y2 = f_u_wallace_rca12_fa9_y0 ^ f_u_wallace_rca12_fa9_f_u_wallace_rca12_and_10_2_y0;
  assign f_u_wallace_rca12_fa9_y3 = f_u_wallace_rca12_fa9_y0 & f_u_wallace_rca12_fa9_f_u_wallace_rca12_and_10_2_y0;
  assign f_u_wallace_rca12_fa9_y4 = f_u_wallace_rca12_fa9_y1 | f_u_wallace_rca12_fa9_y3;
  assign f_u_wallace_rca12_and_11_2_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_11_2_y0 = f_u_wallace_rca12_and_11_2_a_11 & f_u_wallace_rca12_and_11_2_b_2;
  assign f_u_wallace_rca12_and_10_3_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_10_3_y0 = f_u_wallace_rca12_and_10_3_a_10 & f_u_wallace_rca12_and_10_3_b_3;
  assign f_u_wallace_rca12_fa10_f_u_wallace_rca12_fa9_y4 = f_u_wallace_rca12_fa9_y4;
  assign f_u_wallace_rca12_fa10_f_u_wallace_rca12_and_11_2_y0 = f_u_wallace_rca12_and_11_2_y0;
  assign f_u_wallace_rca12_fa10_f_u_wallace_rca12_and_10_3_y0 = f_u_wallace_rca12_and_10_3_y0;
  assign f_u_wallace_rca12_fa10_y0 = f_u_wallace_rca12_fa10_f_u_wallace_rca12_fa9_y4 ^ f_u_wallace_rca12_fa10_f_u_wallace_rca12_and_11_2_y0;
  assign f_u_wallace_rca12_fa10_y1 = f_u_wallace_rca12_fa10_f_u_wallace_rca12_fa9_y4 & f_u_wallace_rca12_fa10_f_u_wallace_rca12_and_11_2_y0;
  assign f_u_wallace_rca12_fa10_y2 = f_u_wallace_rca12_fa10_y0 ^ f_u_wallace_rca12_fa10_f_u_wallace_rca12_and_10_3_y0;
  assign f_u_wallace_rca12_fa10_y3 = f_u_wallace_rca12_fa10_y0 & f_u_wallace_rca12_fa10_f_u_wallace_rca12_and_10_3_y0;
  assign f_u_wallace_rca12_fa10_y4 = f_u_wallace_rca12_fa10_y1 | f_u_wallace_rca12_fa10_y3;
  assign f_u_wallace_rca12_and_11_3_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_11_3_y0 = f_u_wallace_rca12_and_11_3_a_11 & f_u_wallace_rca12_and_11_3_b_3;
  assign f_u_wallace_rca12_and_10_4_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_10_4_y0 = f_u_wallace_rca12_and_10_4_a_10 & f_u_wallace_rca12_and_10_4_b_4;
  assign f_u_wallace_rca12_fa11_f_u_wallace_rca12_fa10_y4 = f_u_wallace_rca12_fa10_y4;
  assign f_u_wallace_rca12_fa11_f_u_wallace_rca12_and_11_3_y0 = f_u_wallace_rca12_and_11_3_y0;
  assign f_u_wallace_rca12_fa11_f_u_wallace_rca12_and_10_4_y0 = f_u_wallace_rca12_and_10_4_y0;
  assign f_u_wallace_rca12_fa11_y0 = f_u_wallace_rca12_fa11_f_u_wallace_rca12_fa10_y4 ^ f_u_wallace_rca12_fa11_f_u_wallace_rca12_and_11_3_y0;
  assign f_u_wallace_rca12_fa11_y1 = f_u_wallace_rca12_fa11_f_u_wallace_rca12_fa10_y4 & f_u_wallace_rca12_fa11_f_u_wallace_rca12_and_11_3_y0;
  assign f_u_wallace_rca12_fa11_y2 = f_u_wallace_rca12_fa11_y0 ^ f_u_wallace_rca12_fa11_f_u_wallace_rca12_and_10_4_y0;
  assign f_u_wallace_rca12_fa11_y3 = f_u_wallace_rca12_fa11_y0 & f_u_wallace_rca12_fa11_f_u_wallace_rca12_and_10_4_y0;
  assign f_u_wallace_rca12_fa11_y4 = f_u_wallace_rca12_fa11_y1 | f_u_wallace_rca12_fa11_y3;
  assign f_u_wallace_rca12_and_11_4_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_11_4_y0 = f_u_wallace_rca12_and_11_4_a_11 & f_u_wallace_rca12_and_11_4_b_4;
  assign f_u_wallace_rca12_and_10_5_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_10_5_y0 = f_u_wallace_rca12_and_10_5_a_10 & f_u_wallace_rca12_and_10_5_b_5;
  assign f_u_wallace_rca12_fa12_f_u_wallace_rca12_fa11_y4 = f_u_wallace_rca12_fa11_y4;
  assign f_u_wallace_rca12_fa12_f_u_wallace_rca12_and_11_4_y0 = f_u_wallace_rca12_and_11_4_y0;
  assign f_u_wallace_rca12_fa12_f_u_wallace_rca12_and_10_5_y0 = f_u_wallace_rca12_and_10_5_y0;
  assign f_u_wallace_rca12_fa12_y0 = f_u_wallace_rca12_fa12_f_u_wallace_rca12_fa11_y4 ^ f_u_wallace_rca12_fa12_f_u_wallace_rca12_and_11_4_y0;
  assign f_u_wallace_rca12_fa12_y1 = f_u_wallace_rca12_fa12_f_u_wallace_rca12_fa11_y4 & f_u_wallace_rca12_fa12_f_u_wallace_rca12_and_11_4_y0;
  assign f_u_wallace_rca12_fa12_y2 = f_u_wallace_rca12_fa12_y0 ^ f_u_wallace_rca12_fa12_f_u_wallace_rca12_and_10_5_y0;
  assign f_u_wallace_rca12_fa12_y3 = f_u_wallace_rca12_fa12_y0 & f_u_wallace_rca12_fa12_f_u_wallace_rca12_and_10_5_y0;
  assign f_u_wallace_rca12_fa12_y4 = f_u_wallace_rca12_fa12_y1 | f_u_wallace_rca12_fa12_y3;
  assign f_u_wallace_rca12_and_11_5_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_11_5_y0 = f_u_wallace_rca12_and_11_5_a_11 & f_u_wallace_rca12_and_11_5_b_5;
  assign f_u_wallace_rca12_and_10_6_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_10_6_y0 = f_u_wallace_rca12_and_10_6_a_10 & f_u_wallace_rca12_and_10_6_b_6;
  assign f_u_wallace_rca12_fa13_f_u_wallace_rca12_fa12_y4 = f_u_wallace_rca12_fa12_y4;
  assign f_u_wallace_rca12_fa13_f_u_wallace_rca12_and_11_5_y0 = f_u_wallace_rca12_and_11_5_y0;
  assign f_u_wallace_rca12_fa13_f_u_wallace_rca12_and_10_6_y0 = f_u_wallace_rca12_and_10_6_y0;
  assign f_u_wallace_rca12_fa13_y0 = f_u_wallace_rca12_fa13_f_u_wallace_rca12_fa12_y4 ^ f_u_wallace_rca12_fa13_f_u_wallace_rca12_and_11_5_y0;
  assign f_u_wallace_rca12_fa13_y1 = f_u_wallace_rca12_fa13_f_u_wallace_rca12_fa12_y4 & f_u_wallace_rca12_fa13_f_u_wallace_rca12_and_11_5_y0;
  assign f_u_wallace_rca12_fa13_y2 = f_u_wallace_rca12_fa13_y0 ^ f_u_wallace_rca12_fa13_f_u_wallace_rca12_and_10_6_y0;
  assign f_u_wallace_rca12_fa13_y3 = f_u_wallace_rca12_fa13_y0 & f_u_wallace_rca12_fa13_f_u_wallace_rca12_and_10_6_y0;
  assign f_u_wallace_rca12_fa13_y4 = f_u_wallace_rca12_fa13_y1 | f_u_wallace_rca12_fa13_y3;
  assign f_u_wallace_rca12_and_11_6_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_11_6_y0 = f_u_wallace_rca12_and_11_6_a_11 & f_u_wallace_rca12_and_11_6_b_6;
  assign f_u_wallace_rca12_and_10_7_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_10_7_y0 = f_u_wallace_rca12_and_10_7_a_10 & f_u_wallace_rca12_and_10_7_b_7;
  assign f_u_wallace_rca12_fa14_f_u_wallace_rca12_fa13_y4 = f_u_wallace_rca12_fa13_y4;
  assign f_u_wallace_rca12_fa14_f_u_wallace_rca12_and_11_6_y0 = f_u_wallace_rca12_and_11_6_y0;
  assign f_u_wallace_rca12_fa14_f_u_wallace_rca12_and_10_7_y0 = f_u_wallace_rca12_and_10_7_y0;
  assign f_u_wallace_rca12_fa14_y0 = f_u_wallace_rca12_fa14_f_u_wallace_rca12_fa13_y4 ^ f_u_wallace_rca12_fa14_f_u_wallace_rca12_and_11_6_y0;
  assign f_u_wallace_rca12_fa14_y1 = f_u_wallace_rca12_fa14_f_u_wallace_rca12_fa13_y4 & f_u_wallace_rca12_fa14_f_u_wallace_rca12_and_11_6_y0;
  assign f_u_wallace_rca12_fa14_y2 = f_u_wallace_rca12_fa14_y0 ^ f_u_wallace_rca12_fa14_f_u_wallace_rca12_and_10_7_y0;
  assign f_u_wallace_rca12_fa14_y3 = f_u_wallace_rca12_fa14_y0 & f_u_wallace_rca12_fa14_f_u_wallace_rca12_and_10_7_y0;
  assign f_u_wallace_rca12_fa14_y4 = f_u_wallace_rca12_fa14_y1 | f_u_wallace_rca12_fa14_y3;
  assign f_u_wallace_rca12_and_11_7_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_11_7_y0 = f_u_wallace_rca12_and_11_7_a_11 & f_u_wallace_rca12_and_11_7_b_7;
  assign f_u_wallace_rca12_and_10_8_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_10_8_y0 = f_u_wallace_rca12_and_10_8_a_10 & f_u_wallace_rca12_and_10_8_b_8;
  assign f_u_wallace_rca12_fa15_f_u_wallace_rca12_fa14_y4 = f_u_wallace_rca12_fa14_y4;
  assign f_u_wallace_rca12_fa15_f_u_wallace_rca12_and_11_7_y0 = f_u_wallace_rca12_and_11_7_y0;
  assign f_u_wallace_rca12_fa15_f_u_wallace_rca12_and_10_8_y0 = f_u_wallace_rca12_and_10_8_y0;
  assign f_u_wallace_rca12_fa15_y0 = f_u_wallace_rca12_fa15_f_u_wallace_rca12_fa14_y4 ^ f_u_wallace_rca12_fa15_f_u_wallace_rca12_and_11_7_y0;
  assign f_u_wallace_rca12_fa15_y1 = f_u_wallace_rca12_fa15_f_u_wallace_rca12_fa14_y4 & f_u_wallace_rca12_fa15_f_u_wallace_rca12_and_11_7_y0;
  assign f_u_wallace_rca12_fa15_y2 = f_u_wallace_rca12_fa15_y0 ^ f_u_wallace_rca12_fa15_f_u_wallace_rca12_and_10_8_y0;
  assign f_u_wallace_rca12_fa15_y3 = f_u_wallace_rca12_fa15_y0 & f_u_wallace_rca12_fa15_f_u_wallace_rca12_and_10_8_y0;
  assign f_u_wallace_rca12_fa15_y4 = f_u_wallace_rca12_fa15_y1 | f_u_wallace_rca12_fa15_y3;
  assign f_u_wallace_rca12_and_11_8_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_11_8_y0 = f_u_wallace_rca12_and_11_8_a_11 & f_u_wallace_rca12_and_11_8_b_8;
  assign f_u_wallace_rca12_and_10_9_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_10_9_y0 = f_u_wallace_rca12_and_10_9_a_10 & f_u_wallace_rca12_and_10_9_b_9;
  assign f_u_wallace_rca12_fa16_f_u_wallace_rca12_fa15_y4 = f_u_wallace_rca12_fa15_y4;
  assign f_u_wallace_rca12_fa16_f_u_wallace_rca12_and_11_8_y0 = f_u_wallace_rca12_and_11_8_y0;
  assign f_u_wallace_rca12_fa16_f_u_wallace_rca12_and_10_9_y0 = f_u_wallace_rca12_and_10_9_y0;
  assign f_u_wallace_rca12_fa16_y0 = f_u_wallace_rca12_fa16_f_u_wallace_rca12_fa15_y4 ^ f_u_wallace_rca12_fa16_f_u_wallace_rca12_and_11_8_y0;
  assign f_u_wallace_rca12_fa16_y1 = f_u_wallace_rca12_fa16_f_u_wallace_rca12_fa15_y4 & f_u_wallace_rca12_fa16_f_u_wallace_rca12_and_11_8_y0;
  assign f_u_wallace_rca12_fa16_y2 = f_u_wallace_rca12_fa16_y0 ^ f_u_wallace_rca12_fa16_f_u_wallace_rca12_and_10_9_y0;
  assign f_u_wallace_rca12_fa16_y3 = f_u_wallace_rca12_fa16_y0 & f_u_wallace_rca12_fa16_f_u_wallace_rca12_and_10_9_y0;
  assign f_u_wallace_rca12_fa16_y4 = f_u_wallace_rca12_fa16_y1 | f_u_wallace_rca12_fa16_y3;
  assign f_u_wallace_rca12_and_11_9_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_11_9_y0 = f_u_wallace_rca12_and_11_9_a_11 & f_u_wallace_rca12_and_11_9_b_9;
  assign f_u_wallace_rca12_and_10_10_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_10_10_y0 = f_u_wallace_rca12_and_10_10_a_10 & f_u_wallace_rca12_and_10_10_b_10;
  assign f_u_wallace_rca12_fa17_f_u_wallace_rca12_fa16_y4 = f_u_wallace_rca12_fa16_y4;
  assign f_u_wallace_rca12_fa17_f_u_wallace_rca12_and_11_9_y0 = f_u_wallace_rca12_and_11_9_y0;
  assign f_u_wallace_rca12_fa17_f_u_wallace_rca12_and_10_10_y0 = f_u_wallace_rca12_and_10_10_y0;
  assign f_u_wallace_rca12_fa17_y0 = f_u_wallace_rca12_fa17_f_u_wallace_rca12_fa16_y4 ^ f_u_wallace_rca12_fa17_f_u_wallace_rca12_and_11_9_y0;
  assign f_u_wallace_rca12_fa17_y1 = f_u_wallace_rca12_fa17_f_u_wallace_rca12_fa16_y4 & f_u_wallace_rca12_fa17_f_u_wallace_rca12_and_11_9_y0;
  assign f_u_wallace_rca12_fa17_y2 = f_u_wallace_rca12_fa17_y0 ^ f_u_wallace_rca12_fa17_f_u_wallace_rca12_and_10_10_y0;
  assign f_u_wallace_rca12_fa17_y3 = f_u_wallace_rca12_fa17_y0 & f_u_wallace_rca12_fa17_f_u_wallace_rca12_and_10_10_y0;
  assign f_u_wallace_rca12_fa17_y4 = f_u_wallace_rca12_fa17_y1 | f_u_wallace_rca12_fa17_y3;
  assign f_u_wallace_rca12_and_1_2_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_1_2_y0 = f_u_wallace_rca12_and_1_2_a_1 & f_u_wallace_rca12_and_1_2_b_2;
  assign f_u_wallace_rca12_and_0_3_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_0_3_y0 = f_u_wallace_rca12_and_0_3_a_0 & f_u_wallace_rca12_and_0_3_b_3;
  assign f_u_wallace_rca12_ha1_f_u_wallace_rca12_and_1_2_y0 = f_u_wallace_rca12_and_1_2_y0;
  assign f_u_wallace_rca12_ha1_f_u_wallace_rca12_and_0_3_y0 = f_u_wallace_rca12_and_0_3_y0;
  assign f_u_wallace_rca12_ha1_y0 = f_u_wallace_rca12_ha1_f_u_wallace_rca12_and_1_2_y0 ^ f_u_wallace_rca12_ha1_f_u_wallace_rca12_and_0_3_y0;
  assign f_u_wallace_rca12_ha1_y1 = f_u_wallace_rca12_ha1_f_u_wallace_rca12_and_1_2_y0 & f_u_wallace_rca12_ha1_f_u_wallace_rca12_and_0_3_y0;
  assign f_u_wallace_rca12_and_2_2_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_2_2_y0 = f_u_wallace_rca12_and_2_2_a_2 & f_u_wallace_rca12_and_2_2_b_2;
  assign f_u_wallace_rca12_and_1_3_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_1_3_y0 = f_u_wallace_rca12_and_1_3_a_1 & f_u_wallace_rca12_and_1_3_b_3;
  assign f_u_wallace_rca12_fa18_f_u_wallace_rca12_ha1_y1 = f_u_wallace_rca12_ha1_y1;
  assign f_u_wallace_rca12_fa18_f_u_wallace_rca12_and_2_2_y0 = f_u_wallace_rca12_and_2_2_y0;
  assign f_u_wallace_rca12_fa18_f_u_wallace_rca12_and_1_3_y0 = f_u_wallace_rca12_and_1_3_y0;
  assign f_u_wallace_rca12_fa18_y0 = f_u_wallace_rca12_fa18_f_u_wallace_rca12_ha1_y1 ^ f_u_wallace_rca12_fa18_f_u_wallace_rca12_and_2_2_y0;
  assign f_u_wallace_rca12_fa18_y1 = f_u_wallace_rca12_fa18_f_u_wallace_rca12_ha1_y1 & f_u_wallace_rca12_fa18_f_u_wallace_rca12_and_2_2_y0;
  assign f_u_wallace_rca12_fa18_y2 = f_u_wallace_rca12_fa18_y0 ^ f_u_wallace_rca12_fa18_f_u_wallace_rca12_and_1_3_y0;
  assign f_u_wallace_rca12_fa18_y3 = f_u_wallace_rca12_fa18_y0 & f_u_wallace_rca12_fa18_f_u_wallace_rca12_and_1_3_y0;
  assign f_u_wallace_rca12_fa18_y4 = f_u_wallace_rca12_fa18_y1 | f_u_wallace_rca12_fa18_y3;
  assign f_u_wallace_rca12_and_3_2_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_3_2_y0 = f_u_wallace_rca12_and_3_2_a_3 & f_u_wallace_rca12_and_3_2_b_2;
  assign f_u_wallace_rca12_and_2_3_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_2_3_y0 = f_u_wallace_rca12_and_2_3_a_2 & f_u_wallace_rca12_and_2_3_b_3;
  assign f_u_wallace_rca12_fa19_f_u_wallace_rca12_fa18_y4 = f_u_wallace_rca12_fa18_y4;
  assign f_u_wallace_rca12_fa19_f_u_wallace_rca12_and_3_2_y0 = f_u_wallace_rca12_and_3_2_y0;
  assign f_u_wallace_rca12_fa19_f_u_wallace_rca12_and_2_3_y0 = f_u_wallace_rca12_and_2_3_y0;
  assign f_u_wallace_rca12_fa19_y0 = f_u_wallace_rca12_fa19_f_u_wallace_rca12_fa18_y4 ^ f_u_wallace_rca12_fa19_f_u_wallace_rca12_and_3_2_y0;
  assign f_u_wallace_rca12_fa19_y1 = f_u_wallace_rca12_fa19_f_u_wallace_rca12_fa18_y4 & f_u_wallace_rca12_fa19_f_u_wallace_rca12_and_3_2_y0;
  assign f_u_wallace_rca12_fa19_y2 = f_u_wallace_rca12_fa19_y0 ^ f_u_wallace_rca12_fa19_f_u_wallace_rca12_and_2_3_y0;
  assign f_u_wallace_rca12_fa19_y3 = f_u_wallace_rca12_fa19_y0 & f_u_wallace_rca12_fa19_f_u_wallace_rca12_and_2_3_y0;
  assign f_u_wallace_rca12_fa19_y4 = f_u_wallace_rca12_fa19_y1 | f_u_wallace_rca12_fa19_y3;
  assign f_u_wallace_rca12_and_4_2_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_4_2_y0 = f_u_wallace_rca12_and_4_2_a_4 & f_u_wallace_rca12_and_4_2_b_2;
  assign f_u_wallace_rca12_and_3_3_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_3_3_y0 = f_u_wallace_rca12_and_3_3_a_3 & f_u_wallace_rca12_and_3_3_b_3;
  assign f_u_wallace_rca12_fa20_f_u_wallace_rca12_fa19_y4 = f_u_wallace_rca12_fa19_y4;
  assign f_u_wallace_rca12_fa20_f_u_wallace_rca12_and_4_2_y0 = f_u_wallace_rca12_and_4_2_y0;
  assign f_u_wallace_rca12_fa20_f_u_wallace_rca12_and_3_3_y0 = f_u_wallace_rca12_and_3_3_y0;
  assign f_u_wallace_rca12_fa20_y0 = f_u_wallace_rca12_fa20_f_u_wallace_rca12_fa19_y4 ^ f_u_wallace_rca12_fa20_f_u_wallace_rca12_and_4_2_y0;
  assign f_u_wallace_rca12_fa20_y1 = f_u_wallace_rca12_fa20_f_u_wallace_rca12_fa19_y4 & f_u_wallace_rca12_fa20_f_u_wallace_rca12_and_4_2_y0;
  assign f_u_wallace_rca12_fa20_y2 = f_u_wallace_rca12_fa20_y0 ^ f_u_wallace_rca12_fa20_f_u_wallace_rca12_and_3_3_y0;
  assign f_u_wallace_rca12_fa20_y3 = f_u_wallace_rca12_fa20_y0 & f_u_wallace_rca12_fa20_f_u_wallace_rca12_and_3_3_y0;
  assign f_u_wallace_rca12_fa20_y4 = f_u_wallace_rca12_fa20_y1 | f_u_wallace_rca12_fa20_y3;
  assign f_u_wallace_rca12_and_5_2_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_5_2_y0 = f_u_wallace_rca12_and_5_2_a_5 & f_u_wallace_rca12_and_5_2_b_2;
  assign f_u_wallace_rca12_and_4_3_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_4_3_y0 = f_u_wallace_rca12_and_4_3_a_4 & f_u_wallace_rca12_and_4_3_b_3;
  assign f_u_wallace_rca12_fa21_f_u_wallace_rca12_fa20_y4 = f_u_wallace_rca12_fa20_y4;
  assign f_u_wallace_rca12_fa21_f_u_wallace_rca12_and_5_2_y0 = f_u_wallace_rca12_and_5_2_y0;
  assign f_u_wallace_rca12_fa21_f_u_wallace_rca12_and_4_3_y0 = f_u_wallace_rca12_and_4_3_y0;
  assign f_u_wallace_rca12_fa21_y0 = f_u_wallace_rca12_fa21_f_u_wallace_rca12_fa20_y4 ^ f_u_wallace_rca12_fa21_f_u_wallace_rca12_and_5_2_y0;
  assign f_u_wallace_rca12_fa21_y1 = f_u_wallace_rca12_fa21_f_u_wallace_rca12_fa20_y4 & f_u_wallace_rca12_fa21_f_u_wallace_rca12_and_5_2_y0;
  assign f_u_wallace_rca12_fa21_y2 = f_u_wallace_rca12_fa21_y0 ^ f_u_wallace_rca12_fa21_f_u_wallace_rca12_and_4_3_y0;
  assign f_u_wallace_rca12_fa21_y3 = f_u_wallace_rca12_fa21_y0 & f_u_wallace_rca12_fa21_f_u_wallace_rca12_and_4_3_y0;
  assign f_u_wallace_rca12_fa21_y4 = f_u_wallace_rca12_fa21_y1 | f_u_wallace_rca12_fa21_y3;
  assign f_u_wallace_rca12_and_6_2_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_6_2_y0 = f_u_wallace_rca12_and_6_2_a_6 & f_u_wallace_rca12_and_6_2_b_2;
  assign f_u_wallace_rca12_and_5_3_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_5_3_y0 = f_u_wallace_rca12_and_5_3_a_5 & f_u_wallace_rca12_and_5_3_b_3;
  assign f_u_wallace_rca12_fa22_f_u_wallace_rca12_fa21_y4 = f_u_wallace_rca12_fa21_y4;
  assign f_u_wallace_rca12_fa22_f_u_wallace_rca12_and_6_2_y0 = f_u_wallace_rca12_and_6_2_y0;
  assign f_u_wallace_rca12_fa22_f_u_wallace_rca12_and_5_3_y0 = f_u_wallace_rca12_and_5_3_y0;
  assign f_u_wallace_rca12_fa22_y0 = f_u_wallace_rca12_fa22_f_u_wallace_rca12_fa21_y4 ^ f_u_wallace_rca12_fa22_f_u_wallace_rca12_and_6_2_y0;
  assign f_u_wallace_rca12_fa22_y1 = f_u_wallace_rca12_fa22_f_u_wallace_rca12_fa21_y4 & f_u_wallace_rca12_fa22_f_u_wallace_rca12_and_6_2_y0;
  assign f_u_wallace_rca12_fa22_y2 = f_u_wallace_rca12_fa22_y0 ^ f_u_wallace_rca12_fa22_f_u_wallace_rca12_and_5_3_y0;
  assign f_u_wallace_rca12_fa22_y3 = f_u_wallace_rca12_fa22_y0 & f_u_wallace_rca12_fa22_f_u_wallace_rca12_and_5_3_y0;
  assign f_u_wallace_rca12_fa22_y4 = f_u_wallace_rca12_fa22_y1 | f_u_wallace_rca12_fa22_y3;
  assign f_u_wallace_rca12_and_7_2_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_7_2_y0 = f_u_wallace_rca12_and_7_2_a_7 & f_u_wallace_rca12_and_7_2_b_2;
  assign f_u_wallace_rca12_and_6_3_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_6_3_y0 = f_u_wallace_rca12_and_6_3_a_6 & f_u_wallace_rca12_and_6_3_b_3;
  assign f_u_wallace_rca12_fa23_f_u_wallace_rca12_fa22_y4 = f_u_wallace_rca12_fa22_y4;
  assign f_u_wallace_rca12_fa23_f_u_wallace_rca12_and_7_2_y0 = f_u_wallace_rca12_and_7_2_y0;
  assign f_u_wallace_rca12_fa23_f_u_wallace_rca12_and_6_3_y0 = f_u_wallace_rca12_and_6_3_y0;
  assign f_u_wallace_rca12_fa23_y0 = f_u_wallace_rca12_fa23_f_u_wallace_rca12_fa22_y4 ^ f_u_wallace_rca12_fa23_f_u_wallace_rca12_and_7_2_y0;
  assign f_u_wallace_rca12_fa23_y1 = f_u_wallace_rca12_fa23_f_u_wallace_rca12_fa22_y4 & f_u_wallace_rca12_fa23_f_u_wallace_rca12_and_7_2_y0;
  assign f_u_wallace_rca12_fa23_y2 = f_u_wallace_rca12_fa23_y0 ^ f_u_wallace_rca12_fa23_f_u_wallace_rca12_and_6_3_y0;
  assign f_u_wallace_rca12_fa23_y3 = f_u_wallace_rca12_fa23_y0 & f_u_wallace_rca12_fa23_f_u_wallace_rca12_and_6_3_y0;
  assign f_u_wallace_rca12_fa23_y4 = f_u_wallace_rca12_fa23_y1 | f_u_wallace_rca12_fa23_y3;
  assign f_u_wallace_rca12_and_8_2_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_8_2_y0 = f_u_wallace_rca12_and_8_2_a_8 & f_u_wallace_rca12_and_8_2_b_2;
  assign f_u_wallace_rca12_and_7_3_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_7_3_y0 = f_u_wallace_rca12_and_7_3_a_7 & f_u_wallace_rca12_and_7_3_b_3;
  assign f_u_wallace_rca12_fa24_f_u_wallace_rca12_fa23_y4 = f_u_wallace_rca12_fa23_y4;
  assign f_u_wallace_rca12_fa24_f_u_wallace_rca12_and_8_2_y0 = f_u_wallace_rca12_and_8_2_y0;
  assign f_u_wallace_rca12_fa24_f_u_wallace_rca12_and_7_3_y0 = f_u_wallace_rca12_and_7_3_y0;
  assign f_u_wallace_rca12_fa24_y0 = f_u_wallace_rca12_fa24_f_u_wallace_rca12_fa23_y4 ^ f_u_wallace_rca12_fa24_f_u_wallace_rca12_and_8_2_y0;
  assign f_u_wallace_rca12_fa24_y1 = f_u_wallace_rca12_fa24_f_u_wallace_rca12_fa23_y4 & f_u_wallace_rca12_fa24_f_u_wallace_rca12_and_8_2_y0;
  assign f_u_wallace_rca12_fa24_y2 = f_u_wallace_rca12_fa24_y0 ^ f_u_wallace_rca12_fa24_f_u_wallace_rca12_and_7_3_y0;
  assign f_u_wallace_rca12_fa24_y3 = f_u_wallace_rca12_fa24_y0 & f_u_wallace_rca12_fa24_f_u_wallace_rca12_and_7_3_y0;
  assign f_u_wallace_rca12_fa24_y4 = f_u_wallace_rca12_fa24_y1 | f_u_wallace_rca12_fa24_y3;
  assign f_u_wallace_rca12_and_9_2_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_9_2_y0 = f_u_wallace_rca12_and_9_2_a_9 & f_u_wallace_rca12_and_9_2_b_2;
  assign f_u_wallace_rca12_and_8_3_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_8_3_y0 = f_u_wallace_rca12_and_8_3_a_8 & f_u_wallace_rca12_and_8_3_b_3;
  assign f_u_wallace_rca12_fa25_f_u_wallace_rca12_fa24_y4 = f_u_wallace_rca12_fa24_y4;
  assign f_u_wallace_rca12_fa25_f_u_wallace_rca12_and_9_2_y0 = f_u_wallace_rca12_and_9_2_y0;
  assign f_u_wallace_rca12_fa25_f_u_wallace_rca12_and_8_3_y0 = f_u_wallace_rca12_and_8_3_y0;
  assign f_u_wallace_rca12_fa25_y0 = f_u_wallace_rca12_fa25_f_u_wallace_rca12_fa24_y4 ^ f_u_wallace_rca12_fa25_f_u_wallace_rca12_and_9_2_y0;
  assign f_u_wallace_rca12_fa25_y1 = f_u_wallace_rca12_fa25_f_u_wallace_rca12_fa24_y4 & f_u_wallace_rca12_fa25_f_u_wallace_rca12_and_9_2_y0;
  assign f_u_wallace_rca12_fa25_y2 = f_u_wallace_rca12_fa25_y0 ^ f_u_wallace_rca12_fa25_f_u_wallace_rca12_and_8_3_y0;
  assign f_u_wallace_rca12_fa25_y3 = f_u_wallace_rca12_fa25_y0 & f_u_wallace_rca12_fa25_f_u_wallace_rca12_and_8_3_y0;
  assign f_u_wallace_rca12_fa25_y4 = f_u_wallace_rca12_fa25_y1 | f_u_wallace_rca12_fa25_y3;
  assign f_u_wallace_rca12_and_9_3_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_3_b_3 = b_3;
  assign f_u_wallace_rca12_and_9_3_y0 = f_u_wallace_rca12_and_9_3_a_9 & f_u_wallace_rca12_and_9_3_b_3;
  assign f_u_wallace_rca12_and_8_4_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_8_4_y0 = f_u_wallace_rca12_and_8_4_a_8 & f_u_wallace_rca12_and_8_4_b_4;
  assign f_u_wallace_rca12_fa26_f_u_wallace_rca12_fa25_y4 = f_u_wallace_rca12_fa25_y4;
  assign f_u_wallace_rca12_fa26_f_u_wallace_rca12_and_9_3_y0 = f_u_wallace_rca12_and_9_3_y0;
  assign f_u_wallace_rca12_fa26_f_u_wallace_rca12_and_8_4_y0 = f_u_wallace_rca12_and_8_4_y0;
  assign f_u_wallace_rca12_fa26_y0 = f_u_wallace_rca12_fa26_f_u_wallace_rca12_fa25_y4 ^ f_u_wallace_rca12_fa26_f_u_wallace_rca12_and_9_3_y0;
  assign f_u_wallace_rca12_fa26_y1 = f_u_wallace_rca12_fa26_f_u_wallace_rca12_fa25_y4 & f_u_wallace_rca12_fa26_f_u_wallace_rca12_and_9_3_y0;
  assign f_u_wallace_rca12_fa26_y2 = f_u_wallace_rca12_fa26_y0 ^ f_u_wallace_rca12_fa26_f_u_wallace_rca12_and_8_4_y0;
  assign f_u_wallace_rca12_fa26_y3 = f_u_wallace_rca12_fa26_y0 & f_u_wallace_rca12_fa26_f_u_wallace_rca12_and_8_4_y0;
  assign f_u_wallace_rca12_fa26_y4 = f_u_wallace_rca12_fa26_y1 | f_u_wallace_rca12_fa26_y3;
  assign f_u_wallace_rca12_and_9_4_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_9_4_y0 = f_u_wallace_rca12_and_9_4_a_9 & f_u_wallace_rca12_and_9_4_b_4;
  assign f_u_wallace_rca12_and_8_5_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_8_5_y0 = f_u_wallace_rca12_and_8_5_a_8 & f_u_wallace_rca12_and_8_5_b_5;
  assign f_u_wallace_rca12_fa27_f_u_wallace_rca12_fa26_y4 = f_u_wallace_rca12_fa26_y4;
  assign f_u_wallace_rca12_fa27_f_u_wallace_rca12_and_9_4_y0 = f_u_wallace_rca12_and_9_4_y0;
  assign f_u_wallace_rca12_fa27_f_u_wallace_rca12_and_8_5_y0 = f_u_wallace_rca12_and_8_5_y0;
  assign f_u_wallace_rca12_fa27_y0 = f_u_wallace_rca12_fa27_f_u_wallace_rca12_fa26_y4 ^ f_u_wallace_rca12_fa27_f_u_wallace_rca12_and_9_4_y0;
  assign f_u_wallace_rca12_fa27_y1 = f_u_wallace_rca12_fa27_f_u_wallace_rca12_fa26_y4 & f_u_wallace_rca12_fa27_f_u_wallace_rca12_and_9_4_y0;
  assign f_u_wallace_rca12_fa27_y2 = f_u_wallace_rca12_fa27_y0 ^ f_u_wallace_rca12_fa27_f_u_wallace_rca12_and_8_5_y0;
  assign f_u_wallace_rca12_fa27_y3 = f_u_wallace_rca12_fa27_y0 & f_u_wallace_rca12_fa27_f_u_wallace_rca12_and_8_5_y0;
  assign f_u_wallace_rca12_fa27_y4 = f_u_wallace_rca12_fa27_y1 | f_u_wallace_rca12_fa27_y3;
  assign f_u_wallace_rca12_and_9_5_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_9_5_y0 = f_u_wallace_rca12_and_9_5_a_9 & f_u_wallace_rca12_and_9_5_b_5;
  assign f_u_wallace_rca12_and_8_6_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_8_6_y0 = f_u_wallace_rca12_and_8_6_a_8 & f_u_wallace_rca12_and_8_6_b_6;
  assign f_u_wallace_rca12_fa28_f_u_wallace_rca12_fa27_y4 = f_u_wallace_rca12_fa27_y4;
  assign f_u_wallace_rca12_fa28_f_u_wallace_rca12_and_9_5_y0 = f_u_wallace_rca12_and_9_5_y0;
  assign f_u_wallace_rca12_fa28_f_u_wallace_rca12_and_8_6_y0 = f_u_wallace_rca12_and_8_6_y0;
  assign f_u_wallace_rca12_fa28_y0 = f_u_wallace_rca12_fa28_f_u_wallace_rca12_fa27_y4 ^ f_u_wallace_rca12_fa28_f_u_wallace_rca12_and_9_5_y0;
  assign f_u_wallace_rca12_fa28_y1 = f_u_wallace_rca12_fa28_f_u_wallace_rca12_fa27_y4 & f_u_wallace_rca12_fa28_f_u_wallace_rca12_and_9_5_y0;
  assign f_u_wallace_rca12_fa28_y2 = f_u_wallace_rca12_fa28_y0 ^ f_u_wallace_rca12_fa28_f_u_wallace_rca12_and_8_6_y0;
  assign f_u_wallace_rca12_fa28_y3 = f_u_wallace_rca12_fa28_y0 & f_u_wallace_rca12_fa28_f_u_wallace_rca12_and_8_6_y0;
  assign f_u_wallace_rca12_fa28_y4 = f_u_wallace_rca12_fa28_y1 | f_u_wallace_rca12_fa28_y3;
  assign f_u_wallace_rca12_and_9_6_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_9_6_y0 = f_u_wallace_rca12_and_9_6_a_9 & f_u_wallace_rca12_and_9_6_b_6;
  assign f_u_wallace_rca12_and_8_7_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_8_7_y0 = f_u_wallace_rca12_and_8_7_a_8 & f_u_wallace_rca12_and_8_7_b_7;
  assign f_u_wallace_rca12_fa29_f_u_wallace_rca12_fa28_y4 = f_u_wallace_rca12_fa28_y4;
  assign f_u_wallace_rca12_fa29_f_u_wallace_rca12_and_9_6_y0 = f_u_wallace_rca12_and_9_6_y0;
  assign f_u_wallace_rca12_fa29_f_u_wallace_rca12_and_8_7_y0 = f_u_wallace_rca12_and_8_7_y0;
  assign f_u_wallace_rca12_fa29_y0 = f_u_wallace_rca12_fa29_f_u_wallace_rca12_fa28_y4 ^ f_u_wallace_rca12_fa29_f_u_wallace_rca12_and_9_6_y0;
  assign f_u_wallace_rca12_fa29_y1 = f_u_wallace_rca12_fa29_f_u_wallace_rca12_fa28_y4 & f_u_wallace_rca12_fa29_f_u_wallace_rca12_and_9_6_y0;
  assign f_u_wallace_rca12_fa29_y2 = f_u_wallace_rca12_fa29_y0 ^ f_u_wallace_rca12_fa29_f_u_wallace_rca12_and_8_7_y0;
  assign f_u_wallace_rca12_fa29_y3 = f_u_wallace_rca12_fa29_y0 & f_u_wallace_rca12_fa29_f_u_wallace_rca12_and_8_7_y0;
  assign f_u_wallace_rca12_fa29_y4 = f_u_wallace_rca12_fa29_y1 | f_u_wallace_rca12_fa29_y3;
  assign f_u_wallace_rca12_and_9_7_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_9_7_y0 = f_u_wallace_rca12_and_9_7_a_9 & f_u_wallace_rca12_and_9_7_b_7;
  assign f_u_wallace_rca12_and_8_8_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_8_8_y0 = f_u_wallace_rca12_and_8_8_a_8 & f_u_wallace_rca12_and_8_8_b_8;
  assign f_u_wallace_rca12_fa30_f_u_wallace_rca12_fa29_y4 = f_u_wallace_rca12_fa29_y4;
  assign f_u_wallace_rca12_fa30_f_u_wallace_rca12_and_9_7_y0 = f_u_wallace_rca12_and_9_7_y0;
  assign f_u_wallace_rca12_fa30_f_u_wallace_rca12_and_8_8_y0 = f_u_wallace_rca12_and_8_8_y0;
  assign f_u_wallace_rca12_fa30_y0 = f_u_wallace_rca12_fa30_f_u_wallace_rca12_fa29_y4 ^ f_u_wallace_rca12_fa30_f_u_wallace_rca12_and_9_7_y0;
  assign f_u_wallace_rca12_fa30_y1 = f_u_wallace_rca12_fa30_f_u_wallace_rca12_fa29_y4 & f_u_wallace_rca12_fa30_f_u_wallace_rca12_and_9_7_y0;
  assign f_u_wallace_rca12_fa30_y2 = f_u_wallace_rca12_fa30_y0 ^ f_u_wallace_rca12_fa30_f_u_wallace_rca12_and_8_8_y0;
  assign f_u_wallace_rca12_fa30_y3 = f_u_wallace_rca12_fa30_y0 & f_u_wallace_rca12_fa30_f_u_wallace_rca12_and_8_8_y0;
  assign f_u_wallace_rca12_fa30_y4 = f_u_wallace_rca12_fa30_y1 | f_u_wallace_rca12_fa30_y3;
  assign f_u_wallace_rca12_and_9_8_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_9_8_y0 = f_u_wallace_rca12_and_9_8_a_9 & f_u_wallace_rca12_and_9_8_b_8;
  assign f_u_wallace_rca12_and_8_9_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_8_9_y0 = f_u_wallace_rca12_and_8_9_a_8 & f_u_wallace_rca12_and_8_9_b_9;
  assign f_u_wallace_rca12_fa31_f_u_wallace_rca12_fa30_y4 = f_u_wallace_rca12_fa30_y4;
  assign f_u_wallace_rca12_fa31_f_u_wallace_rca12_and_9_8_y0 = f_u_wallace_rca12_and_9_8_y0;
  assign f_u_wallace_rca12_fa31_f_u_wallace_rca12_and_8_9_y0 = f_u_wallace_rca12_and_8_9_y0;
  assign f_u_wallace_rca12_fa31_y0 = f_u_wallace_rca12_fa31_f_u_wallace_rca12_fa30_y4 ^ f_u_wallace_rca12_fa31_f_u_wallace_rca12_and_9_8_y0;
  assign f_u_wallace_rca12_fa31_y1 = f_u_wallace_rca12_fa31_f_u_wallace_rca12_fa30_y4 & f_u_wallace_rca12_fa31_f_u_wallace_rca12_and_9_8_y0;
  assign f_u_wallace_rca12_fa31_y2 = f_u_wallace_rca12_fa31_y0 ^ f_u_wallace_rca12_fa31_f_u_wallace_rca12_and_8_9_y0;
  assign f_u_wallace_rca12_fa31_y3 = f_u_wallace_rca12_fa31_y0 & f_u_wallace_rca12_fa31_f_u_wallace_rca12_and_8_9_y0;
  assign f_u_wallace_rca12_fa31_y4 = f_u_wallace_rca12_fa31_y1 | f_u_wallace_rca12_fa31_y3;
  assign f_u_wallace_rca12_and_9_9_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_9_9_y0 = f_u_wallace_rca12_and_9_9_a_9 & f_u_wallace_rca12_and_9_9_b_9;
  assign f_u_wallace_rca12_and_8_10_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_8_10_y0 = f_u_wallace_rca12_and_8_10_a_8 & f_u_wallace_rca12_and_8_10_b_10;
  assign f_u_wallace_rca12_fa32_f_u_wallace_rca12_fa31_y4 = f_u_wallace_rca12_fa31_y4;
  assign f_u_wallace_rca12_fa32_f_u_wallace_rca12_and_9_9_y0 = f_u_wallace_rca12_and_9_9_y0;
  assign f_u_wallace_rca12_fa32_f_u_wallace_rca12_and_8_10_y0 = f_u_wallace_rca12_and_8_10_y0;
  assign f_u_wallace_rca12_fa32_y0 = f_u_wallace_rca12_fa32_f_u_wallace_rca12_fa31_y4 ^ f_u_wallace_rca12_fa32_f_u_wallace_rca12_and_9_9_y0;
  assign f_u_wallace_rca12_fa32_y1 = f_u_wallace_rca12_fa32_f_u_wallace_rca12_fa31_y4 & f_u_wallace_rca12_fa32_f_u_wallace_rca12_and_9_9_y0;
  assign f_u_wallace_rca12_fa32_y2 = f_u_wallace_rca12_fa32_y0 ^ f_u_wallace_rca12_fa32_f_u_wallace_rca12_and_8_10_y0;
  assign f_u_wallace_rca12_fa32_y3 = f_u_wallace_rca12_fa32_y0 & f_u_wallace_rca12_fa32_f_u_wallace_rca12_and_8_10_y0;
  assign f_u_wallace_rca12_fa32_y4 = f_u_wallace_rca12_fa32_y1 | f_u_wallace_rca12_fa32_y3;
  assign f_u_wallace_rca12_and_9_10_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_9_10_y0 = f_u_wallace_rca12_and_9_10_a_9 & f_u_wallace_rca12_and_9_10_b_10;
  assign f_u_wallace_rca12_and_8_11_a_8 = a_8;
  assign f_u_wallace_rca12_and_8_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_8_11_y0 = f_u_wallace_rca12_and_8_11_a_8 & f_u_wallace_rca12_and_8_11_b_11;
  assign f_u_wallace_rca12_fa33_f_u_wallace_rca12_fa32_y4 = f_u_wallace_rca12_fa32_y4;
  assign f_u_wallace_rca12_fa33_f_u_wallace_rca12_and_9_10_y0 = f_u_wallace_rca12_and_9_10_y0;
  assign f_u_wallace_rca12_fa33_f_u_wallace_rca12_and_8_11_y0 = f_u_wallace_rca12_and_8_11_y0;
  assign f_u_wallace_rca12_fa33_y0 = f_u_wallace_rca12_fa33_f_u_wallace_rca12_fa32_y4 ^ f_u_wallace_rca12_fa33_f_u_wallace_rca12_and_9_10_y0;
  assign f_u_wallace_rca12_fa33_y1 = f_u_wallace_rca12_fa33_f_u_wallace_rca12_fa32_y4 & f_u_wallace_rca12_fa33_f_u_wallace_rca12_and_9_10_y0;
  assign f_u_wallace_rca12_fa33_y2 = f_u_wallace_rca12_fa33_y0 ^ f_u_wallace_rca12_fa33_f_u_wallace_rca12_and_8_11_y0;
  assign f_u_wallace_rca12_fa33_y3 = f_u_wallace_rca12_fa33_y0 & f_u_wallace_rca12_fa33_f_u_wallace_rca12_and_8_11_y0;
  assign f_u_wallace_rca12_fa33_y4 = f_u_wallace_rca12_fa33_y1 | f_u_wallace_rca12_fa33_y3;
  assign f_u_wallace_rca12_and_0_4_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_0_4_y0 = f_u_wallace_rca12_and_0_4_a_0 & f_u_wallace_rca12_and_0_4_b_4;
  assign f_u_wallace_rca12_ha2_f_u_wallace_rca12_and_0_4_y0 = f_u_wallace_rca12_and_0_4_y0;
  assign f_u_wallace_rca12_ha2_f_u_wallace_rca12_fa1_y2 = f_u_wallace_rca12_fa1_y2;
  assign f_u_wallace_rca12_ha2_y0 = f_u_wallace_rca12_ha2_f_u_wallace_rca12_and_0_4_y0 ^ f_u_wallace_rca12_ha2_f_u_wallace_rca12_fa1_y2;
  assign f_u_wallace_rca12_ha2_y1 = f_u_wallace_rca12_ha2_f_u_wallace_rca12_and_0_4_y0 & f_u_wallace_rca12_ha2_f_u_wallace_rca12_fa1_y2;
  assign f_u_wallace_rca12_and_1_4_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_1_4_y0 = f_u_wallace_rca12_and_1_4_a_1 & f_u_wallace_rca12_and_1_4_b_4;
  assign f_u_wallace_rca12_and_0_5_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_0_5_y0 = f_u_wallace_rca12_and_0_5_a_0 & f_u_wallace_rca12_and_0_5_b_5;
  assign f_u_wallace_rca12_fa34_f_u_wallace_rca12_ha2_y1 = f_u_wallace_rca12_ha2_y1;
  assign f_u_wallace_rca12_fa34_f_u_wallace_rca12_and_1_4_y0 = f_u_wallace_rca12_and_1_4_y0;
  assign f_u_wallace_rca12_fa34_f_u_wallace_rca12_and_0_5_y0 = f_u_wallace_rca12_and_0_5_y0;
  assign f_u_wallace_rca12_fa34_y0 = f_u_wallace_rca12_fa34_f_u_wallace_rca12_ha2_y1 ^ f_u_wallace_rca12_fa34_f_u_wallace_rca12_and_1_4_y0;
  assign f_u_wallace_rca12_fa34_y1 = f_u_wallace_rca12_fa34_f_u_wallace_rca12_ha2_y1 & f_u_wallace_rca12_fa34_f_u_wallace_rca12_and_1_4_y0;
  assign f_u_wallace_rca12_fa34_y2 = f_u_wallace_rca12_fa34_y0 ^ f_u_wallace_rca12_fa34_f_u_wallace_rca12_and_0_5_y0;
  assign f_u_wallace_rca12_fa34_y3 = f_u_wallace_rca12_fa34_y0 & f_u_wallace_rca12_fa34_f_u_wallace_rca12_and_0_5_y0;
  assign f_u_wallace_rca12_fa34_y4 = f_u_wallace_rca12_fa34_y1 | f_u_wallace_rca12_fa34_y3;
  assign f_u_wallace_rca12_and_2_4_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_2_4_y0 = f_u_wallace_rca12_and_2_4_a_2 & f_u_wallace_rca12_and_2_4_b_4;
  assign f_u_wallace_rca12_and_1_5_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_1_5_y0 = f_u_wallace_rca12_and_1_5_a_1 & f_u_wallace_rca12_and_1_5_b_5;
  assign f_u_wallace_rca12_fa35_f_u_wallace_rca12_fa34_y4 = f_u_wallace_rca12_fa34_y4;
  assign f_u_wallace_rca12_fa35_f_u_wallace_rca12_and_2_4_y0 = f_u_wallace_rca12_and_2_4_y0;
  assign f_u_wallace_rca12_fa35_f_u_wallace_rca12_and_1_5_y0 = f_u_wallace_rca12_and_1_5_y0;
  assign f_u_wallace_rca12_fa35_y0 = f_u_wallace_rca12_fa35_f_u_wallace_rca12_fa34_y4 ^ f_u_wallace_rca12_fa35_f_u_wallace_rca12_and_2_4_y0;
  assign f_u_wallace_rca12_fa35_y1 = f_u_wallace_rca12_fa35_f_u_wallace_rca12_fa34_y4 & f_u_wallace_rca12_fa35_f_u_wallace_rca12_and_2_4_y0;
  assign f_u_wallace_rca12_fa35_y2 = f_u_wallace_rca12_fa35_y0 ^ f_u_wallace_rca12_fa35_f_u_wallace_rca12_and_1_5_y0;
  assign f_u_wallace_rca12_fa35_y3 = f_u_wallace_rca12_fa35_y0 & f_u_wallace_rca12_fa35_f_u_wallace_rca12_and_1_5_y0;
  assign f_u_wallace_rca12_fa35_y4 = f_u_wallace_rca12_fa35_y1 | f_u_wallace_rca12_fa35_y3;
  assign f_u_wallace_rca12_and_3_4_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_3_4_y0 = f_u_wallace_rca12_and_3_4_a_3 & f_u_wallace_rca12_and_3_4_b_4;
  assign f_u_wallace_rca12_and_2_5_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_2_5_y0 = f_u_wallace_rca12_and_2_5_a_2 & f_u_wallace_rca12_and_2_5_b_5;
  assign f_u_wallace_rca12_fa36_f_u_wallace_rca12_fa35_y4 = f_u_wallace_rca12_fa35_y4;
  assign f_u_wallace_rca12_fa36_f_u_wallace_rca12_and_3_4_y0 = f_u_wallace_rca12_and_3_4_y0;
  assign f_u_wallace_rca12_fa36_f_u_wallace_rca12_and_2_5_y0 = f_u_wallace_rca12_and_2_5_y0;
  assign f_u_wallace_rca12_fa36_y0 = f_u_wallace_rca12_fa36_f_u_wallace_rca12_fa35_y4 ^ f_u_wallace_rca12_fa36_f_u_wallace_rca12_and_3_4_y0;
  assign f_u_wallace_rca12_fa36_y1 = f_u_wallace_rca12_fa36_f_u_wallace_rca12_fa35_y4 & f_u_wallace_rca12_fa36_f_u_wallace_rca12_and_3_4_y0;
  assign f_u_wallace_rca12_fa36_y2 = f_u_wallace_rca12_fa36_y0 ^ f_u_wallace_rca12_fa36_f_u_wallace_rca12_and_2_5_y0;
  assign f_u_wallace_rca12_fa36_y3 = f_u_wallace_rca12_fa36_y0 & f_u_wallace_rca12_fa36_f_u_wallace_rca12_and_2_5_y0;
  assign f_u_wallace_rca12_fa36_y4 = f_u_wallace_rca12_fa36_y1 | f_u_wallace_rca12_fa36_y3;
  assign f_u_wallace_rca12_and_4_4_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_4_4_y0 = f_u_wallace_rca12_and_4_4_a_4 & f_u_wallace_rca12_and_4_4_b_4;
  assign f_u_wallace_rca12_and_3_5_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_3_5_y0 = f_u_wallace_rca12_and_3_5_a_3 & f_u_wallace_rca12_and_3_5_b_5;
  assign f_u_wallace_rca12_fa37_f_u_wallace_rca12_fa36_y4 = f_u_wallace_rca12_fa36_y4;
  assign f_u_wallace_rca12_fa37_f_u_wallace_rca12_and_4_4_y0 = f_u_wallace_rca12_and_4_4_y0;
  assign f_u_wallace_rca12_fa37_f_u_wallace_rca12_and_3_5_y0 = f_u_wallace_rca12_and_3_5_y0;
  assign f_u_wallace_rca12_fa37_y0 = f_u_wallace_rca12_fa37_f_u_wallace_rca12_fa36_y4 ^ f_u_wallace_rca12_fa37_f_u_wallace_rca12_and_4_4_y0;
  assign f_u_wallace_rca12_fa37_y1 = f_u_wallace_rca12_fa37_f_u_wallace_rca12_fa36_y4 & f_u_wallace_rca12_fa37_f_u_wallace_rca12_and_4_4_y0;
  assign f_u_wallace_rca12_fa37_y2 = f_u_wallace_rca12_fa37_y0 ^ f_u_wallace_rca12_fa37_f_u_wallace_rca12_and_3_5_y0;
  assign f_u_wallace_rca12_fa37_y3 = f_u_wallace_rca12_fa37_y0 & f_u_wallace_rca12_fa37_f_u_wallace_rca12_and_3_5_y0;
  assign f_u_wallace_rca12_fa37_y4 = f_u_wallace_rca12_fa37_y1 | f_u_wallace_rca12_fa37_y3;
  assign f_u_wallace_rca12_and_5_4_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_5_4_y0 = f_u_wallace_rca12_and_5_4_a_5 & f_u_wallace_rca12_and_5_4_b_4;
  assign f_u_wallace_rca12_and_4_5_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_4_5_y0 = f_u_wallace_rca12_and_4_5_a_4 & f_u_wallace_rca12_and_4_5_b_5;
  assign f_u_wallace_rca12_fa38_f_u_wallace_rca12_fa37_y4 = f_u_wallace_rca12_fa37_y4;
  assign f_u_wallace_rca12_fa38_f_u_wallace_rca12_and_5_4_y0 = f_u_wallace_rca12_and_5_4_y0;
  assign f_u_wallace_rca12_fa38_f_u_wallace_rca12_and_4_5_y0 = f_u_wallace_rca12_and_4_5_y0;
  assign f_u_wallace_rca12_fa38_y0 = f_u_wallace_rca12_fa38_f_u_wallace_rca12_fa37_y4 ^ f_u_wallace_rca12_fa38_f_u_wallace_rca12_and_5_4_y0;
  assign f_u_wallace_rca12_fa38_y1 = f_u_wallace_rca12_fa38_f_u_wallace_rca12_fa37_y4 & f_u_wallace_rca12_fa38_f_u_wallace_rca12_and_5_4_y0;
  assign f_u_wallace_rca12_fa38_y2 = f_u_wallace_rca12_fa38_y0 ^ f_u_wallace_rca12_fa38_f_u_wallace_rca12_and_4_5_y0;
  assign f_u_wallace_rca12_fa38_y3 = f_u_wallace_rca12_fa38_y0 & f_u_wallace_rca12_fa38_f_u_wallace_rca12_and_4_5_y0;
  assign f_u_wallace_rca12_fa38_y4 = f_u_wallace_rca12_fa38_y1 | f_u_wallace_rca12_fa38_y3;
  assign f_u_wallace_rca12_and_6_4_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_6_4_y0 = f_u_wallace_rca12_and_6_4_a_6 & f_u_wallace_rca12_and_6_4_b_4;
  assign f_u_wallace_rca12_and_5_5_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_5_5_y0 = f_u_wallace_rca12_and_5_5_a_5 & f_u_wallace_rca12_and_5_5_b_5;
  assign f_u_wallace_rca12_fa39_f_u_wallace_rca12_fa38_y4 = f_u_wallace_rca12_fa38_y4;
  assign f_u_wallace_rca12_fa39_f_u_wallace_rca12_and_6_4_y0 = f_u_wallace_rca12_and_6_4_y0;
  assign f_u_wallace_rca12_fa39_f_u_wallace_rca12_and_5_5_y0 = f_u_wallace_rca12_and_5_5_y0;
  assign f_u_wallace_rca12_fa39_y0 = f_u_wallace_rca12_fa39_f_u_wallace_rca12_fa38_y4 ^ f_u_wallace_rca12_fa39_f_u_wallace_rca12_and_6_4_y0;
  assign f_u_wallace_rca12_fa39_y1 = f_u_wallace_rca12_fa39_f_u_wallace_rca12_fa38_y4 & f_u_wallace_rca12_fa39_f_u_wallace_rca12_and_6_4_y0;
  assign f_u_wallace_rca12_fa39_y2 = f_u_wallace_rca12_fa39_y0 ^ f_u_wallace_rca12_fa39_f_u_wallace_rca12_and_5_5_y0;
  assign f_u_wallace_rca12_fa39_y3 = f_u_wallace_rca12_fa39_y0 & f_u_wallace_rca12_fa39_f_u_wallace_rca12_and_5_5_y0;
  assign f_u_wallace_rca12_fa39_y4 = f_u_wallace_rca12_fa39_y1 | f_u_wallace_rca12_fa39_y3;
  assign f_u_wallace_rca12_and_7_4_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_4_b_4 = b_4;
  assign f_u_wallace_rca12_and_7_4_y0 = f_u_wallace_rca12_and_7_4_a_7 & f_u_wallace_rca12_and_7_4_b_4;
  assign f_u_wallace_rca12_and_6_5_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_6_5_y0 = f_u_wallace_rca12_and_6_5_a_6 & f_u_wallace_rca12_and_6_5_b_5;
  assign f_u_wallace_rca12_fa40_f_u_wallace_rca12_fa39_y4 = f_u_wallace_rca12_fa39_y4;
  assign f_u_wallace_rca12_fa40_f_u_wallace_rca12_and_7_4_y0 = f_u_wallace_rca12_and_7_4_y0;
  assign f_u_wallace_rca12_fa40_f_u_wallace_rca12_and_6_5_y0 = f_u_wallace_rca12_and_6_5_y0;
  assign f_u_wallace_rca12_fa40_y0 = f_u_wallace_rca12_fa40_f_u_wallace_rca12_fa39_y4 ^ f_u_wallace_rca12_fa40_f_u_wallace_rca12_and_7_4_y0;
  assign f_u_wallace_rca12_fa40_y1 = f_u_wallace_rca12_fa40_f_u_wallace_rca12_fa39_y4 & f_u_wallace_rca12_fa40_f_u_wallace_rca12_and_7_4_y0;
  assign f_u_wallace_rca12_fa40_y2 = f_u_wallace_rca12_fa40_y0 ^ f_u_wallace_rca12_fa40_f_u_wallace_rca12_and_6_5_y0;
  assign f_u_wallace_rca12_fa40_y3 = f_u_wallace_rca12_fa40_y0 & f_u_wallace_rca12_fa40_f_u_wallace_rca12_and_6_5_y0;
  assign f_u_wallace_rca12_fa40_y4 = f_u_wallace_rca12_fa40_y1 | f_u_wallace_rca12_fa40_y3;
  assign f_u_wallace_rca12_and_7_5_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_5_b_5 = b_5;
  assign f_u_wallace_rca12_and_7_5_y0 = f_u_wallace_rca12_and_7_5_a_7 & f_u_wallace_rca12_and_7_5_b_5;
  assign f_u_wallace_rca12_and_6_6_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_6_6_y0 = f_u_wallace_rca12_and_6_6_a_6 & f_u_wallace_rca12_and_6_6_b_6;
  assign f_u_wallace_rca12_fa41_f_u_wallace_rca12_fa40_y4 = f_u_wallace_rca12_fa40_y4;
  assign f_u_wallace_rca12_fa41_f_u_wallace_rca12_and_7_5_y0 = f_u_wallace_rca12_and_7_5_y0;
  assign f_u_wallace_rca12_fa41_f_u_wallace_rca12_and_6_6_y0 = f_u_wallace_rca12_and_6_6_y0;
  assign f_u_wallace_rca12_fa41_y0 = f_u_wallace_rca12_fa41_f_u_wallace_rca12_fa40_y4 ^ f_u_wallace_rca12_fa41_f_u_wallace_rca12_and_7_5_y0;
  assign f_u_wallace_rca12_fa41_y1 = f_u_wallace_rca12_fa41_f_u_wallace_rca12_fa40_y4 & f_u_wallace_rca12_fa41_f_u_wallace_rca12_and_7_5_y0;
  assign f_u_wallace_rca12_fa41_y2 = f_u_wallace_rca12_fa41_y0 ^ f_u_wallace_rca12_fa41_f_u_wallace_rca12_and_6_6_y0;
  assign f_u_wallace_rca12_fa41_y3 = f_u_wallace_rca12_fa41_y0 & f_u_wallace_rca12_fa41_f_u_wallace_rca12_and_6_6_y0;
  assign f_u_wallace_rca12_fa41_y4 = f_u_wallace_rca12_fa41_y1 | f_u_wallace_rca12_fa41_y3;
  assign f_u_wallace_rca12_and_7_6_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_7_6_y0 = f_u_wallace_rca12_and_7_6_a_7 & f_u_wallace_rca12_and_7_6_b_6;
  assign f_u_wallace_rca12_and_6_7_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_6_7_y0 = f_u_wallace_rca12_and_6_7_a_6 & f_u_wallace_rca12_and_6_7_b_7;
  assign f_u_wallace_rca12_fa42_f_u_wallace_rca12_fa41_y4 = f_u_wallace_rca12_fa41_y4;
  assign f_u_wallace_rca12_fa42_f_u_wallace_rca12_and_7_6_y0 = f_u_wallace_rca12_and_7_6_y0;
  assign f_u_wallace_rca12_fa42_f_u_wallace_rca12_and_6_7_y0 = f_u_wallace_rca12_and_6_7_y0;
  assign f_u_wallace_rca12_fa42_y0 = f_u_wallace_rca12_fa42_f_u_wallace_rca12_fa41_y4 ^ f_u_wallace_rca12_fa42_f_u_wallace_rca12_and_7_6_y0;
  assign f_u_wallace_rca12_fa42_y1 = f_u_wallace_rca12_fa42_f_u_wallace_rca12_fa41_y4 & f_u_wallace_rca12_fa42_f_u_wallace_rca12_and_7_6_y0;
  assign f_u_wallace_rca12_fa42_y2 = f_u_wallace_rca12_fa42_y0 ^ f_u_wallace_rca12_fa42_f_u_wallace_rca12_and_6_7_y0;
  assign f_u_wallace_rca12_fa42_y3 = f_u_wallace_rca12_fa42_y0 & f_u_wallace_rca12_fa42_f_u_wallace_rca12_and_6_7_y0;
  assign f_u_wallace_rca12_fa42_y4 = f_u_wallace_rca12_fa42_y1 | f_u_wallace_rca12_fa42_y3;
  assign f_u_wallace_rca12_and_7_7_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_7_7_y0 = f_u_wallace_rca12_and_7_7_a_7 & f_u_wallace_rca12_and_7_7_b_7;
  assign f_u_wallace_rca12_and_6_8_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_6_8_y0 = f_u_wallace_rca12_and_6_8_a_6 & f_u_wallace_rca12_and_6_8_b_8;
  assign f_u_wallace_rca12_fa43_f_u_wallace_rca12_fa42_y4 = f_u_wallace_rca12_fa42_y4;
  assign f_u_wallace_rca12_fa43_f_u_wallace_rca12_and_7_7_y0 = f_u_wallace_rca12_and_7_7_y0;
  assign f_u_wallace_rca12_fa43_f_u_wallace_rca12_and_6_8_y0 = f_u_wallace_rca12_and_6_8_y0;
  assign f_u_wallace_rca12_fa43_y0 = f_u_wallace_rca12_fa43_f_u_wallace_rca12_fa42_y4 ^ f_u_wallace_rca12_fa43_f_u_wallace_rca12_and_7_7_y0;
  assign f_u_wallace_rca12_fa43_y1 = f_u_wallace_rca12_fa43_f_u_wallace_rca12_fa42_y4 & f_u_wallace_rca12_fa43_f_u_wallace_rca12_and_7_7_y0;
  assign f_u_wallace_rca12_fa43_y2 = f_u_wallace_rca12_fa43_y0 ^ f_u_wallace_rca12_fa43_f_u_wallace_rca12_and_6_8_y0;
  assign f_u_wallace_rca12_fa43_y3 = f_u_wallace_rca12_fa43_y0 & f_u_wallace_rca12_fa43_f_u_wallace_rca12_and_6_8_y0;
  assign f_u_wallace_rca12_fa43_y4 = f_u_wallace_rca12_fa43_y1 | f_u_wallace_rca12_fa43_y3;
  assign f_u_wallace_rca12_and_7_8_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_7_8_y0 = f_u_wallace_rca12_and_7_8_a_7 & f_u_wallace_rca12_and_7_8_b_8;
  assign f_u_wallace_rca12_and_6_9_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_6_9_y0 = f_u_wallace_rca12_and_6_9_a_6 & f_u_wallace_rca12_and_6_9_b_9;
  assign f_u_wallace_rca12_fa44_f_u_wallace_rca12_fa43_y4 = f_u_wallace_rca12_fa43_y4;
  assign f_u_wallace_rca12_fa44_f_u_wallace_rca12_and_7_8_y0 = f_u_wallace_rca12_and_7_8_y0;
  assign f_u_wallace_rca12_fa44_f_u_wallace_rca12_and_6_9_y0 = f_u_wallace_rca12_and_6_9_y0;
  assign f_u_wallace_rca12_fa44_y0 = f_u_wallace_rca12_fa44_f_u_wallace_rca12_fa43_y4 ^ f_u_wallace_rca12_fa44_f_u_wallace_rca12_and_7_8_y0;
  assign f_u_wallace_rca12_fa44_y1 = f_u_wallace_rca12_fa44_f_u_wallace_rca12_fa43_y4 & f_u_wallace_rca12_fa44_f_u_wallace_rca12_and_7_8_y0;
  assign f_u_wallace_rca12_fa44_y2 = f_u_wallace_rca12_fa44_y0 ^ f_u_wallace_rca12_fa44_f_u_wallace_rca12_and_6_9_y0;
  assign f_u_wallace_rca12_fa44_y3 = f_u_wallace_rca12_fa44_y0 & f_u_wallace_rca12_fa44_f_u_wallace_rca12_and_6_9_y0;
  assign f_u_wallace_rca12_fa44_y4 = f_u_wallace_rca12_fa44_y1 | f_u_wallace_rca12_fa44_y3;
  assign f_u_wallace_rca12_and_7_9_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_7_9_y0 = f_u_wallace_rca12_and_7_9_a_7 & f_u_wallace_rca12_and_7_9_b_9;
  assign f_u_wallace_rca12_and_6_10_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_6_10_y0 = f_u_wallace_rca12_and_6_10_a_6 & f_u_wallace_rca12_and_6_10_b_10;
  assign f_u_wallace_rca12_fa45_f_u_wallace_rca12_fa44_y4 = f_u_wallace_rca12_fa44_y4;
  assign f_u_wallace_rca12_fa45_f_u_wallace_rca12_and_7_9_y0 = f_u_wallace_rca12_and_7_9_y0;
  assign f_u_wallace_rca12_fa45_f_u_wallace_rca12_and_6_10_y0 = f_u_wallace_rca12_and_6_10_y0;
  assign f_u_wallace_rca12_fa45_y0 = f_u_wallace_rca12_fa45_f_u_wallace_rca12_fa44_y4 ^ f_u_wallace_rca12_fa45_f_u_wallace_rca12_and_7_9_y0;
  assign f_u_wallace_rca12_fa45_y1 = f_u_wallace_rca12_fa45_f_u_wallace_rca12_fa44_y4 & f_u_wallace_rca12_fa45_f_u_wallace_rca12_and_7_9_y0;
  assign f_u_wallace_rca12_fa45_y2 = f_u_wallace_rca12_fa45_y0 ^ f_u_wallace_rca12_fa45_f_u_wallace_rca12_and_6_10_y0;
  assign f_u_wallace_rca12_fa45_y3 = f_u_wallace_rca12_fa45_y0 & f_u_wallace_rca12_fa45_f_u_wallace_rca12_and_6_10_y0;
  assign f_u_wallace_rca12_fa45_y4 = f_u_wallace_rca12_fa45_y1 | f_u_wallace_rca12_fa45_y3;
  assign f_u_wallace_rca12_and_7_10_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_7_10_y0 = f_u_wallace_rca12_and_7_10_a_7 & f_u_wallace_rca12_and_7_10_b_10;
  assign f_u_wallace_rca12_and_6_11_a_6 = a_6;
  assign f_u_wallace_rca12_and_6_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_6_11_y0 = f_u_wallace_rca12_and_6_11_a_6 & f_u_wallace_rca12_and_6_11_b_11;
  assign f_u_wallace_rca12_fa46_f_u_wallace_rca12_fa45_y4 = f_u_wallace_rca12_fa45_y4;
  assign f_u_wallace_rca12_fa46_f_u_wallace_rca12_and_7_10_y0 = f_u_wallace_rca12_and_7_10_y0;
  assign f_u_wallace_rca12_fa46_f_u_wallace_rca12_and_6_11_y0 = f_u_wallace_rca12_and_6_11_y0;
  assign f_u_wallace_rca12_fa46_y0 = f_u_wallace_rca12_fa46_f_u_wallace_rca12_fa45_y4 ^ f_u_wallace_rca12_fa46_f_u_wallace_rca12_and_7_10_y0;
  assign f_u_wallace_rca12_fa46_y1 = f_u_wallace_rca12_fa46_f_u_wallace_rca12_fa45_y4 & f_u_wallace_rca12_fa46_f_u_wallace_rca12_and_7_10_y0;
  assign f_u_wallace_rca12_fa46_y2 = f_u_wallace_rca12_fa46_y0 ^ f_u_wallace_rca12_fa46_f_u_wallace_rca12_and_6_11_y0;
  assign f_u_wallace_rca12_fa46_y3 = f_u_wallace_rca12_fa46_y0 & f_u_wallace_rca12_fa46_f_u_wallace_rca12_and_6_11_y0;
  assign f_u_wallace_rca12_fa46_y4 = f_u_wallace_rca12_fa46_y1 | f_u_wallace_rca12_fa46_y3;
  assign f_u_wallace_rca12_and_7_11_a_7 = a_7;
  assign f_u_wallace_rca12_and_7_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_7_11_y0 = f_u_wallace_rca12_and_7_11_a_7 & f_u_wallace_rca12_and_7_11_b_11;
  assign f_u_wallace_rca12_fa47_f_u_wallace_rca12_fa46_y4 = f_u_wallace_rca12_fa46_y4;
  assign f_u_wallace_rca12_fa47_f_u_wallace_rca12_and_7_11_y0 = f_u_wallace_rca12_and_7_11_y0;
  assign f_u_wallace_rca12_fa47_f_u_wallace_rca12_fa15_y2 = f_u_wallace_rca12_fa15_y2;
  assign f_u_wallace_rca12_fa47_y0 = f_u_wallace_rca12_fa47_f_u_wallace_rca12_fa46_y4 ^ f_u_wallace_rca12_fa47_f_u_wallace_rca12_and_7_11_y0;
  assign f_u_wallace_rca12_fa47_y1 = f_u_wallace_rca12_fa47_f_u_wallace_rca12_fa46_y4 & f_u_wallace_rca12_fa47_f_u_wallace_rca12_and_7_11_y0;
  assign f_u_wallace_rca12_fa47_y2 = f_u_wallace_rca12_fa47_y0 ^ f_u_wallace_rca12_fa47_f_u_wallace_rca12_fa15_y2;
  assign f_u_wallace_rca12_fa47_y3 = f_u_wallace_rca12_fa47_y0 & f_u_wallace_rca12_fa47_f_u_wallace_rca12_fa15_y2;
  assign f_u_wallace_rca12_fa47_y4 = f_u_wallace_rca12_fa47_y1 | f_u_wallace_rca12_fa47_y3;
  assign f_u_wallace_rca12_ha3_f_u_wallace_rca12_fa2_y2 = f_u_wallace_rca12_fa2_y2;
  assign f_u_wallace_rca12_ha3_f_u_wallace_rca12_fa19_y2 = f_u_wallace_rca12_fa19_y2;
  assign f_u_wallace_rca12_ha3_y0 = f_u_wallace_rca12_ha3_f_u_wallace_rca12_fa2_y2 ^ f_u_wallace_rca12_ha3_f_u_wallace_rca12_fa19_y2;
  assign f_u_wallace_rca12_ha3_y1 = f_u_wallace_rca12_ha3_f_u_wallace_rca12_fa2_y2 & f_u_wallace_rca12_ha3_f_u_wallace_rca12_fa19_y2;
  assign f_u_wallace_rca12_and_0_6_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_0_6_y0 = f_u_wallace_rca12_and_0_6_a_0 & f_u_wallace_rca12_and_0_6_b_6;
  assign f_u_wallace_rca12_fa48_f_u_wallace_rca12_ha3_y1 = f_u_wallace_rca12_ha3_y1;
  assign f_u_wallace_rca12_fa48_f_u_wallace_rca12_and_0_6_y0 = f_u_wallace_rca12_and_0_6_y0;
  assign f_u_wallace_rca12_fa48_f_u_wallace_rca12_fa3_y2 = f_u_wallace_rca12_fa3_y2;
  assign f_u_wallace_rca12_fa48_y0 = f_u_wallace_rca12_fa48_f_u_wallace_rca12_ha3_y1 ^ f_u_wallace_rca12_fa48_f_u_wallace_rca12_and_0_6_y0;
  assign f_u_wallace_rca12_fa48_y1 = f_u_wallace_rca12_fa48_f_u_wallace_rca12_ha3_y1 & f_u_wallace_rca12_fa48_f_u_wallace_rca12_and_0_6_y0;
  assign f_u_wallace_rca12_fa48_y2 = f_u_wallace_rca12_fa48_y0 ^ f_u_wallace_rca12_fa48_f_u_wallace_rca12_fa3_y2;
  assign f_u_wallace_rca12_fa48_y3 = f_u_wallace_rca12_fa48_y0 & f_u_wallace_rca12_fa48_f_u_wallace_rca12_fa3_y2;
  assign f_u_wallace_rca12_fa48_y4 = f_u_wallace_rca12_fa48_y1 | f_u_wallace_rca12_fa48_y3;
  assign f_u_wallace_rca12_and_1_6_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_1_6_y0 = f_u_wallace_rca12_and_1_6_a_1 & f_u_wallace_rca12_and_1_6_b_6;
  assign f_u_wallace_rca12_and_0_7_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_0_7_y0 = f_u_wallace_rca12_and_0_7_a_0 & f_u_wallace_rca12_and_0_7_b_7;
  assign f_u_wallace_rca12_fa49_f_u_wallace_rca12_fa48_y4 = f_u_wallace_rca12_fa48_y4;
  assign f_u_wallace_rca12_fa49_f_u_wallace_rca12_and_1_6_y0 = f_u_wallace_rca12_and_1_6_y0;
  assign f_u_wallace_rca12_fa49_f_u_wallace_rca12_and_0_7_y0 = f_u_wallace_rca12_and_0_7_y0;
  assign f_u_wallace_rca12_fa49_y0 = f_u_wallace_rca12_fa49_f_u_wallace_rca12_fa48_y4 ^ f_u_wallace_rca12_fa49_f_u_wallace_rca12_and_1_6_y0;
  assign f_u_wallace_rca12_fa49_y1 = f_u_wallace_rca12_fa49_f_u_wallace_rca12_fa48_y4 & f_u_wallace_rca12_fa49_f_u_wallace_rca12_and_1_6_y0;
  assign f_u_wallace_rca12_fa49_y2 = f_u_wallace_rca12_fa49_y0 ^ f_u_wallace_rca12_fa49_f_u_wallace_rca12_and_0_7_y0;
  assign f_u_wallace_rca12_fa49_y3 = f_u_wallace_rca12_fa49_y0 & f_u_wallace_rca12_fa49_f_u_wallace_rca12_and_0_7_y0;
  assign f_u_wallace_rca12_fa49_y4 = f_u_wallace_rca12_fa49_y1 | f_u_wallace_rca12_fa49_y3;
  assign f_u_wallace_rca12_and_2_6_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_2_6_y0 = f_u_wallace_rca12_and_2_6_a_2 & f_u_wallace_rca12_and_2_6_b_6;
  assign f_u_wallace_rca12_and_1_7_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_1_7_y0 = f_u_wallace_rca12_and_1_7_a_1 & f_u_wallace_rca12_and_1_7_b_7;
  assign f_u_wallace_rca12_fa50_f_u_wallace_rca12_fa49_y4 = f_u_wallace_rca12_fa49_y4;
  assign f_u_wallace_rca12_fa50_f_u_wallace_rca12_and_2_6_y0 = f_u_wallace_rca12_and_2_6_y0;
  assign f_u_wallace_rca12_fa50_f_u_wallace_rca12_and_1_7_y0 = f_u_wallace_rca12_and_1_7_y0;
  assign f_u_wallace_rca12_fa50_y0 = f_u_wallace_rca12_fa50_f_u_wallace_rca12_fa49_y4 ^ f_u_wallace_rca12_fa50_f_u_wallace_rca12_and_2_6_y0;
  assign f_u_wallace_rca12_fa50_y1 = f_u_wallace_rca12_fa50_f_u_wallace_rca12_fa49_y4 & f_u_wallace_rca12_fa50_f_u_wallace_rca12_and_2_6_y0;
  assign f_u_wallace_rca12_fa50_y2 = f_u_wallace_rca12_fa50_y0 ^ f_u_wallace_rca12_fa50_f_u_wallace_rca12_and_1_7_y0;
  assign f_u_wallace_rca12_fa50_y3 = f_u_wallace_rca12_fa50_y0 & f_u_wallace_rca12_fa50_f_u_wallace_rca12_and_1_7_y0;
  assign f_u_wallace_rca12_fa50_y4 = f_u_wallace_rca12_fa50_y1 | f_u_wallace_rca12_fa50_y3;
  assign f_u_wallace_rca12_and_3_6_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_3_6_y0 = f_u_wallace_rca12_and_3_6_a_3 & f_u_wallace_rca12_and_3_6_b_6;
  assign f_u_wallace_rca12_and_2_7_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_2_7_y0 = f_u_wallace_rca12_and_2_7_a_2 & f_u_wallace_rca12_and_2_7_b_7;
  assign f_u_wallace_rca12_fa51_f_u_wallace_rca12_fa50_y4 = f_u_wallace_rca12_fa50_y4;
  assign f_u_wallace_rca12_fa51_f_u_wallace_rca12_and_3_6_y0 = f_u_wallace_rca12_and_3_6_y0;
  assign f_u_wallace_rca12_fa51_f_u_wallace_rca12_and_2_7_y0 = f_u_wallace_rca12_and_2_7_y0;
  assign f_u_wallace_rca12_fa51_y0 = f_u_wallace_rca12_fa51_f_u_wallace_rca12_fa50_y4 ^ f_u_wallace_rca12_fa51_f_u_wallace_rca12_and_3_6_y0;
  assign f_u_wallace_rca12_fa51_y1 = f_u_wallace_rca12_fa51_f_u_wallace_rca12_fa50_y4 & f_u_wallace_rca12_fa51_f_u_wallace_rca12_and_3_6_y0;
  assign f_u_wallace_rca12_fa51_y2 = f_u_wallace_rca12_fa51_y0 ^ f_u_wallace_rca12_fa51_f_u_wallace_rca12_and_2_7_y0;
  assign f_u_wallace_rca12_fa51_y3 = f_u_wallace_rca12_fa51_y0 & f_u_wallace_rca12_fa51_f_u_wallace_rca12_and_2_7_y0;
  assign f_u_wallace_rca12_fa51_y4 = f_u_wallace_rca12_fa51_y1 | f_u_wallace_rca12_fa51_y3;
  assign f_u_wallace_rca12_and_4_6_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_4_6_y0 = f_u_wallace_rca12_and_4_6_a_4 & f_u_wallace_rca12_and_4_6_b_6;
  assign f_u_wallace_rca12_and_3_7_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_3_7_y0 = f_u_wallace_rca12_and_3_7_a_3 & f_u_wallace_rca12_and_3_7_b_7;
  assign f_u_wallace_rca12_fa52_f_u_wallace_rca12_fa51_y4 = f_u_wallace_rca12_fa51_y4;
  assign f_u_wallace_rca12_fa52_f_u_wallace_rca12_and_4_6_y0 = f_u_wallace_rca12_and_4_6_y0;
  assign f_u_wallace_rca12_fa52_f_u_wallace_rca12_and_3_7_y0 = f_u_wallace_rca12_and_3_7_y0;
  assign f_u_wallace_rca12_fa52_y0 = f_u_wallace_rca12_fa52_f_u_wallace_rca12_fa51_y4 ^ f_u_wallace_rca12_fa52_f_u_wallace_rca12_and_4_6_y0;
  assign f_u_wallace_rca12_fa52_y1 = f_u_wallace_rca12_fa52_f_u_wallace_rca12_fa51_y4 & f_u_wallace_rca12_fa52_f_u_wallace_rca12_and_4_6_y0;
  assign f_u_wallace_rca12_fa52_y2 = f_u_wallace_rca12_fa52_y0 ^ f_u_wallace_rca12_fa52_f_u_wallace_rca12_and_3_7_y0;
  assign f_u_wallace_rca12_fa52_y3 = f_u_wallace_rca12_fa52_y0 & f_u_wallace_rca12_fa52_f_u_wallace_rca12_and_3_7_y0;
  assign f_u_wallace_rca12_fa52_y4 = f_u_wallace_rca12_fa52_y1 | f_u_wallace_rca12_fa52_y3;
  assign f_u_wallace_rca12_and_5_6_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_6_b_6 = b_6;
  assign f_u_wallace_rca12_and_5_6_y0 = f_u_wallace_rca12_and_5_6_a_5 & f_u_wallace_rca12_and_5_6_b_6;
  assign f_u_wallace_rca12_and_4_7_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_4_7_y0 = f_u_wallace_rca12_and_4_7_a_4 & f_u_wallace_rca12_and_4_7_b_7;
  assign f_u_wallace_rca12_fa53_f_u_wallace_rca12_fa52_y4 = f_u_wallace_rca12_fa52_y4;
  assign f_u_wallace_rca12_fa53_f_u_wallace_rca12_and_5_6_y0 = f_u_wallace_rca12_and_5_6_y0;
  assign f_u_wallace_rca12_fa53_f_u_wallace_rca12_and_4_7_y0 = f_u_wallace_rca12_and_4_7_y0;
  assign f_u_wallace_rca12_fa53_y0 = f_u_wallace_rca12_fa53_f_u_wallace_rca12_fa52_y4 ^ f_u_wallace_rca12_fa53_f_u_wallace_rca12_and_5_6_y0;
  assign f_u_wallace_rca12_fa53_y1 = f_u_wallace_rca12_fa53_f_u_wallace_rca12_fa52_y4 & f_u_wallace_rca12_fa53_f_u_wallace_rca12_and_5_6_y0;
  assign f_u_wallace_rca12_fa53_y2 = f_u_wallace_rca12_fa53_y0 ^ f_u_wallace_rca12_fa53_f_u_wallace_rca12_and_4_7_y0;
  assign f_u_wallace_rca12_fa53_y3 = f_u_wallace_rca12_fa53_y0 & f_u_wallace_rca12_fa53_f_u_wallace_rca12_and_4_7_y0;
  assign f_u_wallace_rca12_fa53_y4 = f_u_wallace_rca12_fa53_y1 | f_u_wallace_rca12_fa53_y3;
  assign f_u_wallace_rca12_and_5_7_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_7_b_7 = b_7;
  assign f_u_wallace_rca12_and_5_7_y0 = f_u_wallace_rca12_and_5_7_a_5 & f_u_wallace_rca12_and_5_7_b_7;
  assign f_u_wallace_rca12_and_4_8_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_4_8_y0 = f_u_wallace_rca12_and_4_8_a_4 & f_u_wallace_rca12_and_4_8_b_8;
  assign f_u_wallace_rca12_fa54_f_u_wallace_rca12_fa53_y4 = f_u_wallace_rca12_fa53_y4;
  assign f_u_wallace_rca12_fa54_f_u_wallace_rca12_and_5_7_y0 = f_u_wallace_rca12_and_5_7_y0;
  assign f_u_wallace_rca12_fa54_f_u_wallace_rca12_and_4_8_y0 = f_u_wallace_rca12_and_4_8_y0;
  assign f_u_wallace_rca12_fa54_y0 = f_u_wallace_rca12_fa54_f_u_wallace_rca12_fa53_y4 ^ f_u_wallace_rca12_fa54_f_u_wallace_rca12_and_5_7_y0;
  assign f_u_wallace_rca12_fa54_y1 = f_u_wallace_rca12_fa54_f_u_wallace_rca12_fa53_y4 & f_u_wallace_rca12_fa54_f_u_wallace_rca12_and_5_7_y0;
  assign f_u_wallace_rca12_fa54_y2 = f_u_wallace_rca12_fa54_y0 ^ f_u_wallace_rca12_fa54_f_u_wallace_rca12_and_4_8_y0;
  assign f_u_wallace_rca12_fa54_y3 = f_u_wallace_rca12_fa54_y0 & f_u_wallace_rca12_fa54_f_u_wallace_rca12_and_4_8_y0;
  assign f_u_wallace_rca12_fa54_y4 = f_u_wallace_rca12_fa54_y1 | f_u_wallace_rca12_fa54_y3;
  assign f_u_wallace_rca12_and_5_8_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_5_8_y0 = f_u_wallace_rca12_and_5_8_a_5 & f_u_wallace_rca12_and_5_8_b_8;
  assign f_u_wallace_rca12_and_4_9_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_4_9_y0 = f_u_wallace_rca12_and_4_9_a_4 & f_u_wallace_rca12_and_4_9_b_9;
  assign f_u_wallace_rca12_fa55_f_u_wallace_rca12_fa54_y4 = f_u_wallace_rca12_fa54_y4;
  assign f_u_wallace_rca12_fa55_f_u_wallace_rca12_and_5_8_y0 = f_u_wallace_rca12_and_5_8_y0;
  assign f_u_wallace_rca12_fa55_f_u_wallace_rca12_and_4_9_y0 = f_u_wallace_rca12_and_4_9_y0;
  assign f_u_wallace_rca12_fa55_y0 = f_u_wallace_rca12_fa55_f_u_wallace_rca12_fa54_y4 ^ f_u_wallace_rca12_fa55_f_u_wallace_rca12_and_5_8_y0;
  assign f_u_wallace_rca12_fa55_y1 = f_u_wallace_rca12_fa55_f_u_wallace_rca12_fa54_y4 & f_u_wallace_rca12_fa55_f_u_wallace_rca12_and_5_8_y0;
  assign f_u_wallace_rca12_fa55_y2 = f_u_wallace_rca12_fa55_y0 ^ f_u_wallace_rca12_fa55_f_u_wallace_rca12_and_4_9_y0;
  assign f_u_wallace_rca12_fa55_y3 = f_u_wallace_rca12_fa55_y0 & f_u_wallace_rca12_fa55_f_u_wallace_rca12_and_4_9_y0;
  assign f_u_wallace_rca12_fa55_y4 = f_u_wallace_rca12_fa55_y1 | f_u_wallace_rca12_fa55_y3;
  assign f_u_wallace_rca12_and_5_9_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_5_9_y0 = f_u_wallace_rca12_and_5_9_a_5 & f_u_wallace_rca12_and_5_9_b_9;
  assign f_u_wallace_rca12_and_4_10_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_4_10_y0 = f_u_wallace_rca12_and_4_10_a_4 & f_u_wallace_rca12_and_4_10_b_10;
  assign f_u_wallace_rca12_fa56_f_u_wallace_rca12_fa55_y4 = f_u_wallace_rca12_fa55_y4;
  assign f_u_wallace_rca12_fa56_f_u_wallace_rca12_and_5_9_y0 = f_u_wallace_rca12_and_5_9_y0;
  assign f_u_wallace_rca12_fa56_f_u_wallace_rca12_and_4_10_y0 = f_u_wallace_rca12_and_4_10_y0;
  assign f_u_wallace_rca12_fa56_y0 = f_u_wallace_rca12_fa56_f_u_wallace_rca12_fa55_y4 ^ f_u_wallace_rca12_fa56_f_u_wallace_rca12_and_5_9_y0;
  assign f_u_wallace_rca12_fa56_y1 = f_u_wallace_rca12_fa56_f_u_wallace_rca12_fa55_y4 & f_u_wallace_rca12_fa56_f_u_wallace_rca12_and_5_9_y0;
  assign f_u_wallace_rca12_fa56_y2 = f_u_wallace_rca12_fa56_y0 ^ f_u_wallace_rca12_fa56_f_u_wallace_rca12_and_4_10_y0;
  assign f_u_wallace_rca12_fa56_y3 = f_u_wallace_rca12_fa56_y0 & f_u_wallace_rca12_fa56_f_u_wallace_rca12_and_4_10_y0;
  assign f_u_wallace_rca12_fa56_y4 = f_u_wallace_rca12_fa56_y1 | f_u_wallace_rca12_fa56_y3;
  assign f_u_wallace_rca12_and_5_10_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_5_10_y0 = f_u_wallace_rca12_and_5_10_a_5 & f_u_wallace_rca12_and_5_10_b_10;
  assign f_u_wallace_rca12_and_4_11_a_4 = a_4;
  assign f_u_wallace_rca12_and_4_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_4_11_y0 = f_u_wallace_rca12_and_4_11_a_4 & f_u_wallace_rca12_and_4_11_b_11;
  assign f_u_wallace_rca12_fa57_f_u_wallace_rca12_fa56_y4 = f_u_wallace_rca12_fa56_y4;
  assign f_u_wallace_rca12_fa57_f_u_wallace_rca12_and_5_10_y0 = f_u_wallace_rca12_and_5_10_y0;
  assign f_u_wallace_rca12_fa57_f_u_wallace_rca12_and_4_11_y0 = f_u_wallace_rca12_and_4_11_y0;
  assign f_u_wallace_rca12_fa57_y0 = f_u_wallace_rca12_fa57_f_u_wallace_rca12_fa56_y4 ^ f_u_wallace_rca12_fa57_f_u_wallace_rca12_and_5_10_y0;
  assign f_u_wallace_rca12_fa57_y1 = f_u_wallace_rca12_fa57_f_u_wallace_rca12_fa56_y4 & f_u_wallace_rca12_fa57_f_u_wallace_rca12_and_5_10_y0;
  assign f_u_wallace_rca12_fa57_y2 = f_u_wallace_rca12_fa57_y0 ^ f_u_wallace_rca12_fa57_f_u_wallace_rca12_and_4_11_y0;
  assign f_u_wallace_rca12_fa57_y3 = f_u_wallace_rca12_fa57_y0 & f_u_wallace_rca12_fa57_f_u_wallace_rca12_and_4_11_y0;
  assign f_u_wallace_rca12_fa57_y4 = f_u_wallace_rca12_fa57_y1 | f_u_wallace_rca12_fa57_y3;
  assign f_u_wallace_rca12_and_5_11_a_5 = a_5;
  assign f_u_wallace_rca12_and_5_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_5_11_y0 = f_u_wallace_rca12_and_5_11_a_5 & f_u_wallace_rca12_and_5_11_b_11;
  assign f_u_wallace_rca12_fa58_f_u_wallace_rca12_fa57_y4 = f_u_wallace_rca12_fa57_y4;
  assign f_u_wallace_rca12_fa58_f_u_wallace_rca12_and_5_11_y0 = f_u_wallace_rca12_and_5_11_y0;
  assign f_u_wallace_rca12_fa58_f_u_wallace_rca12_fa13_y2 = f_u_wallace_rca12_fa13_y2;
  assign f_u_wallace_rca12_fa58_y0 = f_u_wallace_rca12_fa58_f_u_wallace_rca12_fa57_y4 ^ f_u_wallace_rca12_fa58_f_u_wallace_rca12_and_5_11_y0;
  assign f_u_wallace_rca12_fa58_y1 = f_u_wallace_rca12_fa58_f_u_wallace_rca12_fa57_y4 & f_u_wallace_rca12_fa58_f_u_wallace_rca12_and_5_11_y0;
  assign f_u_wallace_rca12_fa58_y2 = f_u_wallace_rca12_fa58_y0 ^ f_u_wallace_rca12_fa58_f_u_wallace_rca12_fa13_y2;
  assign f_u_wallace_rca12_fa58_y3 = f_u_wallace_rca12_fa58_y0 & f_u_wallace_rca12_fa58_f_u_wallace_rca12_fa13_y2;
  assign f_u_wallace_rca12_fa58_y4 = f_u_wallace_rca12_fa58_y1 | f_u_wallace_rca12_fa58_y3;
  assign f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa58_y4 = f_u_wallace_rca12_fa58_y4;
  assign f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa14_y2 = f_u_wallace_rca12_fa14_y2;
  assign f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa31_y2 = f_u_wallace_rca12_fa31_y2;
  assign f_u_wallace_rca12_fa59_y0 = f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa58_y4 ^ f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa14_y2;
  assign f_u_wallace_rca12_fa59_y1 = f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa58_y4 & f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa14_y2;
  assign f_u_wallace_rca12_fa59_y2 = f_u_wallace_rca12_fa59_y0 ^ f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa31_y2;
  assign f_u_wallace_rca12_fa59_y3 = f_u_wallace_rca12_fa59_y0 & f_u_wallace_rca12_fa59_f_u_wallace_rca12_fa31_y2;
  assign f_u_wallace_rca12_fa59_y4 = f_u_wallace_rca12_fa59_y1 | f_u_wallace_rca12_fa59_y3;
  assign f_u_wallace_rca12_ha4_f_u_wallace_rca12_fa20_y2 = f_u_wallace_rca12_fa20_y2;
  assign f_u_wallace_rca12_ha4_f_u_wallace_rca12_fa35_y2 = f_u_wallace_rca12_fa35_y2;
  assign f_u_wallace_rca12_ha4_y0 = f_u_wallace_rca12_ha4_f_u_wallace_rca12_fa20_y2 ^ f_u_wallace_rca12_ha4_f_u_wallace_rca12_fa35_y2;
  assign f_u_wallace_rca12_ha4_y1 = f_u_wallace_rca12_ha4_f_u_wallace_rca12_fa20_y2 & f_u_wallace_rca12_ha4_f_u_wallace_rca12_fa35_y2;
  assign f_u_wallace_rca12_fa60_f_u_wallace_rca12_ha4_y1 = f_u_wallace_rca12_ha4_y1;
  assign f_u_wallace_rca12_fa60_f_u_wallace_rca12_fa4_y2 = f_u_wallace_rca12_fa4_y2;
  assign f_u_wallace_rca12_fa60_f_u_wallace_rca12_fa21_y2 = f_u_wallace_rca12_fa21_y2;
  assign f_u_wallace_rca12_fa60_y0 = f_u_wallace_rca12_fa60_f_u_wallace_rca12_ha4_y1 ^ f_u_wallace_rca12_fa60_f_u_wallace_rca12_fa4_y2;
  assign f_u_wallace_rca12_fa60_y1 = f_u_wallace_rca12_fa60_f_u_wallace_rca12_ha4_y1 & f_u_wallace_rca12_fa60_f_u_wallace_rca12_fa4_y2;
  assign f_u_wallace_rca12_fa60_y2 = f_u_wallace_rca12_fa60_y0 ^ f_u_wallace_rca12_fa60_f_u_wallace_rca12_fa21_y2;
  assign f_u_wallace_rca12_fa60_y3 = f_u_wallace_rca12_fa60_y0 & f_u_wallace_rca12_fa60_f_u_wallace_rca12_fa21_y2;
  assign f_u_wallace_rca12_fa60_y4 = f_u_wallace_rca12_fa60_y1 | f_u_wallace_rca12_fa60_y3;
  assign f_u_wallace_rca12_and_0_8_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_0_8_y0 = f_u_wallace_rca12_and_0_8_a_0 & f_u_wallace_rca12_and_0_8_b_8;
  assign f_u_wallace_rca12_fa61_f_u_wallace_rca12_fa60_y4 = f_u_wallace_rca12_fa60_y4;
  assign f_u_wallace_rca12_fa61_f_u_wallace_rca12_and_0_8_y0 = f_u_wallace_rca12_and_0_8_y0;
  assign f_u_wallace_rca12_fa61_f_u_wallace_rca12_fa5_y2 = f_u_wallace_rca12_fa5_y2;
  assign f_u_wallace_rca12_fa61_y0 = f_u_wallace_rca12_fa61_f_u_wallace_rca12_fa60_y4 ^ f_u_wallace_rca12_fa61_f_u_wallace_rca12_and_0_8_y0;
  assign f_u_wallace_rca12_fa61_y1 = f_u_wallace_rca12_fa61_f_u_wallace_rca12_fa60_y4 & f_u_wallace_rca12_fa61_f_u_wallace_rca12_and_0_8_y0;
  assign f_u_wallace_rca12_fa61_y2 = f_u_wallace_rca12_fa61_y0 ^ f_u_wallace_rca12_fa61_f_u_wallace_rca12_fa5_y2;
  assign f_u_wallace_rca12_fa61_y3 = f_u_wallace_rca12_fa61_y0 & f_u_wallace_rca12_fa61_f_u_wallace_rca12_fa5_y2;
  assign f_u_wallace_rca12_fa61_y4 = f_u_wallace_rca12_fa61_y1 | f_u_wallace_rca12_fa61_y3;
  assign f_u_wallace_rca12_and_1_8_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_1_8_y0 = f_u_wallace_rca12_and_1_8_a_1 & f_u_wallace_rca12_and_1_8_b_8;
  assign f_u_wallace_rca12_and_0_9_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_0_9_y0 = f_u_wallace_rca12_and_0_9_a_0 & f_u_wallace_rca12_and_0_9_b_9;
  assign f_u_wallace_rca12_fa62_f_u_wallace_rca12_fa61_y4 = f_u_wallace_rca12_fa61_y4;
  assign f_u_wallace_rca12_fa62_f_u_wallace_rca12_and_1_8_y0 = f_u_wallace_rca12_and_1_8_y0;
  assign f_u_wallace_rca12_fa62_f_u_wallace_rca12_and_0_9_y0 = f_u_wallace_rca12_and_0_9_y0;
  assign f_u_wallace_rca12_fa62_y0 = f_u_wallace_rca12_fa62_f_u_wallace_rca12_fa61_y4 ^ f_u_wallace_rca12_fa62_f_u_wallace_rca12_and_1_8_y0;
  assign f_u_wallace_rca12_fa62_y1 = f_u_wallace_rca12_fa62_f_u_wallace_rca12_fa61_y4 & f_u_wallace_rca12_fa62_f_u_wallace_rca12_and_1_8_y0;
  assign f_u_wallace_rca12_fa62_y2 = f_u_wallace_rca12_fa62_y0 ^ f_u_wallace_rca12_fa62_f_u_wallace_rca12_and_0_9_y0;
  assign f_u_wallace_rca12_fa62_y3 = f_u_wallace_rca12_fa62_y0 & f_u_wallace_rca12_fa62_f_u_wallace_rca12_and_0_9_y0;
  assign f_u_wallace_rca12_fa62_y4 = f_u_wallace_rca12_fa62_y1 | f_u_wallace_rca12_fa62_y3;
  assign f_u_wallace_rca12_and_2_8_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_2_8_y0 = f_u_wallace_rca12_and_2_8_a_2 & f_u_wallace_rca12_and_2_8_b_8;
  assign f_u_wallace_rca12_and_1_9_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_1_9_y0 = f_u_wallace_rca12_and_1_9_a_1 & f_u_wallace_rca12_and_1_9_b_9;
  assign f_u_wallace_rca12_fa63_f_u_wallace_rca12_fa62_y4 = f_u_wallace_rca12_fa62_y4;
  assign f_u_wallace_rca12_fa63_f_u_wallace_rca12_and_2_8_y0 = f_u_wallace_rca12_and_2_8_y0;
  assign f_u_wallace_rca12_fa63_f_u_wallace_rca12_and_1_9_y0 = f_u_wallace_rca12_and_1_9_y0;
  assign f_u_wallace_rca12_fa63_y0 = f_u_wallace_rca12_fa63_f_u_wallace_rca12_fa62_y4 ^ f_u_wallace_rca12_fa63_f_u_wallace_rca12_and_2_8_y0;
  assign f_u_wallace_rca12_fa63_y1 = f_u_wallace_rca12_fa63_f_u_wallace_rca12_fa62_y4 & f_u_wallace_rca12_fa63_f_u_wallace_rca12_and_2_8_y0;
  assign f_u_wallace_rca12_fa63_y2 = f_u_wallace_rca12_fa63_y0 ^ f_u_wallace_rca12_fa63_f_u_wallace_rca12_and_1_9_y0;
  assign f_u_wallace_rca12_fa63_y3 = f_u_wallace_rca12_fa63_y0 & f_u_wallace_rca12_fa63_f_u_wallace_rca12_and_1_9_y0;
  assign f_u_wallace_rca12_fa63_y4 = f_u_wallace_rca12_fa63_y1 | f_u_wallace_rca12_fa63_y3;
  assign f_u_wallace_rca12_and_3_8_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_8_b_8 = b_8;
  assign f_u_wallace_rca12_and_3_8_y0 = f_u_wallace_rca12_and_3_8_a_3 & f_u_wallace_rca12_and_3_8_b_8;
  assign f_u_wallace_rca12_and_2_9_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_2_9_y0 = f_u_wallace_rca12_and_2_9_a_2 & f_u_wallace_rca12_and_2_9_b_9;
  assign f_u_wallace_rca12_fa64_f_u_wallace_rca12_fa63_y4 = f_u_wallace_rca12_fa63_y4;
  assign f_u_wallace_rca12_fa64_f_u_wallace_rca12_and_3_8_y0 = f_u_wallace_rca12_and_3_8_y0;
  assign f_u_wallace_rca12_fa64_f_u_wallace_rca12_and_2_9_y0 = f_u_wallace_rca12_and_2_9_y0;
  assign f_u_wallace_rca12_fa64_y0 = f_u_wallace_rca12_fa64_f_u_wallace_rca12_fa63_y4 ^ f_u_wallace_rca12_fa64_f_u_wallace_rca12_and_3_8_y0;
  assign f_u_wallace_rca12_fa64_y1 = f_u_wallace_rca12_fa64_f_u_wallace_rca12_fa63_y4 & f_u_wallace_rca12_fa64_f_u_wallace_rca12_and_3_8_y0;
  assign f_u_wallace_rca12_fa64_y2 = f_u_wallace_rca12_fa64_y0 ^ f_u_wallace_rca12_fa64_f_u_wallace_rca12_and_2_9_y0;
  assign f_u_wallace_rca12_fa64_y3 = f_u_wallace_rca12_fa64_y0 & f_u_wallace_rca12_fa64_f_u_wallace_rca12_and_2_9_y0;
  assign f_u_wallace_rca12_fa64_y4 = f_u_wallace_rca12_fa64_y1 | f_u_wallace_rca12_fa64_y3;
  assign f_u_wallace_rca12_and_3_9_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_9_b_9 = b_9;
  assign f_u_wallace_rca12_and_3_9_y0 = f_u_wallace_rca12_and_3_9_a_3 & f_u_wallace_rca12_and_3_9_b_9;
  assign f_u_wallace_rca12_and_2_10_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_2_10_y0 = f_u_wallace_rca12_and_2_10_a_2 & f_u_wallace_rca12_and_2_10_b_10;
  assign f_u_wallace_rca12_fa65_f_u_wallace_rca12_fa64_y4 = f_u_wallace_rca12_fa64_y4;
  assign f_u_wallace_rca12_fa65_f_u_wallace_rca12_and_3_9_y0 = f_u_wallace_rca12_and_3_9_y0;
  assign f_u_wallace_rca12_fa65_f_u_wallace_rca12_and_2_10_y0 = f_u_wallace_rca12_and_2_10_y0;
  assign f_u_wallace_rca12_fa65_y0 = f_u_wallace_rca12_fa65_f_u_wallace_rca12_fa64_y4 ^ f_u_wallace_rca12_fa65_f_u_wallace_rca12_and_3_9_y0;
  assign f_u_wallace_rca12_fa65_y1 = f_u_wallace_rca12_fa65_f_u_wallace_rca12_fa64_y4 & f_u_wallace_rca12_fa65_f_u_wallace_rca12_and_3_9_y0;
  assign f_u_wallace_rca12_fa65_y2 = f_u_wallace_rca12_fa65_y0 ^ f_u_wallace_rca12_fa65_f_u_wallace_rca12_and_2_10_y0;
  assign f_u_wallace_rca12_fa65_y3 = f_u_wallace_rca12_fa65_y0 & f_u_wallace_rca12_fa65_f_u_wallace_rca12_and_2_10_y0;
  assign f_u_wallace_rca12_fa65_y4 = f_u_wallace_rca12_fa65_y1 | f_u_wallace_rca12_fa65_y3;
  assign f_u_wallace_rca12_and_3_10_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_3_10_y0 = f_u_wallace_rca12_and_3_10_a_3 & f_u_wallace_rca12_and_3_10_b_10;
  assign f_u_wallace_rca12_and_2_11_a_2 = a_2;
  assign f_u_wallace_rca12_and_2_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_2_11_y0 = f_u_wallace_rca12_and_2_11_a_2 & f_u_wallace_rca12_and_2_11_b_11;
  assign f_u_wallace_rca12_fa66_f_u_wallace_rca12_fa65_y4 = f_u_wallace_rca12_fa65_y4;
  assign f_u_wallace_rca12_fa66_f_u_wallace_rca12_and_3_10_y0 = f_u_wallace_rca12_and_3_10_y0;
  assign f_u_wallace_rca12_fa66_f_u_wallace_rca12_and_2_11_y0 = f_u_wallace_rca12_and_2_11_y0;
  assign f_u_wallace_rca12_fa66_y0 = f_u_wallace_rca12_fa66_f_u_wallace_rca12_fa65_y4 ^ f_u_wallace_rca12_fa66_f_u_wallace_rca12_and_3_10_y0;
  assign f_u_wallace_rca12_fa66_y1 = f_u_wallace_rca12_fa66_f_u_wallace_rca12_fa65_y4 & f_u_wallace_rca12_fa66_f_u_wallace_rca12_and_3_10_y0;
  assign f_u_wallace_rca12_fa66_y2 = f_u_wallace_rca12_fa66_y0 ^ f_u_wallace_rca12_fa66_f_u_wallace_rca12_and_2_11_y0;
  assign f_u_wallace_rca12_fa66_y3 = f_u_wallace_rca12_fa66_y0 & f_u_wallace_rca12_fa66_f_u_wallace_rca12_and_2_11_y0;
  assign f_u_wallace_rca12_fa66_y4 = f_u_wallace_rca12_fa66_y1 | f_u_wallace_rca12_fa66_y3;
  assign f_u_wallace_rca12_and_3_11_a_3 = a_3;
  assign f_u_wallace_rca12_and_3_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_3_11_y0 = f_u_wallace_rca12_and_3_11_a_3 & f_u_wallace_rca12_and_3_11_b_11;
  assign f_u_wallace_rca12_fa67_f_u_wallace_rca12_fa66_y4 = f_u_wallace_rca12_fa66_y4;
  assign f_u_wallace_rca12_fa67_f_u_wallace_rca12_and_3_11_y0 = f_u_wallace_rca12_and_3_11_y0;
  assign f_u_wallace_rca12_fa67_f_u_wallace_rca12_fa11_y2 = f_u_wallace_rca12_fa11_y2;
  assign f_u_wallace_rca12_fa67_y0 = f_u_wallace_rca12_fa67_f_u_wallace_rca12_fa66_y4 ^ f_u_wallace_rca12_fa67_f_u_wallace_rca12_and_3_11_y0;
  assign f_u_wallace_rca12_fa67_y1 = f_u_wallace_rca12_fa67_f_u_wallace_rca12_fa66_y4 & f_u_wallace_rca12_fa67_f_u_wallace_rca12_and_3_11_y0;
  assign f_u_wallace_rca12_fa67_y2 = f_u_wallace_rca12_fa67_y0 ^ f_u_wallace_rca12_fa67_f_u_wallace_rca12_fa11_y2;
  assign f_u_wallace_rca12_fa67_y3 = f_u_wallace_rca12_fa67_y0 & f_u_wallace_rca12_fa67_f_u_wallace_rca12_fa11_y2;
  assign f_u_wallace_rca12_fa67_y4 = f_u_wallace_rca12_fa67_y1 | f_u_wallace_rca12_fa67_y3;
  assign f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa67_y4 = f_u_wallace_rca12_fa67_y4;
  assign f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa12_y2 = f_u_wallace_rca12_fa12_y2;
  assign f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa29_y2 = f_u_wallace_rca12_fa29_y2;
  assign f_u_wallace_rca12_fa68_y0 = f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa67_y4 ^ f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa12_y2;
  assign f_u_wallace_rca12_fa68_y1 = f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa67_y4 & f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa12_y2;
  assign f_u_wallace_rca12_fa68_y2 = f_u_wallace_rca12_fa68_y0 ^ f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa29_y2;
  assign f_u_wallace_rca12_fa68_y3 = f_u_wallace_rca12_fa68_y0 & f_u_wallace_rca12_fa68_f_u_wallace_rca12_fa29_y2;
  assign f_u_wallace_rca12_fa68_y4 = f_u_wallace_rca12_fa68_y1 | f_u_wallace_rca12_fa68_y3;
  assign f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa68_y4 = f_u_wallace_rca12_fa68_y4;
  assign f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa30_y2 = f_u_wallace_rca12_fa30_y2;
  assign f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa45_y2 = f_u_wallace_rca12_fa45_y2;
  assign f_u_wallace_rca12_fa69_y0 = f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa68_y4 ^ f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa30_y2;
  assign f_u_wallace_rca12_fa69_y1 = f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa68_y4 & f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa30_y2;
  assign f_u_wallace_rca12_fa69_y2 = f_u_wallace_rca12_fa69_y0 ^ f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa45_y2;
  assign f_u_wallace_rca12_fa69_y3 = f_u_wallace_rca12_fa69_y0 & f_u_wallace_rca12_fa69_f_u_wallace_rca12_fa45_y2;
  assign f_u_wallace_rca12_fa69_y4 = f_u_wallace_rca12_fa69_y1 | f_u_wallace_rca12_fa69_y3;
  assign f_u_wallace_rca12_ha5_f_u_wallace_rca12_fa36_y2 = f_u_wallace_rca12_fa36_y2;
  assign f_u_wallace_rca12_ha5_f_u_wallace_rca12_fa49_y2 = f_u_wallace_rca12_fa49_y2;
  assign f_u_wallace_rca12_ha5_y0 = f_u_wallace_rca12_ha5_f_u_wallace_rca12_fa36_y2 ^ f_u_wallace_rca12_ha5_f_u_wallace_rca12_fa49_y2;
  assign f_u_wallace_rca12_ha5_y1 = f_u_wallace_rca12_ha5_f_u_wallace_rca12_fa36_y2 & f_u_wallace_rca12_ha5_f_u_wallace_rca12_fa49_y2;
  assign f_u_wallace_rca12_fa70_f_u_wallace_rca12_ha5_y1 = f_u_wallace_rca12_ha5_y1;
  assign f_u_wallace_rca12_fa70_f_u_wallace_rca12_fa22_y2 = f_u_wallace_rca12_fa22_y2;
  assign f_u_wallace_rca12_fa70_f_u_wallace_rca12_fa37_y2 = f_u_wallace_rca12_fa37_y2;
  assign f_u_wallace_rca12_fa70_y0 = f_u_wallace_rca12_fa70_f_u_wallace_rca12_ha5_y1 ^ f_u_wallace_rca12_fa70_f_u_wallace_rca12_fa22_y2;
  assign f_u_wallace_rca12_fa70_y1 = f_u_wallace_rca12_fa70_f_u_wallace_rca12_ha5_y1 & f_u_wallace_rca12_fa70_f_u_wallace_rca12_fa22_y2;
  assign f_u_wallace_rca12_fa70_y2 = f_u_wallace_rca12_fa70_y0 ^ f_u_wallace_rca12_fa70_f_u_wallace_rca12_fa37_y2;
  assign f_u_wallace_rca12_fa70_y3 = f_u_wallace_rca12_fa70_y0 & f_u_wallace_rca12_fa70_f_u_wallace_rca12_fa37_y2;
  assign f_u_wallace_rca12_fa70_y4 = f_u_wallace_rca12_fa70_y1 | f_u_wallace_rca12_fa70_y3;
  assign f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa70_y4 = f_u_wallace_rca12_fa70_y4;
  assign f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa6_y2 = f_u_wallace_rca12_fa6_y2;
  assign f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa23_y2 = f_u_wallace_rca12_fa23_y2;
  assign f_u_wallace_rca12_fa71_y0 = f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa70_y4 ^ f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa6_y2;
  assign f_u_wallace_rca12_fa71_y1 = f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa70_y4 & f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa6_y2;
  assign f_u_wallace_rca12_fa71_y2 = f_u_wallace_rca12_fa71_y0 ^ f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa23_y2;
  assign f_u_wallace_rca12_fa71_y3 = f_u_wallace_rca12_fa71_y0 & f_u_wallace_rca12_fa71_f_u_wallace_rca12_fa23_y2;
  assign f_u_wallace_rca12_fa71_y4 = f_u_wallace_rca12_fa71_y1 | f_u_wallace_rca12_fa71_y3;
  assign f_u_wallace_rca12_and_0_10_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_0_10_y0 = f_u_wallace_rca12_and_0_10_a_0 & f_u_wallace_rca12_and_0_10_b_10;
  assign f_u_wallace_rca12_fa72_f_u_wallace_rca12_fa71_y4 = f_u_wallace_rca12_fa71_y4;
  assign f_u_wallace_rca12_fa72_f_u_wallace_rca12_and_0_10_y0 = f_u_wallace_rca12_and_0_10_y0;
  assign f_u_wallace_rca12_fa72_f_u_wallace_rca12_fa7_y2 = f_u_wallace_rca12_fa7_y2;
  assign f_u_wallace_rca12_fa72_y0 = f_u_wallace_rca12_fa72_f_u_wallace_rca12_fa71_y4 ^ f_u_wallace_rca12_fa72_f_u_wallace_rca12_and_0_10_y0;
  assign f_u_wallace_rca12_fa72_y1 = f_u_wallace_rca12_fa72_f_u_wallace_rca12_fa71_y4 & f_u_wallace_rca12_fa72_f_u_wallace_rca12_and_0_10_y0;
  assign f_u_wallace_rca12_fa72_y2 = f_u_wallace_rca12_fa72_y0 ^ f_u_wallace_rca12_fa72_f_u_wallace_rca12_fa7_y2;
  assign f_u_wallace_rca12_fa72_y3 = f_u_wallace_rca12_fa72_y0 & f_u_wallace_rca12_fa72_f_u_wallace_rca12_fa7_y2;
  assign f_u_wallace_rca12_fa72_y4 = f_u_wallace_rca12_fa72_y1 | f_u_wallace_rca12_fa72_y3;
  assign f_u_wallace_rca12_and_1_10_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_1_10_y0 = f_u_wallace_rca12_and_1_10_a_1 & f_u_wallace_rca12_and_1_10_b_10;
  assign f_u_wallace_rca12_and_0_11_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_0_11_y0 = f_u_wallace_rca12_and_0_11_a_0 & f_u_wallace_rca12_and_0_11_b_11;
  assign f_u_wallace_rca12_fa73_f_u_wallace_rca12_fa72_y4 = f_u_wallace_rca12_fa72_y4;
  assign f_u_wallace_rca12_fa73_f_u_wallace_rca12_and_1_10_y0 = f_u_wallace_rca12_and_1_10_y0;
  assign f_u_wallace_rca12_fa73_f_u_wallace_rca12_and_0_11_y0 = f_u_wallace_rca12_and_0_11_y0;
  assign f_u_wallace_rca12_fa73_y0 = f_u_wallace_rca12_fa73_f_u_wallace_rca12_fa72_y4 ^ f_u_wallace_rca12_fa73_f_u_wallace_rca12_and_1_10_y0;
  assign f_u_wallace_rca12_fa73_y1 = f_u_wallace_rca12_fa73_f_u_wallace_rca12_fa72_y4 & f_u_wallace_rca12_fa73_f_u_wallace_rca12_and_1_10_y0;
  assign f_u_wallace_rca12_fa73_y2 = f_u_wallace_rca12_fa73_y0 ^ f_u_wallace_rca12_fa73_f_u_wallace_rca12_and_0_11_y0;
  assign f_u_wallace_rca12_fa73_y3 = f_u_wallace_rca12_fa73_y0 & f_u_wallace_rca12_fa73_f_u_wallace_rca12_and_0_11_y0;
  assign f_u_wallace_rca12_fa73_y4 = f_u_wallace_rca12_fa73_y1 | f_u_wallace_rca12_fa73_y3;
  assign f_u_wallace_rca12_and_1_11_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_1_11_y0 = f_u_wallace_rca12_and_1_11_a_1 & f_u_wallace_rca12_and_1_11_b_11;
  assign f_u_wallace_rca12_fa74_f_u_wallace_rca12_fa73_y4 = f_u_wallace_rca12_fa73_y4;
  assign f_u_wallace_rca12_fa74_f_u_wallace_rca12_and_1_11_y0 = f_u_wallace_rca12_and_1_11_y0;
  assign f_u_wallace_rca12_fa74_f_u_wallace_rca12_fa9_y2 = f_u_wallace_rca12_fa9_y2;
  assign f_u_wallace_rca12_fa74_y0 = f_u_wallace_rca12_fa74_f_u_wallace_rca12_fa73_y4 ^ f_u_wallace_rca12_fa74_f_u_wallace_rca12_and_1_11_y0;
  assign f_u_wallace_rca12_fa74_y1 = f_u_wallace_rca12_fa74_f_u_wallace_rca12_fa73_y4 & f_u_wallace_rca12_fa74_f_u_wallace_rca12_and_1_11_y0;
  assign f_u_wallace_rca12_fa74_y2 = f_u_wallace_rca12_fa74_y0 ^ f_u_wallace_rca12_fa74_f_u_wallace_rca12_fa9_y2;
  assign f_u_wallace_rca12_fa74_y3 = f_u_wallace_rca12_fa74_y0 & f_u_wallace_rca12_fa74_f_u_wallace_rca12_fa9_y2;
  assign f_u_wallace_rca12_fa74_y4 = f_u_wallace_rca12_fa74_y1 | f_u_wallace_rca12_fa74_y3;
  assign f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa74_y4 = f_u_wallace_rca12_fa74_y4;
  assign f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa10_y2 = f_u_wallace_rca12_fa10_y2;
  assign f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa27_y2 = f_u_wallace_rca12_fa27_y2;
  assign f_u_wallace_rca12_fa75_y0 = f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa74_y4 ^ f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa10_y2;
  assign f_u_wallace_rca12_fa75_y1 = f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa74_y4 & f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa10_y2;
  assign f_u_wallace_rca12_fa75_y2 = f_u_wallace_rca12_fa75_y0 ^ f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa27_y2;
  assign f_u_wallace_rca12_fa75_y3 = f_u_wallace_rca12_fa75_y0 & f_u_wallace_rca12_fa75_f_u_wallace_rca12_fa27_y2;
  assign f_u_wallace_rca12_fa75_y4 = f_u_wallace_rca12_fa75_y1 | f_u_wallace_rca12_fa75_y3;
  assign f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa75_y4 = f_u_wallace_rca12_fa75_y4;
  assign f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa28_y2 = f_u_wallace_rca12_fa28_y2;
  assign f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa43_y2 = f_u_wallace_rca12_fa43_y2;
  assign f_u_wallace_rca12_fa76_y0 = f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa75_y4 ^ f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa28_y2;
  assign f_u_wallace_rca12_fa76_y1 = f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa75_y4 & f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa28_y2;
  assign f_u_wallace_rca12_fa76_y2 = f_u_wallace_rca12_fa76_y0 ^ f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa43_y2;
  assign f_u_wallace_rca12_fa76_y3 = f_u_wallace_rca12_fa76_y0 & f_u_wallace_rca12_fa76_f_u_wallace_rca12_fa43_y2;
  assign f_u_wallace_rca12_fa76_y4 = f_u_wallace_rca12_fa76_y1 | f_u_wallace_rca12_fa76_y3;
  assign f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa76_y4 = f_u_wallace_rca12_fa76_y4;
  assign f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa44_y2 = f_u_wallace_rca12_fa44_y2;
  assign f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa57_y2 = f_u_wallace_rca12_fa57_y2;
  assign f_u_wallace_rca12_fa77_y0 = f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa76_y4 ^ f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa44_y2;
  assign f_u_wallace_rca12_fa77_y1 = f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa76_y4 & f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa44_y2;
  assign f_u_wallace_rca12_fa77_y2 = f_u_wallace_rca12_fa77_y0 ^ f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa57_y2;
  assign f_u_wallace_rca12_fa77_y3 = f_u_wallace_rca12_fa77_y0 & f_u_wallace_rca12_fa77_f_u_wallace_rca12_fa57_y2;
  assign f_u_wallace_rca12_fa77_y4 = f_u_wallace_rca12_fa77_y1 | f_u_wallace_rca12_fa77_y3;
  assign f_u_wallace_rca12_ha6_f_u_wallace_rca12_fa50_y2 = f_u_wallace_rca12_fa50_y2;
  assign f_u_wallace_rca12_ha6_f_u_wallace_rca12_fa61_y2 = f_u_wallace_rca12_fa61_y2;
  assign f_u_wallace_rca12_ha6_y0 = f_u_wallace_rca12_ha6_f_u_wallace_rca12_fa50_y2 ^ f_u_wallace_rca12_ha6_f_u_wallace_rca12_fa61_y2;
  assign f_u_wallace_rca12_ha6_y1 = f_u_wallace_rca12_ha6_f_u_wallace_rca12_fa50_y2 & f_u_wallace_rca12_ha6_f_u_wallace_rca12_fa61_y2;
  assign f_u_wallace_rca12_fa78_f_u_wallace_rca12_ha6_y1 = f_u_wallace_rca12_ha6_y1;
  assign f_u_wallace_rca12_fa78_f_u_wallace_rca12_fa38_y2 = f_u_wallace_rca12_fa38_y2;
  assign f_u_wallace_rca12_fa78_f_u_wallace_rca12_fa51_y2 = f_u_wallace_rca12_fa51_y2;
  assign f_u_wallace_rca12_fa78_y0 = f_u_wallace_rca12_fa78_f_u_wallace_rca12_ha6_y1 ^ f_u_wallace_rca12_fa78_f_u_wallace_rca12_fa38_y2;
  assign f_u_wallace_rca12_fa78_y1 = f_u_wallace_rca12_fa78_f_u_wallace_rca12_ha6_y1 & f_u_wallace_rca12_fa78_f_u_wallace_rca12_fa38_y2;
  assign f_u_wallace_rca12_fa78_y2 = f_u_wallace_rca12_fa78_y0 ^ f_u_wallace_rca12_fa78_f_u_wallace_rca12_fa51_y2;
  assign f_u_wallace_rca12_fa78_y3 = f_u_wallace_rca12_fa78_y0 & f_u_wallace_rca12_fa78_f_u_wallace_rca12_fa51_y2;
  assign f_u_wallace_rca12_fa78_y4 = f_u_wallace_rca12_fa78_y1 | f_u_wallace_rca12_fa78_y3;
  assign f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa78_y4 = f_u_wallace_rca12_fa78_y4;
  assign f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa24_y2 = f_u_wallace_rca12_fa24_y2;
  assign f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa39_y2 = f_u_wallace_rca12_fa39_y2;
  assign f_u_wallace_rca12_fa79_y0 = f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa78_y4 ^ f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa24_y2;
  assign f_u_wallace_rca12_fa79_y1 = f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa78_y4 & f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa24_y2;
  assign f_u_wallace_rca12_fa79_y2 = f_u_wallace_rca12_fa79_y0 ^ f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa39_y2;
  assign f_u_wallace_rca12_fa79_y3 = f_u_wallace_rca12_fa79_y0 & f_u_wallace_rca12_fa79_f_u_wallace_rca12_fa39_y2;
  assign f_u_wallace_rca12_fa79_y4 = f_u_wallace_rca12_fa79_y1 | f_u_wallace_rca12_fa79_y3;
  assign f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa79_y4 = f_u_wallace_rca12_fa79_y4;
  assign f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa8_y2 = f_u_wallace_rca12_fa8_y2;
  assign f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa25_y2 = f_u_wallace_rca12_fa25_y2;
  assign f_u_wallace_rca12_fa80_y0 = f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa79_y4 ^ f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa8_y2;
  assign f_u_wallace_rca12_fa80_y1 = f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa79_y4 & f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa8_y2;
  assign f_u_wallace_rca12_fa80_y2 = f_u_wallace_rca12_fa80_y0 ^ f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa25_y2;
  assign f_u_wallace_rca12_fa80_y3 = f_u_wallace_rca12_fa80_y0 & f_u_wallace_rca12_fa80_f_u_wallace_rca12_fa25_y2;
  assign f_u_wallace_rca12_fa80_y4 = f_u_wallace_rca12_fa80_y1 | f_u_wallace_rca12_fa80_y3;
  assign f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa80_y4 = f_u_wallace_rca12_fa80_y4;
  assign f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa26_y2 = f_u_wallace_rca12_fa26_y2;
  assign f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa41_y2 = f_u_wallace_rca12_fa41_y2;
  assign f_u_wallace_rca12_fa81_y0 = f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa80_y4 ^ f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa26_y2;
  assign f_u_wallace_rca12_fa81_y1 = f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa80_y4 & f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa26_y2;
  assign f_u_wallace_rca12_fa81_y2 = f_u_wallace_rca12_fa81_y0 ^ f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa41_y2;
  assign f_u_wallace_rca12_fa81_y3 = f_u_wallace_rca12_fa81_y0 & f_u_wallace_rca12_fa81_f_u_wallace_rca12_fa41_y2;
  assign f_u_wallace_rca12_fa81_y4 = f_u_wallace_rca12_fa81_y1 | f_u_wallace_rca12_fa81_y3;
  assign f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa81_y4 = f_u_wallace_rca12_fa81_y4;
  assign f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa42_y2 = f_u_wallace_rca12_fa42_y2;
  assign f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa55_y2 = f_u_wallace_rca12_fa55_y2;
  assign f_u_wallace_rca12_fa82_y0 = f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa81_y4 ^ f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa42_y2;
  assign f_u_wallace_rca12_fa82_y1 = f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa81_y4 & f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa42_y2;
  assign f_u_wallace_rca12_fa82_y2 = f_u_wallace_rca12_fa82_y0 ^ f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa55_y2;
  assign f_u_wallace_rca12_fa82_y3 = f_u_wallace_rca12_fa82_y0 & f_u_wallace_rca12_fa82_f_u_wallace_rca12_fa55_y2;
  assign f_u_wallace_rca12_fa82_y4 = f_u_wallace_rca12_fa82_y1 | f_u_wallace_rca12_fa82_y3;
  assign f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa82_y4 = f_u_wallace_rca12_fa82_y4;
  assign f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa56_y2 = f_u_wallace_rca12_fa56_y2;
  assign f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa67_y2 = f_u_wallace_rca12_fa67_y2;
  assign f_u_wallace_rca12_fa83_y0 = f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa82_y4 ^ f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa56_y2;
  assign f_u_wallace_rca12_fa83_y1 = f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa82_y4 & f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa56_y2;
  assign f_u_wallace_rca12_fa83_y2 = f_u_wallace_rca12_fa83_y0 ^ f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa67_y2;
  assign f_u_wallace_rca12_fa83_y3 = f_u_wallace_rca12_fa83_y0 & f_u_wallace_rca12_fa83_f_u_wallace_rca12_fa67_y2;
  assign f_u_wallace_rca12_fa83_y4 = f_u_wallace_rca12_fa83_y1 | f_u_wallace_rca12_fa83_y3;
  assign f_u_wallace_rca12_ha7_f_u_wallace_rca12_fa62_y2 = f_u_wallace_rca12_fa62_y2;
  assign f_u_wallace_rca12_ha7_f_u_wallace_rca12_fa71_y2 = f_u_wallace_rca12_fa71_y2;
  assign f_u_wallace_rca12_ha7_y0 = f_u_wallace_rca12_ha7_f_u_wallace_rca12_fa62_y2 ^ f_u_wallace_rca12_ha7_f_u_wallace_rca12_fa71_y2;
  assign f_u_wallace_rca12_ha7_y1 = f_u_wallace_rca12_ha7_f_u_wallace_rca12_fa62_y2 & f_u_wallace_rca12_ha7_f_u_wallace_rca12_fa71_y2;
  assign f_u_wallace_rca12_fa84_f_u_wallace_rca12_ha7_y1 = f_u_wallace_rca12_ha7_y1;
  assign f_u_wallace_rca12_fa84_f_u_wallace_rca12_fa52_y2 = f_u_wallace_rca12_fa52_y2;
  assign f_u_wallace_rca12_fa84_f_u_wallace_rca12_fa63_y2 = f_u_wallace_rca12_fa63_y2;
  assign f_u_wallace_rca12_fa84_y0 = f_u_wallace_rca12_fa84_f_u_wallace_rca12_ha7_y1 ^ f_u_wallace_rca12_fa84_f_u_wallace_rca12_fa52_y2;
  assign f_u_wallace_rca12_fa84_y1 = f_u_wallace_rca12_fa84_f_u_wallace_rca12_ha7_y1 & f_u_wallace_rca12_fa84_f_u_wallace_rca12_fa52_y2;
  assign f_u_wallace_rca12_fa84_y2 = f_u_wallace_rca12_fa84_y0 ^ f_u_wallace_rca12_fa84_f_u_wallace_rca12_fa63_y2;
  assign f_u_wallace_rca12_fa84_y3 = f_u_wallace_rca12_fa84_y0 & f_u_wallace_rca12_fa84_f_u_wallace_rca12_fa63_y2;
  assign f_u_wallace_rca12_fa84_y4 = f_u_wallace_rca12_fa84_y1 | f_u_wallace_rca12_fa84_y3;
  assign f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa84_y4 = f_u_wallace_rca12_fa84_y4;
  assign f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa40_y2 = f_u_wallace_rca12_fa40_y2;
  assign f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa53_y2 = f_u_wallace_rca12_fa53_y2;
  assign f_u_wallace_rca12_fa85_y0 = f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa84_y4 ^ f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa40_y2;
  assign f_u_wallace_rca12_fa85_y1 = f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa84_y4 & f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa40_y2;
  assign f_u_wallace_rca12_fa85_y2 = f_u_wallace_rca12_fa85_y0 ^ f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa53_y2;
  assign f_u_wallace_rca12_fa85_y3 = f_u_wallace_rca12_fa85_y0 & f_u_wallace_rca12_fa85_f_u_wallace_rca12_fa53_y2;
  assign f_u_wallace_rca12_fa85_y4 = f_u_wallace_rca12_fa85_y1 | f_u_wallace_rca12_fa85_y3;
  assign f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa85_y4 = f_u_wallace_rca12_fa85_y4;
  assign f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa54_y2 = f_u_wallace_rca12_fa54_y2;
  assign f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa65_y2 = f_u_wallace_rca12_fa65_y2;
  assign f_u_wallace_rca12_fa86_y0 = f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa85_y4 ^ f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa54_y2;
  assign f_u_wallace_rca12_fa86_y1 = f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa85_y4 & f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa54_y2;
  assign f_u_wallace_rca12_fa86_y2 = f_u_wallace_rca12_fa86_y0 ^ f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa65_y2;
  assign f_u_wallace_rca12_fa86_y3 = f_u_wallace_rca12_fa86_y0 & f_u_wallace_rca12_fa86_f_u_wallace_rca12_fa65_y2;
  assign f_u_wallace_rca12_fa86_y4 = f_u_wallace_rca12_fa86_y1 | f_u_wallace_rca12_fa86_y3;
  assign f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa86_y4 = f_u_wallace_rca12_fa86_y4;
  assign f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa66_y2 = f_u_wallace_rca12_fa66_y2;
  assign f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa75_y2 = f_u_wallace_rca12_fa75_y2;
  assign f_u_wallace_rca12_fa87_y0 = f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa86_y4 ^ f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa66_y2;
  assign f_u_wallace_rca12_fa87_y1 = f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa86_y4 & f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa66_y2;
  assign f_u_wallace_rca12_fa87_y2 = f_u_wallace_rca12_fa87_y0 ^ f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa75_y2;
  assign f_u_wallace_rca12_fa87_y3 = f_u_wallace_rca12_fa87_y0 & f_u_wallace_rca12_fa87_f_u_wallace_rca12_fa75_y2;
  assign f_u_wallace_rca12_fa87_y4 = f_u_wallace_rca12_fa87_y1 | f_u_wallace_rca12_fa87_y3;
  assign f_u_wallace_rca12_ha8_f_u_wallace_rca12_fa72_y2 = f_u_wallace_rca12_fa72_y2;
  assign f_u_wallace_rca12_ha8_f_u_wallace_rca12_fa79_y2 = f_u_wallace_rca12_fa79_y2;
  assign f_u_wallace_rca12_ha8_y0 = f_u_wallace_rca12_ha8_f_u_wallace_rca12_fa72_y2 ^ f_u_wallace_rca12_ha8_f_u_wallace_rca12_fa79_y2;
  assign f_u_wallace_rca12_ha8_y1 = f_u_wallace_rca12_ha8_f_u_wallace_rca12_fa72_y2 & f_u_wallace_rca12_ha8_f_u_wallace_rca12_fa79_y2;
  assign f_u_wallace_rca12_fa88_f_u_wallace_rca12_ha8_y1 = f_u_wallace_rca12_ha8_y1;
  assign f_u_wallace_rca12_fa88_f_u_wallace_rca12_fa64_y2 = f_u_wallace_rca12_fa64_y2;
  assign f_u_wallace_rca12_fa88_f_u_wallace_rca12_fa73_y2 = f_u_wallace_rca12_fa73_y2;
  assign f_u_wallace_rca12_fa88_y0 = f_u_wallace_rca12_fa88_f_u_wallace_rca12_ha8_y1 ^ f_u_wallace_rca12_fa88_f_u_wallace_rca12_fa64_y2;
  assign f_u_wallace_rca12_fa88_y1 = f_u_wallace_rca12_fa88_f_u_wallace_rca12_ha8_y1 & f_u_wallace_rca12_fa88_f_u_wallace_rca12_fa64_y2;
  assign f_u_wallace_rca12_fa88_y2 = f_u_wallace_rca12_fa88_y0 ^ f_u_wallace_rca12_fa88_f_u_wallace_rca12_fa73_y2;
  assign f_u_wallace_rca12_fa88_y3 = f_u_wallace_rca12_fa88_y0 & f_u_wallace_rca12_fa88_f_u_wallace_rca12_fa73_y2;
  assign f_u_wallace_rca12_fa88_y4 = f_u_wallace_rca12_fa88_y1 | f_u_wallace_rca12_fa88_y3;
  assign f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa88_y4 = f_u_wallace_rca12_fa88_y4;
  assign f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa74_y2 = f_u_wallace_rca12_fa74_y2;
  assign f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa81_y2 = f_u_wallace_rca12_fa81_y2;
  assign f_u_wallace_rca12_fa89_y0 = f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa88_y4 ^ f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa74_y2;
  assign f_u_wallace_rca12_fa89_y1 = f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa88_y4 & f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa74_y2;
  assign f_u_wallace_rca12_fa89_y2 = f_u_wallace_rca12_fa89_y0 ^ f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa81_y2;
  assign f_u_wallace_rca12_fa89_y3 = f_u_wallace_rca12_fa89_y0 & f_u_wallace_rca12_fa89_f_u_wallace_rca12_fa81_y2;
  assign f_u_wallace_rca12_fa89_y4 = f_u_wallace_rca12_fa89_y1 | f_u_wallace_rca12_fa89_y3;
  assign f_u_wallace_rca12_ha9_f_u_wallace_rca12_fa80_y2 = f_u_wallace_rca12_fa80_y2;
  assign f_u_wallace_rca12_ha9_f_u_wallace_rca12_fa85_y2 = f_u_wallace_rca12_fa85_y2;
  assign f_u_wallace_rca12_ha9_y0 = f_u_wallace_rca12_ha9_f_u_wallace_rca12_fa80_y2 ^ f_u_wallace_rca12_ha9_f_u_wallace_rca12_fa85_y2;
  assign f_u_wallace_rca12_ha9_y1 = f_u_wallace_rca12_ha9_f_u_wallace_rca12_fa80_y2 & f_u_wallace_rca12_ha9_f_u_wallace_rca12_fa85_y2;
  assign f_u_wallace_rca12_ha10_f_u_wallace_rca12_ha9_y1 = f_u_wallace_rca12_ha9_y1;
  assign f_u_wallace_rca12_ha10_f_u_wallace_rca12_fa86_y2 = f_u_wallace_rca12_fa86_y2;
  assign f_u_wallace_rca12_ha10_y0 = f_u_wallace_rca12_ha10_f_u_wallace_rca12_ha9_y1 ^ f_u_wallace_rca12_ha10_f_u_wallace_rca12_fa86_y2;
  assign f_u_wallace_rca12_ha10_y1 = f_u_wallace_rca12_ha10_f_u_wallace_rca12_ha9_y1 & f_u_wallace_rca12_ha10_f_u_wallace_rca12_fa86_y2;
  assign f_u_wallace_rca12_fa90_f_u_wallace_rca12_ha10_y1 = f_u_wallace_rca12_ha10_y1;
  assign f_u_wallace_rca12_fa90_f_u_wallace_rca12_fa89_y4 = f_u_wallace_rca12_fa89_y4;
  assign f_u_wallace_rca12_fa90_f_u_wallace_rca12_fa82_y2 = f_u_wallace_rca12_fa82_y2;
  assign f_u_wallace_rca12_fa90_y0 = f_u_wallace_rca12_fa90_f_u_wallace_rca12_ha10_y1 ^ f_u_wallace_rca12_fa90_f_u_wallace_rca12_fa89_y4;
  assign f_u_wallace_rca12_fa90_y1 = f_u_wallace_rca12_fa90_f_u_wallace_rca12_ha10_y1 & f_u_wallace_rca12_fa90_f_u_wallace_rca12_fa89_y4;
  assign f_u_wallace_rca12_fa90_y2 = f_u_wallace_rca12_fa90_y0 ^ f_u_wallace_rca12_fa90_f_u_wallace_rca12_fa82_y2;
  assign f_u_wallace_rca12_fa90_y3 = f_u_wallace_rca12_fa90_y0 & f_u_wallace_rca12_fa90_f_u_wallace_rca12_fa82_y2;
  assign f_u_wallace_rca12_fa90_y4 = f_u_wallace_rca12_fa90_y1 | f_u_wallace_rca12_fa90_y3;
  assign f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa90_y4 = f_u_wallace_rca12_fa90_y4;
  assign f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa87_y4 = f_u_wallace_rca12_fa87_y4;
  assign f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa76_y2 = f_u_wallace_rca12_fa76_y2;
  assign f_u_wallace_rca12_fa91_y0 = f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa90_y4 ^ f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa87_y4;
  assign f_u_wallace_rca12_fa91_y1 = f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa90_y4 & f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa87_y4;
  assign f_u_wallace_rca12_fa91_y2 = f_u_wallace_rca12_fa91_y0 ^ f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa76_y2;
  assign f_u_wallace_rca12_fa91_y3 = f_u_wallace_rca12_fa91_y0 & f_u_wallace_rca12_fa91_f_u_wallace_rca12_fa76_y2;
  assign f_u_wallace_rca12_fa91_y4 = f_u_wallace_rca12_fa91_y1 | f_u_wallace_rca12_fa91_y3;
  assign f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa91_y4 = f_u_wallace_rca12_fa91_y4;
  assign f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa83_y4 = f_u_wallace_rca12_fa83_y4;
  assign f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa68_y2 = f_u_wallace_rca12_fa68_y2;
  assign f_u_wallace_rca12_fa92_y0 = f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa91_y4 ^ f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa83_y4;
  assign f_u_wallace_rca12_fa92_y1 = f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa91_y4 & f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa83_y4;
  assign f_u_wallace_rca12_fa92_y2 = f_u_wallace_rca12_fa92_y0 ^ f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa68_y2;
  assign f_u_wallace_rca12_fa92_y3 = f_u_wallace_rca12_fa92_y0 & f_u_wallace_rca12_fa92_f_u_wallace_rca12_fa68_y2;
  assign f_u_wallace_rca12_fa92_y4 = f_u_wallace_rca12_fa92_y1 | f_u_wallace_rca12_fa92_y3;
  assign f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa92_y4 = f_u_wallace_rca12_fa92_y4;
  assign f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa77_y4 = f_u_wallace_rca12_fa77_y4;
  assign f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa58_y2 = f_u_wallace_rca12_fa58_y2;
  assign f_u_wallace_rca12_fa93_y0 = f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa92_y4 ^ f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa77_y4;
  assign f_u_wallace_rca12_fa93_y1 = f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa92_y4 & f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa77_y4;
  assign f_u_wallace_rca12_fa93_y2 = f_u_wallace_rca12_fa93_y0 ^ f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa58_y2;
  assign f_u_wallace_rca12_fa93_y3 = f_u_wallace_rca12_fa93_y0 & f_u_wallace_rca12_fa93_f_u_wallace_rca12_fa58_y2;
  assign f_u_wallace_rca12_fa93_y4 = f_u_wallace_rca12_fa93_y1 | f_u_wallace_rca12_fa93_y3;
  assign f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa93_y4 = f_u_wallace_rca12_fa93_y4;
  assign f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa69_y4 = f_u_wallace_rca12_fa69_y4;
  assign f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa46_y2 = f_u_wallace_rca12_fa46_y2;
  assign f_u_wallace_rca12_fa94_y0 = f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa93_y4 ^ f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa69_y4;
  assign f_u_wallace_rca12_fa94_y1 = f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa93_y4 & f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa69_y4;
  assign f_u_wallace_rca12_fa94_y2 = f_u_wallace_rca12_fa94_y0 ^ f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa46_y2;
  assign f_u_wallace_rca12_fa94_y3 = f_u_wallace_rca12_fa94_y0 & f_u_wallace_rca12_fa94_f_u_wallace_rca12_fa46_y2;
  assign f_u_wallace_rca12_fa94_y4 = f_u_wallace_rca12_fa94_y1 | f_u_wallace_rca12_fa94_y3;
  assign f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa94_y4 = f_u_wallace_rca12_fa94_y4;
  assign f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa59_y4 = f_u_wallace_rca12_fa59_y4;
  assign f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa32_y2 = f_u_wallace_rca12_fa32_y2;
  assign f_u_wallace_rca12_fa95_y0 = f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa94_y4 ^ f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa59_y4;
  assign f_u_wallace_rca12_fa95_y1 = f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa94_y4 & f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa59_y4;
  assign f_u_wallace_rca12_fa95_y2 = f_u_wallace_rca12_fa95_y0 ^ f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa32_y2;
  assign f_u_wallace_rca12_fa95_y3 = f_u_wallace_rca12_fa95_y0 & f_u_wallace_rca12_fa95_f_u_wallace_rca12_fa32_y2;
  assign f_u_wallace_rca12_fa95_y4 = f_u_wallace_rca12_fa95_y1 | f_u_wallace_rca12_fa95_y3;
  assign f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa95_y4 = f_u_wallace_rca12_fa95_y4;
  assign f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa47_y4 = f_u_wallace_rca12_fa47_y4;
  assign f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa16_y2 = f_u_wallace_rca12_fa16_y2;
  assign f_u_wallace_rca12_fa96_y0 = f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa95_y4 ^ f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa47_y4;
  assign f_u_wallace_rca12_fa96_y1 = f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa95_y4 & f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa47_y4;
  assign f_u_wallace_rca12_fa96_y2 = f_u_wallace_rca12_fa96_y0 ^ f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa16_y2;
  assign f_u_wallace_rca12_fa96_y3 = f_u_wallace_rca12_fa96_y0 & f_u_wallace_rca12_fa96_f_u_wallace_rca12_fa16_y2;
  assign f_u_wallace_rca12_fa96_y4 = f_u_wallace_rca12_fa96_y1 | f_u_wallace_rca12_fa96_y3;
  assign f_u_wallace_rca12_and_9_11_a_9 = a_9;
  assign f_u_wallace_rca12_and_9_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_9_11_y0 = f_u_wallace_rca12_and_9_11_a_9 & f_u_wallace_rca12_and_9_11_b_11;
  assign f_u_wallace_rca12_fa97_f_u_wallace_rca12_fa96_y4 = f_u_wallace_rca12_fa96_y4;
  assign f_u_wallace_rca12_fa97_f_u_wallace_rca12_fa33_y4 = f_u_wallace_rca12_fa33_y4;
  assign f_u_wallace_rca12_fa97_f_u_wallace_rca12_and_9_11_y0 = f_u_wallace_rca12_and_9_11_y0;
  assign f_u_wallace_rca12_fa97_y0 = f_u_wallace_rca12_fa97_f_u_wallace_rca12_fa96_y4 ^ f_u_wallace_rca12_fa97_f_u_wallace_rca12_fa33_y4;
  assign f_u_wallace_rca12_fa97_y1 = f_u_wallace_rca12_fa97_f_u_wallace_rca12_fa96_y4 & f_u_wallace_rca12_fa97_f_u_wallace_rca12_fa33_y4;
  assign f_u_wallace_rca12_fa97_y2 = f_u_wallace_rca12_fa97_y0 ^ f_u_wallace_rca12_fa97_f_u_wallace_rca12_and_9_11_y0;
  assign f_u_wallace_rca12_fa97_y3 = f_u_wallace_rca12_fa97_y0 & f_u_wallace_rca12_fa97_f_u_wallace_rca12_and_9_11_y0;
  assign f_u_wallace_rca12_fa97_y4 = f_u_wallace_rca12_fa97_y1 | f_u_wallace_rca12_fa97_y3;
  assign f_u_wallace_rca12_and_11_10_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_10_b_10 = b_10;
  assign f_u_wallace_rca12_and_11_10_y0 = f_u_wallace_rca12_and_11_10_a_11 & f_u_wallace_rca12_and_11_10_b_10;
  assign f_u_wallace_rca12_fa98_f_u_wallace_rca12_fa97_y4 = f_u_wallace_rca12_fa97_y4;
  assign f_u_wallace_rca12_fa98_f_u_wallace_rca12_fa17_y4 = f_u_wallace_rca12_fa17_y4;
  assign f_u_wallace_rca12_fa98_f_u_wallace_rca12_and_11_10_y0 = f_u_wallace_rca12_and_11_10_y0;
  assign f_u_wallace_rca12_fa98_y0 = f_u_wallace_rca12_fa98_f_u_wallace_rca12_fa97_y4 ^ f_u_wallace_rca12_fa98_f_u_wallace_rca12_fa17_y4;
  assign f_u_wallace_rca12_fa98_y1 = f_u_wallace_rca12_fa98_f_u_wallace_rca12_fa97_y4 & f_u_wallace_rca12_fa98_f_u_wallace_rca12_fa17_y4;
  assign f_u_wallace_rca12_fa98_y2 = f_u_wallace_rca12_fa98_y0 ^ f_u_wallace_rca12_fa98_f_u_wallace_rca12_and_11_10_y0;
  assign f_u_wallace_rca12_fa98_y3 = f_u_wallace_rca12_fa98_y0 & f_u_wallace_rca12_fa98_f_u_wallace_rca12_and_11_10_y0;
  assign f_u_wallace_rca12_fa98_y4 = f_u_wallace_rca12_fa98_y1 | f_u_wallace_rca12_fa98_y3;
  assign f_u_wallace_rca12_and_0_0_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_0_0_y0 = f_u_wallace_rca12_and_0_0_a_0 & f_u_wallace_rca12_and_0_0_b_0;
  assign f_u_wallace_rca12_and_1_0_a_1 = a_1;
  assign f_u_wallace_rca12_and_1_0_b_0 = b_0;
  assign f_u_wallace_rca12_and_1_0_y0 = f_u_wallace_rca12_and_1_0_a_1 & f_u_wallace_rca12_and_1_0_b_0;
  assign f_u_wallace_rca12_and_0_2_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_2_b_2 = b_2;
  assign f_u_wallace_rca12_and_0_2_y0 = f_u_wallace_rca12_and_0_2_a_0 & f_u_wallace_rca12_and_0_2_b_2;
  assign f_u_wallace_rca12_and_10_11_a_10 = a_10;
  assign f_u_wallace_rca12_and_10_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_10_11_y0 = f_u_wallace_rca12_and_10_11_a_10 & f_u_wallace_rca12_and_10_11_b_11;
  assign f_u_wallace_rca12_and_0_1_a_0 = a_0;
  assign f_u_wallace_rca12_and_0_1_b_1 = b_1;
  assign f_u_wallace_rca12_and_0_1_y0 = f_u_wallace_rca12_and_0_1_a_0 & f_u_wallace_rca12_and_0_1_b_1;
  assign f_u_wallace_rca12_and_11_11_a_11 = a_11;
  assign f_u_wallace_rca12_and_11_11_b_11 = b_11;
  assign f_u_wallace_rca12_and_11_11_y0 = f_u_wallace_rca12_and_11_11_a_11 & f_u_wallace_rca12_and_11_11_b_11;
  assign f_u_wallace_rca12_u_rca22_ha_f_u_wallace_rca12_and_1_0_y0 = f_u_wallace_rca12_and_1_0_y0;
  assign f_u_wallace_rca12_u_rca22_ha_f_u_wallace_rca12_and_0_1_y0 = f_u_wallace_rca12_and_0_1_y0;
  assign f_u_wallace_rca12_u_rca22_ha_y0 = f_u_wallace_rca12_u_rca22_ha_f_u_wallace_rca12_and_1_0_y0 ^ f_u_wallace_rca12_u_rca22_ha_f_u_wallace_rca12_and_0_1_y0;
  assign f_u_wallace_rca12_u_rca22_ha_y1 = f_u_wallace_rca12_u_rca22_ha_f_u_wallace_rca12_and_1_0_y0 & f_u_wallace_rca12_u_rca22_ha_f_u_wallace_rca12_and_0_1_y0;
  assign f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_and_0_2_y0 = f_u_wallace_rca12_and_0_2_y0;
  assign f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_ha0_y0 = f_u_wallace_rca12_ha0_y0;
  assign f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_u_rca22_ha_y1 = f_u_wallace_rca12_u_rca22_ha_y1;
  assign f_u_wallace_rca12_u_rca22_fa1_y0 = f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_and_0_2_y0 ^ f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_ha0_y0;
  assign f_u_wallace_rca12_u_rca22_fa1_y1 = f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_and_0_2_y0 & f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_ha0_y0;
  assign f_u_wallace_rca12_u_rca22_fa1_y2 = f_u_wallace_rca12_u_rca22_fa1_y0 ^ f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_u_rca22_ha_y1;
  assign f_u_wallace_rca12_u_rca22_fa1_y3 = f_u_wallace_rca12_u_rca22_fa1_y0 & f_u_wallace_rca12_u_rca22_fa1_f_u_wallace_rca12_u_rca22_ha_y1;
  assign f_u_wallace_rca12_u_rca22_fa1_y4 = f_u_wallace_rca12_u_rca22_fa1_y1 | f_u_wallace_rca12_u_rca22_fa1_y3;
  assign f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_fa0_y2 = f_u_wallace_rca12_fa0_y2;
  assign f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_ha1_y0 = f_u_wallace_rca12_ha1_y0;
  assign f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_u_rca22_fa1_y4 = f_u_wallace_rca12_u_rca22_fa1_y4;
  assign f_u_wallace_rca12_u_rca22_fa2_y0 = f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_fa0_y2 ^ f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_ha1_y0;
  assign f_u_wallace_rca12_u_rca22_fa2_y1 = f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_fa0_y2 & f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_ha1_y0;
  assign f_u_wallace_rca12_u_rca22_fa2_y2 = f_u_wallace_rca12_u_rca22_fa2_y0 ^ f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_u_rca22_fa1_y4;
  assign f_u_wallace_rca12_u_rca22_fa2_y3 = f_u_wallace_rca12_u_rca22_fa2_y0 & f_u_wallace_rca12_u_rca22_fa2_f_u_wallace_rca12_u_rca22_fa1_y4;
  assign f_u_wallace_rca12_u_rca22_fa2_y4 = f_u_wallace_rca12_u_rca22_fa2_y1 | f_u_wallace_rca12_u_rca22_fa2_y3;
  assign f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_fa18_y2 = f_u_wallace_rca12_fa18_y2;
  assign f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_ha2_y0 = f_u_wallace_rca12_ha2_y0;
  assign f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_u_rca22_fa2_y4 = f_u_wallace_rca12_u_rca22_fa2_y4;
  assign f_u_wallace_rca12_u_rca22_fa3_y0 = f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_fa18_y2 ^ f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_ha2_y0;
  assign f_u_wallace_rca12_u_rca22_fa3_y1 = f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_fa18_y2 & f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_ha2_y0;
  assign f_u_wallace_rca12_u_rca22_fa3_y2 = f_u_wallace_rca12_u_rca22_fa3_y0 ^ f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_u_rca22_fa2_y4;
  assign f_u_wallace_rca12_u_rca22_fa3_y3 = f_u_wallace_rca12_u_rca22_fa3_y0 & f_u_wallace_rca12_u_rca22_fa3_f_u_wallace_rca12_u_rca22_fa2_y4;
  assign f_u_wallace_rca12_u_rca22_fa3_y4 = f_u_wallace_rca12_u_rca22_fa3_y1 | f_u_wallace_rca12_u_rca22_fa3_y3;
  assign f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_fa34_y2 = f_u_wallace_rca12_fa34_y2;
  assign f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_ha3_y0 = f_u_wallace_rca12_ha3_y0;
  assign f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_u_rca22_fa3_y4 = f_u_wallace_rca12_u_rca22_fa3_y4;
  assign f_u_wallace_rca12_u_rca22_fa4_y0 = f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_fa34_y2 ^ f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_ha3_y0;
  assign f_u_wallace_rca12_u_rca22_fa4_y1 = f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_fa34_y2 & f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_ha3_y0;
  assign f_u_wallace_rca12_u_rca22_fa4_y2 = f_u_wallace_rca12_u_rca22_fa4_y0 ^ f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_u_rca22_fa3_y4;
  assign f_u_wallace_rca12_u_rca22_fa4_y3 = f_u_wallace_rca12_u_rca22_fa4_y0 & f_u_wallace_rca12_u_rca22_fa4_f_u_wallace_rca12_u_rca22_fa3_y4;
  assign f_u_wallace_rca12_u_rca22_fa4_y4 = f_u_wallace_rca12_u_rca22_fa4_y1 | f_u_wallace_rca12_u_rca22_fa4_y3;
  assign f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_fa48_y2 = f_u_wallace_rca12_fa48_y2;
  assign f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_ha4_y0 = f_u_wallace_rca12_ha4_y0;
  assign f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_u_rca22_fa4_y4 = f_u_wallace_rca12_u_rca22_fa4_y4;
  assign f_u_wallace_rca12_u_rca22_fa5_y0 = f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_fa48_y2 ^ f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_ha4_y0;
  assign f_u_wallace_rca12_u_rca22_fa5_y1 = f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_fa48_y2 & f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_ha4_y0;
  assign f_u_wallace_rca12_u_rca22_fa5_y2 = f_u_wallace_rca12_u_rca22_fa5_y0 ^ f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_u_rca22_fa4_y4;
  assign f_u_wallace_rca12_u_rca22_fa5_y3 = f_u_wallace_rca12_u_rca22_fa5_y0 & f_u_wallace_rca12_u_rca22_fa5_f_u_wallace_rca12_u_rca22_fa4_y4;
  assign f_u_wallace_rca12_u_rca22_fa5_y4 = f_u_wallace_rca12_u_rca22_fa5_y1 | f_u_wallace_rca12_u_rca22_fa5_y3;
  assign f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_fa60_y2 = f_u_wallace_rca12_fa60_y2;
  assign f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_ha5_y0 = f_u_wallace_rca12_ha5_y0;
  assign f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_u_rca22_fa5_y4 = f_u_wallace_rca12_u_rca22_fa5_y4;
  assign f_u_wallace_rca12_u_rca22_fa6_y0 = f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_fa60_y2 ^ f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_ha5_y0;
  assign f_u_wallace_rca12_u_rca22_fa6_y1 = f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_fa60_y2 & f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_ha5_y0;
  assign f_u_wallace_rca12_u_rca22_fa6_y2 = f_u_wallace_rca12_u_rca22_fa6_y0 ^ f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_u_rca22_fa5_y4;
  assign f_u_wallace_rca12_u_rca22_fa6_y3 = f_u_wallace_rca12_u_rca22_fa6_y0 & f_u_wallace_rca12_u_rca22_fa6_f_u_wallace_rca12_u_rca22_fa5_y4;
  assign f_u_wallace_rca12_u_rca22_fa6_y4 = f_u_wallace_rca12_u_rca22_fa6_y1 | f_u_wallace_rca12_u_rca22_fa6_y3;
  assign f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_fa70_y2 = f_u_wallace_rca12_fa70_y2;
  assign f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_ha6_y0 = f_u_wallace_rca12_ha6_y0;
  assign f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_u_rca22_fa6_y4 = f_u_wallace_rca12_u_rca22_fa6_y4;
  assign f_u_wallace_rca12_u_rca22_fa7_y0 = f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_fa70_y2 ^ f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_ha6_y0;
  assign f_u_wallace_rca12_u_rca22_fa7_y1 = f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_fa70_y2 & f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_ha6_y0;
  assign f_u_wallace_rca12_u_rca22_fa7_y2 = f_u_wallace_rca12_u_rca22_fa7_y0 ^ f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_u_rca22_fa6_y4;
  assign f_u_wallace_rca12_u_rca22_fa7_y3 = f_u_wallace_rca12_u_rca22_fa7_y0 & f_u_wallace_rca12_u_rca22_fa7_f_u_wallace_rca12_u_rca22_fa6_y4;
  assign f_u_wallace_rca12_u_rca22_fa7_y4 = f_u_wallace_rca12_u_rca22_fa7_y1 | f_u_wallace_rca12_u_rca22_fa7_y3;
  assign f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_fa78_y2 = f_u_wallace_rca12_fa78_y2;
  assign f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_ha7_y0 = f_u_wallace_rca12_ha7_y0;
  assign f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_u_rca22_fa7_y4 = f_u_wallace_rca12_u_rca22_fa7_y4;
  assign f_u_wallace_rca12_u_rca22_fa8_y0 = f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_fa78_y2 ^ f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_ha7_y0;
  assign f_u_wallace_rca12_u_rca22_fa8_y1 = f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_fa78_y2 & f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_ha7_y0;
  assign f_u_wallace_rca12_u_rca22_fa8_y2 = f_u_wallace_rca12_u_rca22_fa8_y0 ^ f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_u_rca22_fa7_y4;
  assign f_u_wallace_rca12_u_rca22_fa8_y3 = f_u_wallace_rca12_u_rca22_fa8_y0 & f_u_wallace_rca12_u_rca22_fa8_f_u_wallace_rca12_u_rca22_fa7_y4;
  assign f_u_wallace_rca12_u_rca22_fa8_y4 = f_u_wallace_rca12_u_rca22_fa8_y1 | f_u_wallace_rca12_u_rca22_fa8_y3;
  assign f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_fa84_y2 = f_u_wallace_rca12_fa84_y2;
  assign f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_ha8_y0 = f_u_wallace_rca12_ha8_y0;
  assign f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_u_rca22_fa8_y4 = f_u_wallace_rca12_u_rca22_fa8_y4;
  assign f_u_wallace_rca12_u_rca22_fa9_y0 = f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_fa84_y2 ^ f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_ha8_y0;
  assign f_u_wallace_rca12_u_rca22_fa9_y1 = f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_fa84_y2 & f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_ha8_y0;
  assign f_u_wallace_rca12_u_rca22_fa9_y2 = f_u_wallace_rca12_u_rca22_fa9_y0 ^ f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_u_rca22_fa8_y4;
  assign f_u_wallace_rca12_u_rca22_fa9_y3 = f_u_wallace_rca12_u_rca22_fa9_y0 & f_u_wallace_rca12_u_rca22_fa9_f_u_wallace_rca12_u_rca22_fa8_y4;
  assign f_u_wallace_rca12_u_rca22_fa9_y4 = f_u_wallace_rca12_u_rca22_fa9_y1 | f_u_wallace_rca12_u_rca22_fa9_y3;
  assign f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_fa88_y2 = f_u_wallace_rca12_fa88_y2;
  assign f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_ha9_y0 = f_u_wallace_rca12_ha9_y0;
  assign f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_u_rca22_fa9_y4 = f_u_wallace_rca12_u_rca22_fa9_y4;
  assign f_u_wallace_rca12_u_rca22_fa10_y0 = f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_fa88_y2 ^ f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_ha9_y0;
  assign f_u_wallace_rca12_u_rca22_fa10_y1 = f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_fa88_y2 & f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_ha9_y0;
  assign f_u_wallace_rca12_u_rca22_fa10_y2 = f_u_wallace_rca12_u_rca22_fa10_y0 ^ f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_u_rca22_fa9_y4;
  assign f_u_wallace_rca12_u_rca22_fa10_y3 = f_u_wallace_rca12_u_rca22_fa10_y0 & f_u_wallace_rca12_u_rca22_fa10_f_u_wallace_rca12_u_rca22_fa9_y4;
  assign f_u_wallace_rca12_u_rca22_fa10_y4 = f_u_wallace_rca12_u_rca22_fa10_y1 | f_u_wallace_rca12_u_rca22_fa10_y3;
  assign f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_fa89_y2 = f_u_wallace_rca12_fa89_y2;
  assign f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_ha10_y0 = f_u_wallace_rca12_ha10_y0;
  assign f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_u_rca22_fa10_y4 = f_u_wallace_rca12_u_rca22_fa10_y4;
  assign f_u_wallace_rca12_u_rca22_fa11_y0 = f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_fa89_y2 ^ f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_ha10_y0;
  assign f_u_wallace_rca12_u_rca22_fa11_y1 = f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_fa89_y2 & f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_ha10_y0;
  assign f_u_wallace_rca12_u_rca22_fa11_y2 = f_u_wallace_rca12_u_rca22_fa11_y0 ^ f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_u_rca22_fa10_y4;
  assign f_u_wallace_rca12_u_rca22_fa11_y3 = f_u_wallace_rca12_u_rca22_fa11_y0 & f_u_wallace_rca12_u_rca22_fa11_f_u_wallace_rca12_u_rca22_fa10_y4;
  assign f_u_wallace_rca12_u_rca22_fa11_y4 = f_u_wallace_rca12_u_rca22_fa11_y1 | f_u_wallace_rca12_u_rca22_fa11_y3;
  assign f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_fa87_y2 = f_u_wallace_rca12_fa87_y2;
  assign f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_fa90_y2 = f_u_wallace_rca12_fa90_y2;
  assign f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_u_rca22_fa11_y4 = f_u_wallace_rca12_u_rca22_fa11_y4;
  assign f_u_wallace_rca12_u_rca22_fa12_y0 = f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_fa87_y2 ^ f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_fa90_y2;
  assign f_u_wallace_rca12_u_rca22_fa12_y1 = f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_fa87_y2 & f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_fa90_y2;
  assign f_u_wallace_rca12_u_rca22_fa12_y2 = f_u_wallace_rca12_u_rca22_fa12_y0 ^ f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_u_rca22_fa11_y4;
  assign f_u_wallace_rca12_u_rca22_fa12_y3 = f_u_wallace_rca12_u_rca22_fa12_y0 & f_u_wallace_rca12_u_rca22_fa12_f_u_wallace_rca12_u_rca22_fa11_y4;
  assign f_u_wallace_rca12_u_rca22_fa12_y4 = f_u_wallace_rca12_u_rca22_fa12_y1 | f_u_wallace_rca12_u_rca22_fa12_y3;
  assign f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_fa83_y2 = f_u_wallace_rca12_fa83_y2;
  assign f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_fa91_y2 = f_u_wallace_rca12_fa91_y2;
  assign f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_u_rca22_fa12_y4 = f_u_wallace_rca12_u_rca22_fa12_y4;
  assign f_u_wallace_rca12_u_rca22_fa13_y0 = f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_fa83_y2 ^ f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_fa91_y2;
  assign f_u_wallace_rca12_u_rca22_fa13_y1 = f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_fa83_y2 & f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_fa91_y2;
  assign f_u_wallace_rca12_u_rca22_fa13_y2 = f_u_wallace_rca12_u_rca22_fa13_y0 ^ f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_u_rca22_fa12_y4;
  assign f_u_wallace_rca12_u_rca22_fa13_y3 = f_u_wallace_rca12_u_rca22_fa13_y0 & f_u_wallace_rca12_u_rca22_fa13_f_u_wallace_rca12_u_rca22_fa12_y4;
  assign f_u_wallace_rca12_u_rca22_fa13_y4 = f_u_wallace_rca12_u_rca22_fa13_y1 | f_u_wallace_rca12_u_rca22_fa13_y3;
  assign f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_fa77_y2 = f_u_wallace_rca12_fa77_y2;
  assign f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_fa92_y2 = f_u_wallace_rca12_fa92_y2;
  assign f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_u_rca22_fa13_y4 = f_u_wallace_rca12_u_rca22_fa13_y4;
  assign f_u_wallace_rca12_u_rca22_fa14_y0 = f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_fa77_y2 ^ f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_fa92_y2;
  assign f_u_wallace_rca12_u_rca22_fa14_y1 = f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_fa77_y2 & f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_fa92_y2;
  assign f_u_wallace_rca12_u_rca22_fa14_y2 = f_u_wallace_rca12_u_rca22_fa14_y0 ^ f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_u_rca22_fa13_y4;
  assign f_u_wallace_rca12_u_rca22_fa14_y3 = f_u_wallace_rca12_u_rca22_fa14_y0 & f_u_wallace_rca12_u_rca22_fa14_f_u_wallace_rca12_u_rca22_fa13_y4;
  assign f_u_wallace_rca12_u_rca22_fa14_y4 = f_u_wallace_rca12_u_rca22_fa14_y1 | f_u_wallace_rca12_u_rca22_fa14_y3;
  assign f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_fa69_y2 = f_u_wallace_rca12_fa69_y2;
  assign f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_fa93_y2 = f_u_wallace_rca12_fa93_y2;
  assign f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_u_rca22_fa14_y4 = f_u_wallace_rca12_u_rca22_fa14_y4;
  assign f_u_wallace_rca12_u_rca22_fa15_y0 = f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_fa69_y2 ^ f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_fa93_y2;
  assign f_u_wallace_rca12_u_rca22_fa15_y1 = f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_fa69_y2 & f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_fa93_y2;
  assign f_u_wallace_rca12_u_rca22_fa15_y2 = f_u_wallace_rca12_u_rca22_fa15_y0 ^ f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_u_rca22_fa14_y4;
  assign f_u_wallace_rca12_u_rca22_fa15_y3 = f_u_wallace_rca12_u_rca22_fa15_y0 & f_u_wallace_rca12_u_rca22_fa15_f_u_wallace_rca12_u_rca22_fa14_y4;
  assign f_u_wallace_rca12_u_rca22_fa15_y4 = f_u_wallace_rca12_u_rca22_fa15_y1 | f_u_wallace_rca12_u_rca22_fa15_y3;
  assign f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_fa59_y2 = f_u_wallace_rca12_fa59_y2;
  assign f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_fa94_y2 = f_u_wallace_rca12_fa94_y2;
  assign f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_u_rca22_fa15_y4 = f_u_wallace_rca12_u_rca22_fa15_y4;
  assign f_u_wallace_rca12_u_rca22_fa16_y0 = f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_fa59_y2 ^ f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_fa94_y2;
  assign f_u_wallace_rca12_u_rca22_fa16_y1 = f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_fa59_y2 & f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_fa94_y2;
  assign f_u_wallace_rca12_u_rca22_fa16_y2 = f_u_wallace_rca12_u_rca22_fa16_y0 ^ f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_u_rca22_fa15_y4;
  assign f_u_wallace_rca12_u_rca22_fa16_y3 = f_u_wallace_rca12_u_rca22_fa16_y0 & f_u_wallace_rca12_u_rca22_fa16_f_u_wallace_rca12_u_rca22_fa15_y4;
  assign f_u_wallace_rca12_u_rca22_fa16_y4 = f_u_wallace_rca12_u_rca22_fa16_y1 | f_u_wallace_rca12_u_rca22_fa16_y3;
  assign f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_fa47_y2 = f_u_wallace_rca12_fa47_y2;
  assign f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_fa95_y2 = f_u_wallace_rca12_fa95_y2;
  assign f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_u_rca22_fa16_y4 = f_u_wallace_rca12_u_rca22_fa16_y4;
  assign f_u_wallace_rca12_u_rca22_fa17_y0 = f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_fa47_y2 ^ f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_fa95_y2;
  assign f_u_wallace_rca12_u_rca22_fa17_y1 = f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_fa47_y2 & f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_fa95_y2;
  assign f_u_wallace_rca12_u_rca22_fa17_y2 = f_u_wallace_rca12_u_rca22_fa17_y0 ^ f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_u_rca22_fa16_y4;
  assign f_u_wallace_rca12_u_rca22_fa17_y3 = f_u_wallace_rca12_u_rca22_fa17_y0 & f_u_wallace_rca12_u_rca22_fa17_f_u_wallace_rca12_u_rca22_fa16_y4;
  assign f_u_wallace_rca12_u_rca22_fa17_y4 = f_u_wallace_rca12_u_rca22_fa17_y1 | f_u_wallace_rca12_u_rca22_fa17_y3;
  assign f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_fa33_y2 = f_u_wallace_rca12_fa33_y2;
  assign f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_fa96_y2 = f_u_wallace_rca12_fa96_y2;
  assign f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_u_rca22_fa17_y4 = f_u_wallace_rca12_u_rca22_fa17_y4;
  assign f_u_wallace_rca12_u_rca22_fa18_y0 = f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_fa33_y2 ^ f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_fa96_y2;
  assign f_u_wallace_rca12_u_rca22_fa18_y1 = f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_fa33_y2 & f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_fa96_y2;
  assign f_u_wallace_rca12_u_rca22_fa18_y2 = f_u_wallace_rca12_u_rca22_fa18_y0 ^ f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_u_rca22_fa17_y4;
  assign f_u_wallace_rca12_u_rca22_fa18_y3 = f_u_wallace_rca12_u_rca22_fa18_y0 & f_u_wallace_rca12_u_rca22_fa18_f_u_wallace_rca12_u_rca22_fa17_y4;
  assign f_u_wallace_rca12_u_rca22_fa18_y4 = f_u_wallace_rca12_u_rca22_fa18_y1 | f_u_wallace_rca12_u_rca22_fa18_y3;
  assign f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_fa17_y2 = f_u_wallace_rca12_fa17_y2;
  assign f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_fa97_y2 = f_u_wallace_rca12_fa97_y2;
  assign f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_u_rca22_fa18_y4 = f_u_wallace_rca12_u_rca22_fa18_y4;
  assign f_u_wallace_rca12_u_rca22_fa19_y0 = f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_fa17_y2 ^ f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_fa97_y2;
  assign f_u_wallace_rca12_u_rca22_fa19_y1 = f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_fa17_y2 & f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_fa97_y2;
  assign f_u_wallace_rca12_u_rca22_fa19_y2 = f_u_wallace_rca12_u_rca22_fa19_y0 ^ f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_u_rca22_fa18_y4;
  assign f_u_wallace_rca12_u_rca22_fa19_y3 = f_u_wallace_rca12_u_rca22_fa19_y0 & f_u_wallace_rca12_u_rca22_fa19_f_u_wallace_rca12_u_rca22_fa18_y4;
  assign f_u_wallace_rca12_u_rca22_fa19_y4 = f_u_wallace_rca12_u_rca22_fa19_y1 | f_u_wallace_rca12_u_rca22_fa19_y3;
  assign f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_and_10_11_y0 = f_u_wallace_rca12_and_10_11_y0;
  assign f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_fa98_y2 = f_u_wallace_rca12_fa98_y2;
  assign f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_u_rca22_fa19_y4 = f_u_wallace_rca12_u_rca22_fa19_y4;
  assign f_u_wallace_rca12_u_rca22_fa20_y0 = f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_and_10_11_y0 ^ f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_fa98_y2;
  assign f_u_wallace_rca12_u_rca22_fa20_y1 = f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_and_10_11_y0 & f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_fa98_y2;
  assign f_u_wallace_rca12_u_rca22_fa20_y2 = f_u_wallace_rca12_u_rca22_fa20_y0 ^ f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_u_rca22_fa19_y4;
  assign f_u_wallace_rca12_u_rca22_fa20_y3 = f_u_wallace_rca12_u_rca22_fa20_y0 & f_u_wallace_rca12_u_rca22_fa20_f_u_wallace_rca12_u_rca22_fa19_y4;
  assign f_u_wallace_rca12_u_rca22_fa20_y4 = f_u_wallace_rca12_u_rca22_fa20_y1 | f_u_wallace_rca12_u_rca22_fa20_y3;
  assign f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_fa98_y4 = f_u_wallace_rca12_fa98_y4;
  assign f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_and_11_11_y0 = f_u_wallace_rca12_and_11_11_y0;
  assign f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_u_rca22_fa20_y4 = f_u_wallace_rca12_u_rca22_fa20_y4;
  assign f_u_wallace_rca12_u_rca22_fa21_y0 = f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_fa98_y4 ^ f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_and_11_11_y0;
  assign f_u_wallace_rca12_u_rca22_fa21_y1 = f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_fa98_y4 & f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_and_11_11_y0;
  assign f_u_wallace_rca12_u_rca22_fa21_y2 = f_u_wallace_rca12_u_rca22_fa21_y0 ^ f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_u_rca22_fa20_y4;
  assign f_u_wallace_rca12_u_rca22_fa21_y3 = f_u_wallace_rca12_u_rca22_fa21_y0 & f_u_wallace_rca12_u_rca22_fa21_f_u_wallace_rca12_u_rca22_fa20_y4;
  assign f_u_wallace_rca12_u_rca22_fa21_y4 = f_u_wallace_rca12_u_rca22_fa21_y1 | f_u_wallace_rca12_u_rca22_fa21_y3;

  assign out[0] = f_u_wallace_rca12_and_0_0_y0;
  assign out[1] = f_u_wallace_rca12_u_rca22_ha_y0;
  assign out[2] = f_u_wallace_rca12_u_rca22_fa1_y2;
  assign out[3] = f_u_wallace_rca12_u_rca22_fa2_y2;
  assign out[4] = f_u_wallace_rca12_u_rca22_fa3_y2;
  assign out[5] = f_u_wallace_rca12_u_rca22_fa4_y2;
  assign out[6] = f_u_wallace_rca12_u_rca22_fa5_y2;
  assign out[7] = f_u_wallace_rca12_u_rca22_fa6_y2;
  assign out[8] = f_u_wallace_rca12_u_rca22_fa7_y2;
  assign out[9] = f_u_wallace_rca12_u_rca22_fa8_y2;
  assign out[10] = f_u_wallace_rca12_u_rca22_fa9_y2;
  assign out[11] = f_u_wallace_rca12_u_rca22_fa10_y2;
  assign out[12] = f_u_wallace_rca12_u_rca22_fa11_y2;
  assign out[13] = f_u_wallace_rca12_u_rca22_fa12_y2;
  assign out[14] = f_u_wallace_rca12_u_rca22_fa13_y2;
  assign out[15] = f_u_wallace_rca12_u_rca22_fa14_y2;
  assign out[16] = f_u_wallace_rca12_u_rca22_fa15_y2;
  assign out[17] = f_u_wallace_rca12_u_rca22_fa16_y2;
  assign out[18] = f_u_wallace_rca12_u_rca22_fa17_y2;
  assign out[19] = f_u_wallace_rca12_u_rca22_fa18_y2;
  assign out[20] = f_u_wallace_rca12_u_rca22_fa19_y2;
  assign out[21] = f_u_wallace_rca12_u_rca22_fa20_y2;
  assign out[22] = f_u_wallace_rca12_u_rca22_fa21_y2;
  assign out[23] = f_u_wallace_rca12_u_rca22_fa21_y4;
endmodule