module f_u_arrbam8_h6_v6(input [7:0] a, input [7:0] b, output [15:0] f_u_arrbam8_h6_v6_out);
  wire f_u_arrbam8_h6_v6_and0_6;
  wire f_u_arrbam8_h6_v6_and1_6;
  wire f_u_arrbam8_h6_v6_and2_6;
  wire f_u_arrbam8_h6_v6_and3_6;
  wire f_u_arrbam8_h6_v6_and4_6;
  wire f_u_arrbam8_h6_v6_and5_6;
  wire f_u_arrbam8_h6_v6_and6_6;
  wire f_u_arrbam8_h6_v6_and7_6;
  wire f_u_arrbam8_h6_v6_and0_7;
  wire f_u_arrbam8_h6_v6_ha0_7_xor0;
  wire f_u_arrbam8_h6_v6_ha0_7_and0;
  wire f_u_arrbam8_h6_v6_and1_7;
  wire f_u_arrbam8_h6_v6_fa1_7_xor0;
  wire f_u_arrbam8_h6_v6_fa1_7_and0;
  wire f_u_arrbam8_h6_v6_fa1_7_xor1;
  wire f_u_arrbam8_h6_v6_fa1_7_and1;
  wire f_u_arrbam8_h6_v6_fa1_7_or0;
  wire f_u_arrbam8_h6_v6_and2_7;
  wire f_u_arrbam8_h6_v6_fa2_7_xor0;
  wire f_u_arrbam8_h6_v6_fa2_7_and0;
  wire f_u_arrbam8_h6_v6_fa2_7_xor1;
  wire f_u_arrbam8_h6_v6_fa2_7_and1;
  wire f_u_arrbam8_h6_v6_fa2_7_or0;
  wire f_u_arrbam8_h6_v6_and3_7;
  wire f_u_arrbam8_h6_v6_fa3_7_xor0;
  wire f_u_arrbam8_h6_v6_fa3_7_and0;
  wire f_u_arrbam8_h6_v6_fa3_7_xor1;
  wire f_u_arrbam8_h6_v6_fa3_7_and1;
  wire f_u_arrbam8_h6_v6_fa3_7_or0;
  wire f_u_arrbam8_h6_v6_and4_7;
  wire f_u_arrbam8_h6_v6_fa4_7_xor0;
  wire f_u_arrbam8_h6_v6_fa4_7_and0;
  wire f_u_arrbam8_h6_v6_fa4_7_xor1;
  wire f_u_arrbam8_h6_v6_fa4_7_and1;
  wire f_u_arrbam8_h6_v6_fa4_7_or0;
  wire f_u_arrbam8_h6_v6_and5_7;
  wire f_u_arrbam8_h6_v6_fa5_7_xor0;
  wire f_u_arrbam8_h6_v6_fa5_7_and0;
  wire f_u_arrbam8_h6_v6_fa5_7_xor1;
  wire f_u_arrbam8_h6_v6_fa5_7_and1;
  wire f_u_arrbam8_h6_v6_fa5_7_or0;
  wire f_u_arrbam8_h6_v6_and6_7;
  wire f_u_arrbam8_h6_v6_fa6_7_xor0;
  wire f_u_arrbam8_h6_v6_fa6_7_and0;
  wire f_u_arrbam8_h6_v6_fa6_7_xor1;
  wire f_u_arrbam8_h6_v6_fa6_7_and1;
  wire f_u_arrbam8_h6_v6_fa6_7_or0;
  wire f_u_arrbam8_h6_v6_and7_7;
  wire f_u_arrbam8_h6_v6_ha7_7_xor0;
  wire f_u_arrbam8_h6_v6_ha7_7_and0;

  assign f_u_arrbam8_h6_v6_and0_6 = a[0] & b[6];
  assign f_u_arrbam8_h6_v6_and1_6 = a[1] & b[6];
  assign f_u_arrbam8_h6_v6_and2_6 = a[2] & b[6];
  assign f_u_arrbam8_h6_v6_and3_6 = a[3] & b[6];
  assign f_u_arrbam8_h6_v6_and4_6 = a[4] & b[6];
  assign f_u_arrbam8_h6_v6_and5_6 = a[5] & b[6];
  assign f_u_arrbam8_h6_v6_and6_6 = a[6] & b[6];
  assign f_u_arrbam8_h6_v6_and7_6 = a[7] & b[6];
  assign f_u_arrbam8_h6_v6_and0_7 = a[0] & b[7];
  assign f_u_arrbam8_h6_v6_ha0_7_xor0 = f_u_arrbam8_h6_v6_and0_7 ^ f_u_arrbam8_h6_v6_and1_6;
  assign f_u_arrbam8_h6_v6_ha0_7_and0 = f_u_arrbam8_h6_v6_and0_7 & f_u_arrbam8_h6_v6_and1_6;
  assign f_u_arrbam8_h6_v6_and1_7 = a[1] & b[7];
  assign f_u_arrbam8_h6_v6_fa1_7_xor0 = f_u_arrbam8_h6_v6_and1_7 ^ f_u_arrbam8_h6_v6_and2_6;
  assign f_u_arrbam8_h6_v6_fa1_7_and0 = f_u_arrbam8_h6_v6_and1_7 & f_u_arrbam8_h6_v6_and2_6;
  assign f_u_arrbam8_h6_v6_fa1_7_xor1 = f_u_arrbam8_h6_v6_fa1_7_xor0 ^ f_u_arrbam8_h6_v6_ha0_7_and0;
  assign f_u_arrbam8_h6_v6_fa1_7_and1 = f_u_arrbam8_h6_v6_fa1_7_xor0 & f_u_arrbam8_h6_v6_ha0_7_and0;
  assign f_u_arrbam8_h6_v6_fa1_7_or0 = f_u_arrbam8_h6_v6_fa1_7_and0 | f_u_arrbam8_h6_v6_fa1_7_and1;
  assign f_u_arrbam8_h6_v6_and2_7 = a[2] & b[7];
  assign f_u_arrbam8_h6_v6_fa2_7_xor0 = f_u_arrbam8_h6_v6_and2_7 ^ f_u_arrbam8_h6_v6_and3_6;
  assign f_u_arrbam8_h6_v6_fa2_7_and0 = f_u_arrbam8_h6_v6_and2_7 & f_u_arrbam8_h6_v6_and3_6;
  assign f_u_arrbam8_h6_v6_fa2_7_xor1 = f_u_arrbam8_h6_v6_fa2_7_xor0 ^ f_u_arrbam8_h6_v6_fa1_7_or0;
  assign f_u_arrbam8_h6_v6_fa2_7_and1 = f_u_arrbam8_h6_v6_fa2_7_xor0 & f_u_arrbam8_h6_v6_fa1_7_or0;
  assign f_u_arrbam8_h6_v6_fa2_7_or0 = f_u_arrbam8_h6_v6_fa2_7_and0 | f_u_arrbam8_h6_v6_fa2_7_and1;
  assign f_u_arrbam8_h6_v6_and3_7 = a[3] & b[7];
  assign f_u_arrbam8_h6_v6_fa3_7_xor0 = f_u_arrbam8_h6_v6_and3_7 ^ f_u_arrbam8_h6_v6_and4_6;
  assign f_u_arrbam8_h6_v6_fa3_7_and0 = f_u_arrbam8_h6_v6_and3_7 & f_u_arrbam8_h6_v6_and4_6;
  assign f_u_arrbam8_h6_v6_fa3_7_xor1 = f_u_arrbam8_h6_v6_fa3_7_xor0 ^ f_u_arrbam8_h6_v6_fa2_7_or0;
  assign f_u_arrbam8_h6_v6_fa3_7_and1 = f_u_arrbam8_h6_v6_fa3_7_xor0 & f_u_arrbam8_h6_v6_fa2_7_or0;
  assign f_u_arrbam8_h6_v6_fa3_7_or0 = f_u_arrbam8_h6_v6_fa3_7_and0 | f_u_arrbam8_h6_v6_fa3_7_and1;
  assign f_u_arrbam8_h6_v6_and4_7 = a[4] & b[7];
  assign f_u_arrbam8_h6_v6_fa4_7_xor0 = f_u_arrbam8_h6_v6_and4_7 ^ f_u_arrbam8_h6_v6_and5_6;
  assign f_u_arrbam8_h6_v6_fa4_7_and0 = f_u_arrbam8_h6_v6_and4_7 & f_u_arrbam8_h6_v6_and5_6;
  assign f_u_arrbam8_h6_v6_fa4_7_xor1 = f_u_arrbam8_h6_v6_fa4_7_xor0 ^ f_u_arrbam8_h6_v6_fa3_7_or0;
  assign f_u_arrbam8_h6_v6_fa4_7_and1 = f_u_arrbam8_h6_v6_fa4_7_xor0 & f_u_arrbam8_h6_v6_fa3_7_or0;
  assign f_u_arrbam8_h6_v6_fa4_7_or0 = f_u_arrbam8_h6_v6_fa4_7_and0 | f_u_arrbam8_h6_v6_fa4_7_and1;
  assign f_u_arrbam8_h6_v6_and5_7 = a[5] & b[7];
  assign f_u_arrbam8_h6_v6_fa5_7_xor0 = f_u_arrbam8_h6_v6_and5_7 ^ f_u_arrbam8_h6_v6_and6_6;
  assign f_u_arrbam8_h6_v6_fa5_7_and0 = f_u_arrbam8_h6_v6_and5_7 & f_u_arrbam8_h6_v6_and6_6;
  assign f_u_arrbam8_h6_v6_fa5_7_xor1 = f_u_arrbam8_h6_v6_fa5_7_xor0 ^ f_u_arrbam8_h6_v6_fa4_7_or0;
  assign f_u_arrbam8_h6_v6_fa5_7_and1 = f_u_arrbam8_h6_v6_fa5_7_xor0 & f_u_arrbam8_h6_v6_fa4_7_or0;
  assign f_u_arrbam8_h6_v6_fa5_7_or0 = f_u_arrbam8_h6_v6_fa5_7_and0 | f_u_arrbam8_h6_v6_fa5_7_and1;
  assign f_u_arrbam8_h6_v6_and6_7 = a[6] & b[7];
  assign f_u_arrbam8_h6_v6_fa6_7_xor0 = f_u_arrbam8_h6_v6_and6_7 ^ f_u_arrbam8_h6_v6_and7_6;
  assign f_u_arrbam8_h6_v6_fa6_7_and0 = f_u_arrbam8_h6_v6_and6_7 & f_u_arrbam8_h6_v6_and7_6;
  assign f_u_arrbam8_h6_v6_fa6_7_xor1 = f_u_arrbam8_h6_v6_fa6_7_xor0 ^ f_u_arrbam8_h6_v6_fa5_7_or0;
  assign f_u_arrbam8_h6_v6_fa6_7_and1 = f_u_arrbam8_h6_v6_fa6_7_xor0 & f_u_arrbam8_h6_v6_fa5_7_or0;
  assign f_u_arrbam8_h6_v6_fa6_7_or0 = f_u_arrbam8_h6_v6_fa6_7_and0 | f_u_arrbam8_h6_v6_fa6_7_and1;
  assign f_u_arrbam8_h6_v6_and7_7 = a[7] & b[7];
  assign f_u_arrbam8_h6_v6_ha7_7_xor0 = f_u_arrbam8_h6_v6_and7_7 ^ f_u_arrbam8_h6_v6_fa6_7_or0;
  assign f_u_arrbam8_h6_v6_ha7_7_and0 = f_u_arrbam8_h6_v6_and7_7 & f_u_arrbam8_h6_v6_fa6_7_or0;

  assign f_u_arrbam8_h6_v6_out[0] = 1'b0;
  assign f_u_arrbam8_h6_v6_out[1] = 1'b0;
  assign f_u_arrbam8_h6_v6_out[2] = 1'b0;
  assign f_u_arrbam8_h6_v6_out[3] = 1'b0;
  assign f_u_arrbam8_h6_v6_out[4] = 1'b0;
  assign f_u_arrbam8_h6_v6_out[5] = 1'b0;
  assign f_u_arrbam8_h6_v6_out[6] = f_u_arrbam8_h6_v6_and0_6;
  assign f_u_arrbam8_h6_v6_out[7] = f_u_arrbam8_h6_v6_ha0_7_xor0;
  assign f_u_arrbam8_h6_v6_out[8] = f_u_arrbam8_h6_v6_fa1_7_xor1;
  assign f_u_arrbam8_h6_v6_out[9] = f_u_arrbam8_h6_v6_fa2_7_xor1;
  assign f_u_arrbam8_h6_v6_out[10] = f_u_arrbam8_h6_v6_fa3_7_xor1;
  assign f_u_arrbam8_h6_v6_out[11] = f_u_arrbam8_h6_v6_fa4_7_xor1;
  assign f_u_arrbam8_h6_v6_out[12] = f_u_arrbam8_h6_v6_fa5_7_xor1;
  assign f_u_arrbam8_h6_v6_out[13] = f_u_arrbam8_h6_v6_fa6_7_xor1;
  assign f_u_arrbam8_h6_v6_out[14] = f_u_arrbam8_h6_v6_ha7_7_xor0;
  assign f_u_arrbam8_h6_v6_out[15] = f_u_arrbam8_h6_v6_ha7_7_and0;
endmodule