module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module fs(input [0:0] a, input [0:0] b, input [0:0] bin, output [0:0] fs_xor1, output [0:0] fs_or0);
  wire [0:0] fs_xor0;
  wire [0:0] fs_not0;
  wire [0:0] fs_and0;
  wire [0:0] fs_not1;
  wire [0:0] fs_and1;
  xor_gate xor_gate_fs_xor0(.a(a[0]), .b(b[0]), .out(fs_xor0));
  not_gate not_gate_fs_not0(.a(a[0]), .out(fs_not0));
  and_gate and_gate_fs_and0(.a(fs_not0[0]), .b(b[0]), .out(fs_and0));
  xor_gate xor_gate_fs_xor1(.a(bin[0]), .b(fs_xor0[0]), .out(fs_xor1));
  not_gate not_gate_fs_not1(.a(fs_xor0[0]), .out(fs_not1));
  and_gate and_gate_fs_and1(.a(fs_not1[0]), .b(bin[0]), .out(fs_and1));
  or_gate or_gate_fs_or0(.a(fs_and1[0]), .b(fs_and0[0]), .out(fs_or0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module h_arrdiv8(input [7:0] a, input [7:0] b, output [7:0] h_arrdiv8_out);
  wire [0:0] h_arrdiv8_fs0_xor0;
  wire [0:0] h_arrdiv8_fs0_and0;
  wire [0:0] h_arrdiv8_fs1_xor1;
  wire [0:0] h_arrdiv8_fs1_or0;
  wire [0:0] h_arrdiv8_fs2_xor1;
  wire [0:0] h_arrdiv8_fs2_or0;
  wire [0:0] h_arrdiv8_fs3_xor1;
  wire [0:0] h_arrdiv8_fs3_or0;
  wire [0:0] h_arrdiv8_fs4_xor1;
  wire [0:0] h_arrdiv8_fs4_or0;
  wire [0:0] h_arrdiv8_fs5_xor1;
  wire [0:0] h_arrdiv8_fs5_or0;
  wire [0:0] h_arrdiv8_fs6_xor1;
  wire [0:0] h_arrdiv8_fs6_or0;
  wire [0:0] h_arrdiv8_fs7_xor1;
  wire [0:0] h_arrdiv8_fs7_or0;
  wire [0:0] h_arrdiv8_mux2to10_xor0;
  wire [0:0] h_arrdiv8_mux2to11_and1;
  wire [0:0] h_arrdiv8_mux2to12_and1;
  wire [0:0] h_arrdiv8_mux2to13_and1;
  wire [0:0] h_arrdiv8_mux2to14_and1;
  wire [0:0] h_arrdiv8_mux2to15_and1;
  wire [0:0] h_arrdiv8_mux2to16_and1;
  wire [0:0] h_arrdiv8_not0;
  wire [0:0] h_arrdiv8_fs8_xor0;
  wire [0:0] h_arrdiv8_fs8_and0;
  wire [0:0] h_arrdiv8_fs9_xor1;
  wire [0:0] h_arrdiv8_fs9_or0;
  wire [0:0] h_arrdiv8_fs10_xor1;
  wire [0:0] h_arrdiv8_fs10_or0;
  wire [0:0] h_arrdiv8_fs11_xor1;
  wire [0:0] h_arrdiv8_fs11_or0;
  wire [0:0] h_arrdiv8_fs12_xor1;
  wire [0:0] h_arrdiv8_fs12_or0;
  wire [0:0] h_arrdiv8_fs13_xor1;
  wire [0:0] h_arrdiv8_fs13_or0;
  wire [0:0] h_arrdiv8_fs14_xor1;
  wire [0:0] h_arrdiv8_fs14_or0;
  wire [0:0] h_arrdiv8_fs15_xor1;
  wire [0:0] h_arrdiv8_fs15_or0;
  wire [0:0] h_arrdiv8_mux2to17_xor0;
  wire [0:0] h_arrdiv8_mux2to18_xor0;
  wire [0:0] h_arrdiv8_mux2to19_xor0;
  wire [0:0] h_arrdiv8_mux2to110_xor0;
  wire [0:0] h_arrdiv8_mux2to111_xor0;
  wire [0:0] h_arrdiv8_mux2to112_xor0;
  wire [0:0] h_arrdiv8_mux2to113_xor0;
  wire [0:0] h_arrdiv8_not1;
  wire [0:0] h_arrdiv8_fs16_xor0;
  wire [0:0] h_arrdiv8_fs16_and0;
  wire [0:0] h_arrdiv8_fs17_xor1;
  wire [0:0] h_arrdiv8_fs17_or0;
  wire [0:0] h_arrdiv8_fs18_xor1;
  wire [0:0] h_arrdiv8_fs18_or0;
  wire [0:0] h_arrdiv8_fs19_xor1;
  wire [0:0] h_arrdiv8_fs19_or0;
  wire [0:0] h_arrdiv8_fs20_xor1;
  wire [0:0] h_arrdiv8_fs20_or0;
  wire [0:0] h_arrdiv8_fs21_xor1;
  wire [0:0] h_arrdiv8_fs21_or0;
  wire [0:0] h_arrdiv8_fs22_xor1;
  wire [0:0] h_arrdiv8_fs22_or0;
  wire [0:0] h_arrdiv8_fs23_xor1;
  wire [0:0] h_arrdiv8_fs23_or0;
  wire [0:0] h_arrdiv8_mux2to114_xor0;
  wire [0:0] h_arrdiv8_mux2to115_xor0;
  wire [0:0] h_arrdiv8_mux2to116_xor0;
  wire [0:0] h_arrdiv8_mux2to117_xor0;
  wire [0:0] h_arrdiv8_mux2to118_xor0;
  wire [0:0] h_arrdiv8_mux2to119_xor0;
  wire [0:0] h_arrdiv8_mux2to120_xor0;
  wire [0:0] h_arrdiv8_not2;
  wire [0:0] h_arrdiv8_fs24_xor0;
  wire [0:0] h_arrdiv8_fs24_and0;
  wire [0:0] h_arrdiv8_fs25_xor1;
  wire [0:0] h_arrdiv8_fs25_or0;
  wire [0:0] h_arrdiv8_fs26_xor1;
  wire [0:0] h_arrdiv8_fs26_or0;
  wire [0:0] h_arrdiv8_fs27_xor1;
  wire [0:0] h_arrdiv8_fs27_or0;
  wire [0:0] h_arrdiv8_fs28_xor1;
  wire [0:0] h_arrdiv8_fs28_or0;
  wire [0:0] h_arrdiv8_fs29_xor1;
  wire [0:0] h_arrdiv8_fs29_or0;
  wire [0:0] h_arrdiv8_fs30_xor1;
  wire [0:0] h_arrdiv8_fs30_or0;
  wire [0:0] h_arrdiv8_fs31_xor1;
  wire [0:0] h_arrdiv8_fs31_or0;
  wire [0:0] h_arrdiv8_mux2to121_xor0;
  wire [0:0] h_arrdiv8_mux2to122_xor0;
  wire [0:0] h_arrdiv8_mux2to123_xor0;
  wire [0:0] h_arrdiv8_mux2to124_xor0;
  wire [0:0] h_arrdiv8_mux2to125_xor0;
  wire [0:0] h_arrdiv8_mux2to126_xor0;
  wire [0:0] h_arrdiv8_mux2to127_xor0;
  wire [0:0] h_arrdiv8_not3;
  wire [0:0] h_arrdiv8_fs32_xor0;
  wire [0:0] h_arrdiv8_fs32_and0;
  wire [0:0] h_arrdiv8_fs33_xor1;
  wire [0:0] h_arrdiv8_fs33_or0;
  wire [0:0] h_arrdiv8_fs34_xor1;
  wire [0:0] h_arrdiv8_fs34_or0;
  wire [0:0] h_arrdiv8_fs35_xor1;
  wire [0:0] h_arrdiv8_fs35_or0;
  wire [0:0] h_arrdiv8_fs36_xor1;
  wire [0:0] h_arrdiv8_fs36_or0;
  wire [0:0] h_arrdiv8_fs37_xor1;
  wire [0:0] h_arrdiv8_fs37_or0;
  wire [0:0] h_arrdiv8_fs38_xor1;
  wire [0:0] h_arrdiv8_fs38_or0;
  wire [0:0] h_arrdiv8_fs39_xor1;
  wire [0:0] h_arrdiv8_fs39_or0;
  wire [0:0] h_arrdiv8_mux2to128_xor0;
  wire [0:0] h_arrdiv8_mux2to129_xor0;
  wire [0:0] h_arrdiv8_mux2to130_xor0;
  wire [0:0] h_arrdiv8_mux2to131_xor0;
  wire [0:0] h_arrdiv8_mux2to132_xor0;
  wire [0:0] h_arrdiv8_mux2to133_xor0;
  wire [0:0] h_arrdiv8_mux2to134_xor0;
  wire [0:0] h_arrdiv8_not4;
  wire [0:0] h_arrdiv8_fs40_xor0;
  wire [0:0] h_arrdiv8_fs40_and0;
  wire [0:0] h_arrdiv8_fs41_xor1;
  wire [0:0] h_arrdiv8_fs41_or0;
  wire [0:0] h_arrdiv8_fs42_xor1;
  wire [0:0] h_arrdiv8_fs42_or0;
  wire [0:0] h_arrdiv8_fs43_xor1;
  wire [0:0] h_arrdiv8_fs43_or0;
  wire [0:0] h_arrdiv8_fs44_xor1;
  wire [0:0] h_arrdiv8_fs44_or0;
  wire [0:0] h_arrdiv8_fs45_xor1;
  wire [0:0] h_arrdiv8_fs45_or0;
  wire [0:0] h_arrdiv8_fs46_xor1;
  wire [0:0] h_arrdiv8_fs46_or0;
  wire [0:0] h_arrdiv8_fs47_xor1;
  wire [0:0] h_arrdiv8_fs47_or0;
  wire [0:0] h_arrdiv8_mux2to135_xor0;
  wire [0:0] h_arrdiv8_mux2to136_xor0;
  wire [0:0] h_arrdiv8_mux2to137_xor0;
  wire [0:0] h_arrdiv8_mux2to138_xor0;
  wire [0:0] h_arrdiv8_mux2to139_xor0;
  wire [0:0] h_arrdiv8_mux2to140_xor0;
  wire [0:0] h_arrdiv8_mux2to141_xor0;
  wire [0:0] h_arrdiv8_not5;
  wire [0:0] h_arrdiv8_fs48_xor0;
  wire [0:0] h_arrdiv8_fs48_and0;
  wire [0:0] h_arrdiv8_fs49_xor1;
  wire [0:0] h_arrdiv8_fs49_or0;
  wire [0:0] h_arrdiv8_fs50_xor1;
  wire [0:0] h_arrdiv8_fs50_or0;
  wire [0:0] h_arrdiv8_fs51_xor1;
  wire [0:0] h_arrdiv8_fs51_or0;
  wire [0:0] h_arrdiv8_fs52_xor1;
  wire [0:0] h_arrdiv8_fs52_or0;
  wire [0:0] h_arrdiv8_fs53_xor1;
  wire [0:0] h_arrdiv8_fs53_or0;
  wire [0:0] h_arrdiv8_fs54_xor1;
  wire [0:0] h_arrdiv8_fs54_or0;
  wire [0:0] h_arrdiv8_fs55_xor1;
  wire [0:0] h_arrdiv8_fs55_or0;
  wire [0:0] h_arrdiv8_mux2to142_xor0;
  wire [0:0] h_arrdiv8_mux2to143_xor0;
  wire [0:0] h_arrdiv8_mux2to144_xor0;
  wire [0:0] h_arrdiv8_mux2to145_xor0;
  wire [0:0] h_arrdiv8_mux2to146_xor0;
  wire [0:0] h_arrdiv8_mux2to147_xor0;
  wire [0:0] h_arrdiv8_mux2to148_xor0;
  wire [0:0] h_arrdiv8_not6;
  wire [0:0] h_arrdiv8_fs56_xor0;
  wire [0:0] h_arrdiv8_fs56_and0;
  wire [0:0] h_arrdiv8_fs57_xor1;
  wire [0:0] h_arrdiv8_fs57_or0;
  wire [0:0] h_arrdiv8_fs58_xor1;
  wire [0:0] h_arrdiv8_fs58_or0;
  wire [0:0] h_arrdiv8_fs59_xor1;
  wire [0:0] h_arrdiv8_fs59_or0;
  wire [0:0] h_arrdiv8_fs60_xor1;
  wire [0:0] h_arrdiv8_fs60_or0;
  wire [0:0] h_arrdiv8_fs61_xor1;
  wire [0:0] h_arrdiv8_fs61_or0;
  wire [0:0] h_arrdiv8_fs62_xor1;
  wire [0:0] h_arrdiv8_fs62_or0;
  wire [0:0] h_arrdiv8_fs63_xor1;
  wire [0:0] h_arrdiv8_fs63_or0;
  wire [0:0] h_arrdiv8_not7;

  fs fs_h_arrdiv8_fs0_out(.a(a[7]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv8_fs0_xor0), .fs_or0(h_arrdiv8_fs0_and0));
  fs fs_h_arrdiv8_fs1_out(.a(1'b0), .b(b[1]), .bin(h_arrdiv8_fs0_and0[0]), .fs_xor1(h_arrdiv8_fs1_xor1), .fs_or0(h_arrdiv8_fs1_or0));
  fs fs_h_arrdiv8_fs2_out(.a(1'b0), .b(b[2]), .bin(h_arrdiv8_fs1_or0[0]), .fs_xor1(h_arrdiv8_fs2_xor1), .fs_or0(h_arrdiv8_fs2_or0));
  fs fs_h_arrdiv8_fs3_out(.a(1'b0), .b(b[3]), .bin(h_arrdiv8_fs2_or0[0]), .fs_xor1(h_arrdiv8_fs3_xor1), .fs_or0(h_arrdiv8_fs3_or0));
  fs fs_h_arrdiv8_fs4_out(.a(1'b0), .b(b[4]), .bin(h_arrdiv8_fs3_or0[0]), .fs_xor1(h_arrdiv8_fs4_xor1), .fs_or0(h_arrdiv8_fs4_or0));
  fs fs_h_arrdiv8_fs5_out(.a(1'b0), .b(b[5]), .bin(h_arrdiv8_fs4_or0[0]), .fs_xor1(h_arrdiv8_fs5_xor1), .fs_or0(h_arrdiv8_fs5_or0));
  fs fs_h_arrdiv8_fs6_out(.a(1'b0), .b(b[6]), .bin(h_arrdiv8_fs5_or0[0]), .fs_xor1(h_arrdiv8_fs6_xor1), .fs_or0(h_arrdiv8_fs6_or0));
  fs fs_h_arrdiv8_fs7_out(.a(1'b0), .b(b[7]), .bin(h_arrdiv8_fs6_or0[0]), .fs_xor1(h_arrdiv8_fs7_xor1), .fs_or0(h_arrdiv8_fs7_or0));
  mux2to1 mux2to1_h_arrdiv8_mux2to10_out(.d0(h_arrdiv8_fs0_xor0[0]), .d1(a[7]), .sel(h_arrdiv8_fs7_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to10_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to11_out(.d0(h_arrdiv8_fs1_xor1[0]), .d1(1'b0), .sel(h_arrdiv8_fs7_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to11_and1));
  mux2to1 mux2to1_h_arrdiv8_mux2to12_out(.d0(h_arrdiv8_fs2_xor1[0]), .d1(1'b0), .sel(h_arrdiv8_fs7_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to12_and1));
  mux2to1 mux2to1_h_arrdiv8_mux2to13_out(.d0(h_arrdiv8_fs3_xor1[0]), .d1(1'b0), .sel(h_arrdiv8_fs7_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to13_and1));
  mux2to1 mux2to1_h_arrdiv8_mux2to14_out(.d0(h_arrdiv8_fs4_xor1[0]), .d1(1'b0), .sel(h_arrdiv8_fs7_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to14_and1));
  mux2to1 mux2to1_h_arrdiv8_mux2to15_out(.d0(h_arrdiv8_fs5_xor1[0]), .d1(1'b0), .sel(h_arrdiv8_fs7_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to15_and1));
  mux2to1 mux2to1_h_arrdiv8_mux2to16_out(.d0(h_arrdiv8_fs6_xor1[0]), .d1(1'b0), .sel(h_arrdiv8_fs7_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to16_and1));
  not_gate not_gate_h_arrdiv8_not0(.a(h_arrdiv8_fs7_or0[0]), .out(h_arrdiv8_not0));
  fs fs_h_arrdiv8_fs8_out(.a(a[6]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv8_fs8_xor0), .fs_or0(h_arrdiv8_fs8_and0));
  fs fs_h_arrdiv8_fs9_out(.a(h_arrdiv8_mux2to10_xor0[0]), .b(b[1]), .bin(h_arrdiv8_fs8_and0[0]), .fs_xor1(h_arrdiv8_fs9_xor1), .fs_or0(h_arrdiv8_fs9_or0));
  fs fs_h_arrdiv8_fs10_out(.a(h_arrdiv8_mux2to11_and1[0]), .b(b[2]), .bin(h_arrdiv8_fs9_or0[0]), .fs_xor1(h_arrdiv8_fs10_xor1), .fs_or0(h_arrdiv8_fs10_or0));
  fs fs_h_arrdiv8_fs11_out(.a(h_arrdiv8_mux2to12_and1[0]), .b(b[3]), .bin(h_arrdiv8_fs10_or0[0]), .fs_xor1(h_arrdiv8_fs11_xor1), .fs_or0(h_arrdiv8_fs11_or0));
  fs fs_h_arrdiv8_fs12_out(.a(h_arrdiv8_mux2to13_and1[0]), .b(b[4]), .bin(h_arrdiv8_fs11_or0[0]), .fs_xor1(h_arrdiv8_fs12_xor1), .fs_or0(h_arrdiv8_fs12_or0));
  fs fs_h_arrdiv8_fs13_out(.a(h_arrdiv8_mux2to14_and1[0]), .b(b[5]), .bin(h_arrdiv8_fs12_or0[0]), .fs_xor1(h_arrdiv8_fs13_xor1), .fs_or0(h_arrdiv8_fs13_or0));
  fs fs_h_arrdiv8_fs14_out(.a(h_arrdiv8_mux2to15_and1[0]), .b(b[6]), .bin(h_arrdiv8_fs13_or0[0]), .fs_xor1(h_arrdiv8_fs14_xor1), .fs_or0(h_arrdiv8_fs14_or0));
  fs fs_h_arrdiv8_fs15_out(.a(h_arrdiv8_mux2to16_and1[0]), .b(b[7]), .bin(h_arrdiv8_fs14_or0[0]), .fs_xor1(h_arrdiv8_fs15_xor1), .fs_or0(h_arrdiv8_fs15_or0));
  mux2to1 mux2to1_h_arrdiv8_mux2to17_out(.d0(h_arrdiv8_fs8_xor0[0]), .d1(a[6]), .sel(h_arrdiv8_fs15_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to17_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to18_out(.d0(h_arrdiv8_fs9_xor1[0]), .d1(h_arrdiv8_mux2to10_xor0[0]), .sel(h_arrdiv8_fs15_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to18_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to19_out(.d0(h_arrdiv8_fs10_xor1[0]), .d1(h_arrdiv8_mux2to11_and1[0]), .sel(h_arrdiv8_fs15_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to19_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to110_out(.d0(h_arrdiv8_fs11_xor1[0]), .d1(h_arrdiv8_mux2to12_and1[0]), .sel(h_arrdiv8_fs15_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to110_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to111_out(.d0(h_arrdiv8_fs12_xor1[0]), .d1(h_arrdiv8_mux2to13_and1[0]), .sel(h_arrdiv8_fs15_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to111_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to112_out(.d0(h_arrdiv8_fs13_xor1[0]), .d1(h_arrdiv8_mux2to14_and1[0]), .sel(h_arrdiv8_fs15_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to112_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to113_out(.d0(h_arrdiv8_fs14_xor1[0]), .d1(h_arrdiv8_mux2to15_and1[0]), .sel(h_arrdiv8_fs15_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to113_xor0));
  not_gate not_gate_h_arrdiv8_not1(.a(h_arrdiv8_fs15_or0[0]), .out(h_arrdiv8_not1));
  fs fs_h_arrdiv8_fs16_out(.a(a[5]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv8_fs16_xor0), .fs_or0(h_arrdiv8_fs16_and0));
  fs fs_h_arrdiv8_fs17_out(.a(h_arrdiv8_mux2to17_xor0[0]), .b(b[1]), .bin(h_arrdiv8_fs16_and0[0]), .fs_xor1(h_arrdiv8_fs17_xor1), .fs_or0(h_arrdiv8_fs17_or0));
  fs fs_h_arrdiv8_fs18_out(.a(h_arrdiv8_mux2to18_xor0[0]), .b(b[2]), .bin(h_arrdiv8_fs17_or0[0]), .fs_xor1(h_arrdiv8_fs18_xor1), .fs_or0(h_arrdiv8_fs18_or0));
  fs fs_h_arrdiv8_fs19_out(.a(h_arrdiv8_mux2to19_xor0[0]), .b(b[3]), .bin(h_arrdiv8_fs18_or0[0]), .fs_xor1(h_arrdiv8_fs19_xor1), .fs_or0(h_arrdiv8_fs19_or0));
  fs fs_h_arrdiv8_fs20_out(.a(h_arrdiv8_mux2to110_xor0[0]), .b(b[4]), .bin(h_arrdiv8_fs19_or0[0]), .fs_xor1(h_arrdiv8_fs20_xor1), .fs_or0(h_arrdiv8_fs20_or0));
  fs fs_h_arrdiv8_fs21_out(.a(h_arrdiv8_mux2to111_xor0[0]), .b(b[5]), .bin(h_arrdiv8_fs20_or0[0]), .fs_xor1(h_arrdiv8_fs21_xor1), .fs_or0(h_arrdiv8_fs21_or0));
  fs fs_h_arrdiv8_fs22_out(.a(h_arrdiv8_mux2to112_xor0[0]), .b(b[6]), .bin(h_arrdiv8_fs21_or0[0]), .fs_xor1(h_arrdiv8_fs22_xor1), .fs_or0(h_arrdiv8_fs22_or0));
  fs fs_h_arrdiv8_fs23_out(.a(h_arrdiv8_mux2to113_xor0[0]), .b(b[7]), .bin(h_arrdiv8_fs22_or0[0]), .fs_xor1(h_arrdiv8_fs23_xor1), .fs_or0(h_arrdiv8_fs23_or0));
  mux2to1 mux2to1_h_arrdiv8_mux2to114_out(.d0(h_arrdiv8_fs16_xor0[0]), .d1(a[5]), .sel(h_arrdiv8_fs23_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to114_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to115_out(.d0(h_arrdiv8_fs17_xor1[0]), .d1(h_arrdiv8_mux2to17_xor0[0]), .sel(h_arrdiv8_fs23_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to115_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to116_out(.d0(h_arrdiv8_fs18_xor1[0]), .d1(h_arrdiv8_mux2to18_xor0[0]), .sel(h_arrdiv8_fs23_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to116_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to117_out(.d0(h_arrdiv8_fs19_xor1[0]), .d1(h_arrdiv8_mux2to19_xor0[0]), .sel(h_arrdiv8_fs23_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to117_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to118_out(.d0(h_arrdiv8_fs20_xor1[0]), .d1(h_arrdiv8_mux2to110_xor0[0]), .sel(h_arrdiv8_fs23_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to118_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to119_out(.d0(h_arrdiv8_fs21_xor1[0]), .d1(h_arrdiv8_mux2to111_xor0[0]), .sel(h_arrdiv8_fs23_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to119_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to120_out(.d0(h_arrdiv8_fs22_xor1[0]), .d1(h_arrdiv8_mux2to112_xor0[0]), .sel(h_arrdiv8_fs23_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to120_xor0));
  not_gate not_gate_h_arrdiv8_not2(.a(h_arrdiv8_fs23_or0[0]), .out(h_arrdiv8_not2));
  fs fs_h_arrdiv8_fs24_out(.a(a[4]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv8_fs24_xor0), .fs_or0(h_arrdiv8_fs24_and0));
  fs fs_h_arrdiv8_fs25_out(.a(h_arrdiv8_mux2to114_xor0[0]), .b(b[1]), .bin(h_arrdiv8_fs24_and0[0]), .fs_xor1(h_arrdiv8_fs25_xor1), .fs_or0(h_arrdiv8_fs25_or0));
  fs fs_h_arrdiv8_fs26_out(.a(h_arrdiv8_mux2to115_xor0[0]), .b(b[2]), .bin(h_arrdiv8_fs25_or0[0]), .fs_xor1(h_arrdiv8_fs26_xor1), .fs_or0(h_arrdiv8_fs26_or0));
  fs fs_h_arrdiv8_fs27_out(.a(h_arrdiv8_mux2to116_xor0[0]), .b(b[3]), .bin(h_arrdiv8_fs26_or0[0]), .fs_xor1(h_arrdiv8_fs27_xor1), .fs_or0(h_arrdiv8_fs27_or0));
  fs fs_h_arrdiv8_fs28_out(.a(h_arrdiv8_mux2to117_xor0[0]), .b(b[4]), .bin(h_arrdiv8_fs27_or0[0]), .fs_xor1(h_arrdiv8_fs28_xor1), .fs_or0(h_arrdiv8_fs28_or0));
  fs fs_h_arrdiv8_fs29_out(.a(h_arrdiv8_mux2to118_xor0[0]), .b(b[5]), .bin(h_arrdiv8_fs28_or0[0]), .fs_xor1(h_arrdiv8_fs29_xor1), .fs_or0(h_arrdiv8_fs29_or0));
  fs fs_h_arrdiv8_fs30_out(.a(h_arrdiv8_mux2to119_xor0[0]), .b(b[6]), .bin(h_arrdiv8_fs29_or0[0]), .fs_xor1(h_arrdiv8_fs30_xor1), .fs_or0(h_arrdiv8_fs30_or0));
  fs fs_h_arrdiv8_fs31_out(.a(h_arrdiv8_mux2to120_xor0[0]), .b(b[7]), .bin(h_arrdiv8_fs30_or0[0]), .fs_xor1(h_arrdiv8_fs31_xor1), .fs_or0(h_arrdiv8_fs31_or0));
  mux2to1 mux2to1_h_arrdiv8_mux2to121_out(.d0(h_arrdiv8_fs24_xor0[0]), .d1(a[4]), .sel(h_arrdiv8_fs31_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to121_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to122_out(.d0(h_arrdiv8_fs25_xor1[0]), .d1(h_arrdiv8_mux2to114_xor0[0]), .sel(h_arrdiv8_fs31_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to122_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to123_out(.d0(h_arrdiv8_fs26_xor1[0]), .d1(h_arrdiv8_mux2to115_xor0[0]), .sel(h_arrdiv8_fs31_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to123_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to124_out(.d0(h_arrdiv8_fs27_xor1[0]), .d1(h_arrdiv8_mux2to116_xor0[0]), .sel(h_arrdiv8_fs31_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to124_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to125_out(.d0(h_arrdiv8_fs28_xor1[0]), .d1(h_arrdiv8_mux2to117_xor0[0]), .sel(h_arrdiv8_fs31_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to125_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to126_out(.d0(h_arrdiv8_fs29_xor1[0]), .d1(h_arrdiv8_mux2to118_xor0[0]), .sel(h_arrdiv8_fs31_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to126_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to127_out(.d0(h_arrdiv8_fs30_xor1[0]), .d1(h_arrdiv8_mux2to119_xor0[0]), .sel(h_arrdiv8_fs31_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to127_xor0));
  not_gate not_gate_h_arrdiv8_not3(.a(h_arrdiv8_fs31_or0[0]), .out(h_arrdiv8_not3));
  fs fs_h_arrdiv8_fs32_out(.a(a[3]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv8_fs32_xor0), .fs_or0(h_arrdiv8_fs32_and0));
  fs fs_h_arrdiv8_fs33_out(.a(h_arrdiv8_mux2to121_xor0[0]), .b(b[1]), .bin(h_arrdiv8_fs32_and0[0]), .fs_xor1(h_arrdiv8_fs33_xor1), .fs_or0(h_arrdiv8_fs33_or0));
  fs fs_h_arrdiv8_fs34_out(.a(h_arrdiv8_mux2to122_xor0[0]), .b(b[2]), .bin(h_arrdiv8_fs33_or0[0]), .fs_xor1(h_arrdiv8_fs34_xor1), .fs_or0(h_arrdiv8_fs34_or0));
  fs fs_h_arrdiv8_fs35_out(.a(h_arrdiv8_mux2to123_xor0[0]), .b(b[3]), .bin(h_arrdiv8_fs34_or0[0]), .fs_xor1(h_arrdiv8_fs35_xor1), .fs_or0(h_arrdiv8_fs35_or0));
  fs fs_h_arrdiv8_fs36_out(.a(h_arrdiv8_mux2to124_xor0[0]), .b(b[4]), .bin(h_arrdiv8_fs35_or0[0]), .fs_xor1(h_arrdiv8_fs36_xor1), .fs_or0(h_arrdiv8_fs36_or0));
  fs fs_h_arrdiv8_fs37_out(.a(h_arrdiv8_mux2to125_xor0[0]), .b(b[5]), .bin(h_arrdiv8_fs36_or0[0]), .fs_xor1(h_arrdiv8_fs37_xor1), .fs_or0(h_arrdiv8_fs37_or0));
  fs fs_h_arrdiv8_fs38_out(.a(h_arrdiv8_mux2to126_xor0[0]), .b(b[6]), .bin(h_arrdiv8_fs37_or0[0]), .fs_xor1(h_arrdiv8_fs38_xor1), .fs_or0(h_arrdiv8_fs38_or0));
  fs fs_h_arrdiv8_fs39_out(.a(h_arrdiv8_mux2to127_xor0[0]), .b(b[7]), .bin(h_arrdiv8_fs38_or0[0]), .fs_xor1(h_arrdiv8_fs39_xor1), .fs_or0(h_arrdiv8_fs39_or0));
  mux2to1 mux2to1_h_arrdiv8_mux2to128_out(.d0(h_arrdiv8_fs32_xor0[0]), .d1(a[3]), .sel(h_arrdiv8_fs39_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to128_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to129_out(.d0(h_arrdiv8_fs33_xor1[0]), .d1(h_arrdiv8_mux2to121_xor0[0]), .sel(h_arrdiv8_fs39_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to129_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to130_out(.d0(h_arrdiv8_fs34_xor1[0]), .d1(h_arrdiv8_mux2to122_xor0[0]), .sel(h_arrdiv8_fs39_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to130_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to131_out(.d0(h_arrdiv8_fs35_xor1[0]), .d1(h_arrdiv8_mux2to123_xor0[0]), .sel(h_arrdiv8_fs39_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to131_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to132_out(.d0(h_arrdiv8_fs36_xor1[0]), .d1(h_arrdiv8_mux2to124_xor0[0]), .sel(h_arrdiv8_fs39_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to132_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to133_out(.d0(h_arrdiv8_fs37_xor1[0]), .d1(h_arrdiv8_mux2to125_xor0[0]), .sel(h_arrdiv8_fs39_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to133_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to134_out(.d0(h_arrdiv8_fs38_xor1[0]), .d1(h_arrdiv8_mux2to126_xor0[0]), .sel(h_arrdiv8_fs39_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to134_xor0));
  not_gate not_gate_h_arrdiv8_not4(.a(h_arrdiv8_fs39_or0[0]), .out(h_arrdiv8_not4));
  fs fs_h_arrdiv8_fs40_out(.a(a[2]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv8_fs40_xor0), .fs_or0(h_arrdiv8_fs40_and0));
  fs fs_h_arrdiv8_fs41_out(.a(h_arrdiv8_mux2to128_xor0[0]), .b(b[1]), .bin(h_arrdiv8_fs40_and0[0]), .fs_xor1(h_arrdiv8_fs41_xor1), .fs_or0(h_arrdiv8_fs41_or0));
  fs fs_h_arrdiv8_fs42_out(.a(h_arrdiv8_mux2to129_xor0[0]), .b(b[2]), .bin(h_arrdiv8_fs41_or0[0]), .fs_xor1(h_arrdiv8_fs42_xor1), .fs_or0(h_arrdiv8_fs42_or0));
  fs fs_h_arrdiv8_fs43_out(.a(h_arrdiv8_mux2to130_xor0[0]), .b(b[3]), .bin(h_arrdiv8_fs42_or0[0]), .fs_xor1(h_arrdiv8_fs43_xor1), .fs_or0(h_arrdiv8_fs43_or0));
  fs fs_h_arrdiv8_fs44_out(.a(h_arrdiv8_mux2to131_xor0[0]), .b(b[4]), .bin(h_arrdiv8_fs43_or0[0]), .fs_xor1(h_arrdiv8_fs44_xor1), .fs_or0(h_arrdiv8_fs44_or0));
  fs fs_h_arrdiv8_fs45_out(.a(h_arrdiv8_mux2to132_xor0[0]), .b(b[5]), .bin(h_arrdiv8_fs44_or0[0]), .fs_xor1(h_arrdiv8_fs45_xor1), .fs_or0(h_arrdiv8_fs45_or0));
  fs fs_h_arrdiv8_fs46_out(.a(h_arrdiv8_mux2to133_xor0[0]), .b(b[6]), .bin(h_arrdiv8_fs45_or0[0]), .fs_xor1(h_arrdiv8_fs46_xor1), .fs_or0(h_arrdiv8_fs46_or0));
  fs fs_h_arrdiv8_fs47_out(.a(h_arrdiv8_mux2to134_xor0[0]), .b(b[7]), .bin(h_arrdiv8_fs46_or0[0]), .fs_xor1(h_arrdiv8_fs47_xor1), .fs_or0(h_arrdiv8_fs47_or0));
  mux2to1 mux2to1_h_arrdiv8_mux2to135_out(.d0(h_arrdiv8_fs40_xor0[0]), .d1(a[2]), .sel(h_arrdiv8_fs47_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to135_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to136_out(.d0(h_arrdiv8_fs41_xor1[0]), .d1(h_arrdiv8_mux2to128_xor0[0]), .sel(h_arrdiv8_fs47_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to136_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to137_out(.d0(h_arrdiv8_fs42_xor1[0]), .d1(h_arrdiv8_mux2to129_xor0[0]), .sel(h_arrdiv8_fs47_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to137_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to138_out(.d0(h_arrdiv8_fs43_xor1[0]), .d1(h_arrdiv8_mux2to130_xor0[0]), .sel(h_arrdiv8_fs47_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to138_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to139_out(.d0(h_arrdiv8_fs44_xor1[0]), .d1(h_arrdiv8_mux2to131_xor0[0]), .sel(h_arrdiv8_fs47_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to139_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to140_out(.d0(h_arrdiv8_fs45_xor1[0]), .d1(h_arrdiv8_mux2to132_xor0[0]), .sel(h_arrdiv8_fs47_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to140_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to141_out(.d0(h_arrdiv8_fs46_xor1[0]), .d1(h_arrdiv8_mux2to133_xor0[0]), .sel(h_arrdiv8_fs47_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to141_xor0));
  not_gate not_gate_h_arrdiv8_not5(.a(h_arrdiv8_fs47_or0[0]), .out(h_arrdiv8_not5));
  fs fs_h_arrdiv8_fs48_out(.a(a[1]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv8_fs48_xor0), .fs_or0(h_arrdiv8_fs48_and0));
  fs fs_h_arrdiv8_fs49_out(.a(h_arrdiv8_mux2to135_xor0[0]), .b(b[1]), .bin(h_arrdiv8_fs48_and0[0]), .fs_xor1(h_arrdiv8_fs49_xor1), .fs_or0(h_arrdiv8_fs49_or0));
  fs fs_h_arrdiv8_fs50_out(.a(h_arrdiv8_mux2to136_xor0[0]), .b(b[2]), .bin(h_arrdiv8_fs49_or0[0]), .fs_xor1(h_arrdiv8_fs50_xor1), .fs_or0(h_arrdiv8_fs50_or0));
  fs fs_h_arrdiv8_fs51_out(.a(h_arrdiv8_mux2to137_xor0[0]), .b(b[3]), .bin(h_arrdiv8_fs50_or0[0]), .fs_xor1(h_arrdiv8_fs51_xor1), .fs_or0(h_arrdiv8_fs51_or0));
  fs fs_h_arrdiv8_fs52_out(.a(h_arrdiv8_mux2to138_xor0[0]), .b(b[4]), .bin(h_arrdiv8_fs51_or0[0]), .fs_xor1(h_arrdiv8_fs52_xor1), .fs_or0(h_arrdiv8_fs52_or0));
  fs fs_h_arrdiv8_fs53_out(.a(h_arrdiv8_mux2to139_xor0[0]), .b(b[5]), .bin(h_arrdiv8_fs52_or0[0]), .fs_xor1(h_arrdiv8_fs53_xor1), .fs_or0(h_arrdiv8_fs53_or0));
  fs fs_h_arrdiv8_fs54_out(.a(h_arrdiv8_mux2to140_xor0[0]), .b(b[6]), .bin(h_arrdiv8_fs53_or0[0]), .fs_xor1(h_arrdiv8_fs54_xor1), .fs_or0(h_arrdiv8_fs54_or0));
  fs fs_h_arrdiv8_fs55_out(.a(h_arrdiv8_mux2to141_xor0[0]), .b(b[7]), .bin(h_arrdiv8_fs54_or0[0]), .fs_xor1(h_arrdiv8_fs55_xor1), .fs_or0(h_arrdiv8_fs55_or0));
  mux2to1 mux2to1_h_arrdiv8_mux2to142_out(.d0(h_arrdiv8_fs48_xor0[0]), .d1(a[1]), .sel(h_arrdiv8_fs55_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to142_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to143_out(.d0(h_arrdiv8_fs49_xor1[0]), .d1(h_arrdiv8_mux2to135_xor0[0]), .sel(h_arrdiv8_fs55_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to143_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to144_out(.d0(h_arrdiv8_fs50_xor1[0]), .d1(h_arrdiv8_mux2to136_xor0[0]), .sel(h_arrdiv8_fs55_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to144_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to145_out(.d0(h_arrdiv8_fs51_xor1[0]), .d1(h_arrdiv8_mux2to137_xor0[0]), .sel(h_arrdiv8_fs55_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to145_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to146_out(.d0(h_arrdiv8_fs52_xor1[0]), .d1(h_arrdiv8_mux2to138_xor0[0]), .sel(h_arrdiv8_fs55_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to146_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to147_out(.d0(h_arrdiv8_fs53_xor1[0]), .d1(h_arrdiv8_mux2to139_xor0[0]), .sel(h_arrdiv8_fs55_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to147_xor0));
  mux2to1 mux2to1_h_arrdiv8_mux2to148_out(.d0(h_arrdiv8_fs54_xor1[0]), .d1(h_arrdiv8_mux2to140_xor0[0]), .sel(h_arrdiv8_fs55_or0[0]), .mux2to1_xor0(h_arrdiv8_mux2to148_xor0));
  not_gate not_gate_h_arrdiv8_not6(.a(h_arrdiv8_fs55_or0[0]), .out(h_arrdiv8_not6));
  fs fs_h_arrdiv8_fs56_out(.a(a[0]), .b(b[0]), .bin(1'b0), .fs_xor1(h_arrdiv8_fs56_xor0), .fs_or0(h_arrdiv8_fs56_and0));
  fs fs_h_arrdiv8_fs57_out(.a(h_arrdiv8_mux2to142_xor0[0]), .b(b[1]), .bin(h_arrdiv8_fs56_and0[0]), .fs_xor1(h_arrdiv8_fs57_xor1), .fs_or0(h_arrdiv8_fs57_or0));
  fs fs_h_arrdiv8_fs58_out(.a(h_arrdiv8_mux2to143_xor0[0]), .b(b[2]), .bin(h_arrdiv8_fs57_or0[0]), .fs_xor1(h_arrdiv8_fs58_xor1), .fs_or0(h_arrdiv8_fs58_or0));
  fs fs_h_arrdiv8_fs59_out(.a(h_arrdiv8_mux2to144_xor0[0]), .b(b[3]), .bin(h_arrdiv8_fs58_or0[0]), .fs_xor1(h_arrdiv8_fs59_xor1), .fs_or0(h_arrdiv8_fs59_or0));
  fs fs_h_arrdiv8_fs60_out(.a(h_arrdiv8_mux2to145_xor0[0]), .b(b[4]), .bin(h_arrdiv8_fs59_or0[0]), .fs_xor1(h_arrdiv8_fs60_xor1), .fs_or0(h_arrdiv8_fs60_or0));
  fs fs_h_arrdiv8_fs61_out(.a(h_arrdiv8_mux2to146_xor0[0]), .b(b[5]), .bin(h_arrdiv8_fs60_or0[0]), .fs_xor1(h_arrdiv8_fs61_xor1), .fs_or0(h_arrdiv8_fs61_or0));
  fs fs_h_arrdiv8_fs62_out(.a(h_arrdiv8_mux2to147_xor0[0]), .b(b[6]), .bin(h_arrdiv8_fs61_or0[0]), .fs_xor1(h_arrdiv8_fs62_xor1), .fs_or0(h_arrdiv8_fs62_or0));
  fs fs_h_arrdiv8_fs63_out(.a(h_arrdiv8_mux2to148_xor0[0]), .b(b[7]), .bin(h_arrdiv8_fs62_or0[0]), .fs_xor1(h_arrdiv8_fs63_xor1), .fs_or0(h_arrdiv8_fs63_or0));
  not_gate not_gate_h_arrdiv8_not7(.a(h_arrdiv8_fs63_or0[0]), .out(h_arrdiv8_not7));

  assign h_arrdiv8_out[0] = h_arrdiv8_not7[0];
  assign h_arrdiv8_out[1] = h_arrdiv8_not6[0];
  assign h_arrdiv8_out[2] = h_arrdiv8_not5[0];
  assign h_arrdiv8_out[3] = h_arrdiv8_not4[0];
  assign h_arrdiv8_out[4] = h_arrdiv8_not3[0];
  assign h_arrdiv8_out[5] = h_arrdiv8_not2[0];
  assign h_arrdiv8_out[6] = h_arrdiv8_not1[0];
  assign h_arrdiv8_out[7] = h_arrdiv8_not0[0];
endmodule