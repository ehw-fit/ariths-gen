module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(a[0], b[0], pg_logic_or0);
  and_gate and_gate_pg_logic_and0(a[0], b[0], pg_logic_and0);
  xor_gate xor_gate_pg_logic_xor0(a[0], b[0], pg_logic_xor0);
endmodule

module h_s_cla12(input [11:0] a, input [11:0] b, output [12:0] h_s_cla12_out);
  wire [0:0] h_s_cla12_pg_logic0_or0;
  wire [0:0] h_s_cla12_pg_logic0_and0;
  wire [0:0] h_s_cla12_pg_logic0_xor0;
  wire [0:0] h_s_cla12_pg_logic1_or0;
  wire [0:0] h_s_cla12_pg_logic1_and0;
  wire [0:0] h_s_cla12_pg_logic1_xor0;
  wire [0:0] h_s_cla12_xor1;
  wire [0:0] h_s_cla12_and0;
  wire [0:0] h_s_cla12_or0;
  wire [0:0] h_s_cla12_pg_logic2_or0;
  wire [0:0] h_s_cla12_pg_logic2_and0;
  wire [0:0] h_s_cla12_pg_logic2_xor0;
  wire [0:0] h_s_cla12_xor2;
  wire [0:0] h_s_cla12_and1;
  wire [0:0] h_s_cla12_and2;
  wire [0:0] h_s_cla12_and3;
  wire [0:0] h_s_cla12_and4;
  wire [0:0] h_s_cla12_or1;
  wire [0:0] h_s_cla12_or2;
  wire [0:0] h_s_cla12_pg_logic3_or0;
  wire [0:0] h_s_cla12_pg_logic3_and0;
  wire [0:0] h_s_cla12_pg_logic3_xor0;
  wire [0:0] h_s_cla12_xor3;
  wire [0:0] h_s_cla12_and5;
  wire [0:0] h_s_cla12_and6;
  wire [0:0] h_s_cla12_and7;
  wire [0:0] h_s_cla12_and8;
  wire [0:0] h_s_cla12_and9;
  wire [0:0] h_s_cla12_and10;
  wire [0:0] h_s_cla12_and11;
  wire [0:0] h_s_cla12_or3;
  wire [0:0] h_s_cla12_or4;
  wire [0:0] h_s_cla12_or5;
  wire [0:0] h_s_cla12_pg_logic4_or0;
  wire [0:0] h_s_cla12_pg_logic4_and0;
  wire [0:0] h_s_cla12_pg_logic4_xor0;
  wire [0:0] h_s_cla12_xor4;
  wire [0:0] h_s_cla12_and12;
  wire [0:0] h_s_cla12_or6;
  wire [0:0] h_s_cla12_pg_logic5_or0;
  wire [0:0] h_s_cla12_pg_logic5_and0;
  wire [0:0] h_s_cla12_pg_logic5_xor0;
  wire [0:0] h_s_cla12_xor5;
  wire [0:0] h_s_cla12_and13;
  wire [0:0] h_s_cla12_and14;
  wire [0:0] h_s_cla12_and15;
  wire [0:0] h_s_cla12_or7;
  wire [0:0] h_s_cla12_or8;
  wire [0:0] h_s_cla12_pg_logic6_or0;
  wire [0:0] h_s_cla12_pg_logic6_and0;
  wire [0:0] h_s_cla12_pg_logic6_xor0;
  wire [0:0] h_s_cla12_xor6;
  wire [0:0] h_s_cla12_and16;
  wire [0:0] h_s_cla12_and17;
  wire [0:0] h_s_cla12_and18;
  wire [0:0] h_s_cla12_and19;
  wire [0:0] h_s_cla12_and20;
  wire [0:0] h_s_cla12_and21;
  wire [0:0] h_s_cla12_or9;
  wire [0:0] h_s_cla12_or10;
  wire [0:0] h_s_cla12_or11;
  wire [0:0] h_s_cla12_pg_logic7_or0;
  wire [0:0] h_s_cla12_pg_logic7_and0;
  wire [0:0] h_s_cla12_pg_logic7_xor0;
  wire [0:0] h_s_cla12_xor7;
  wire [0:0] h_s_cla12_and22;
  wire [0:0] h_s_cla12_and23;
  wire [0:0] h_s_cla12_and24;
  wire [0:0] h_s_cla12_and25;
  wire [0:0] h_s_cla12_and26;
  wire [0:0] h_s_cla12_and27;
  wire [0:0] h_s_cla12_and28;
  wire [0:0] h_s_cla12_and29;
  wire [0:0] h_s_cla12_and30;
  wire [0:0] h_s_cla12_and31;
  wire [0:0] h_s_cla12_or12;
  wire [0:0] h_s_cla12_or13;
  wire [0:0] h_s_cla12_or14;
  wire [0:0] h_s_cla12_or15;
  wire [0:0] h_s_cla12_pg_logic8_or0;
  wire [0:0] h_s_cla12_pg_logic8_and0;
  wire [0:0] h_s_cla12_pg_logic8_xor0;
  wire [0:0] h_s_cla12_xor8;
  wire [0:0] h_s_cla12_and32;
  wire [0:0] h_s_cla12_or16;
  wire [0:0] h_s_cla12_pg_logic9_or0;
  wire [0:0] h_s_cla12_pg_logic9_and0;
  wire [0:0] h_s_cla12_pg_logic9_xor0;
  wire [0:0] h_s_cla12_xor9;
  wire [0:0] h_s_cla12_and33;
  wire [0:0] h_s_cla12_and34;
  wire [0:0] h_s_cla12_and35;
  wire [0:0] h_s_cla12_or17;
  wire [0:0] h_s_cla12_or18;
  wire [0:0] h_s_cla12_pg_logic10_or0;
  wire [0:0] h_s_cla12_pg_logic10_and0;
  wire [0:0] h_s_cla12_pg_logic10_xor0;
  wire [0:0] h_s_cla12_xor10;
  wire [0:0] h_s_cla12_and36;
  wire [0:0] h_s_cla12_and37;
  wire [0:0] h_s_cla12_and38;
  wire [0:0] h_s_cla12_and39;
  wire [0:0] h_s_cla12_and40;
  wire [0:0] h_s_cla12_and41;
  wire [0:0] h_s_cla12_or19;
  wire [0:0] h_s_cla12_or20;
  wire [0:0] h_s_cla12_or21;
  wire [0:0] h_s_cla12_pg_logic11_or0;
  wire [0:0] h_s_cla12_pg_logic11_and0;
  wire [0:0] h_s_cla12_pg_logic11_xor0;
  wire [0:0] h_s_cla12_xor11;
  wire [0:0] h_s_cla12_and42;
  wire [0:0] h_s_cla12_and43;
  wire [0:0] h_s_cla12_and44;
  wire [0:0] h_s_cla12_and45;
  wire [0:0] h_s_cla12_and46;
  wire [0:0] h_s_cla12_and47;
  wire [0:0] h_s_cla12_and48;
  wire [0:0] h_s_cla12_and49;
  wire [0:0] h_s_cla12_and50;
  wire [0:0] h_s_cla12_and51;
  wire [0:0] h_s_cla12_or22;
  wire [0:0] h_s_cla12_or23;
  wire [0:0] h_s_cla12_or24;
  wire [0:0] h_s_cla12_or25;
  wire [0:0] h_s_cla12_xor12;
  wire [0:0] h_s_cla12_xor13;

  pg_logic pg_logic_h_s_cla12_pg_logic0_out(a[0], b[0], h_s_cla12_pg_logic0_or0, h_s_cla12_pg_logic0_and0, h_s_cla12_pg_logic0_xor0);
  pg_logic pg_logic_h_s_cla12_pg_logic1_out(a[1], b[1], h_s_cla12_pg_logic1_or0, h_s_cla12_pg_logic1_and0, h_s_cla12_pg_logic1_xor0);
  xor_gate xor_gate_h_s_cla12_xor1(h_s_cla12_pg_logic1_xor0[0], h_s_cla12_pg_logic0_and0[0], h_s_cla12_xor1);
  and_gate and_gate_h_s_cla12_and0(h_s_cla12_pg_logic0_and0[0], h_s_cla12_pg_logic1_or0[0], h_s_cla12_and0);
  or_gate or_gate_h_s_cla12_or0(h_s_cla12_pg_logic1_and0[0], h_s_cla12_and0[0], h_s_cla12_or0);
  pg_logic pg_logic_h_s_cla12_pg_logic2_out(a[2], b[2], h_s_cla12_pg_logic2_or0, h_s_cla12_pg_logic2_and0, h_s_cla12_pg_logic2_xor0);
  xor_gate xor_gate_h_s_cla12_xor2(h_s_cla12_pg_logic2_xor0[0], h_s_cla12_or0[0], h_s_cla12_xor2);
  and_gate and_gate_h_s_cla12_and1(h_s_cla12_pg_logic2_or0[0], h_s_cla12_pg_logic0_or0[0], h_s_cla12_and1);
  and_gate and_gate_h_s_cla12_and2(h_s_cla12_pg_logic0_and0[0], h_s_cla12_pg_logic2_or0[0], h_s_cla12_and2);
  and_gate and_gate_h_s_cla12_and3(h_s_cla12_and2[0], h_s_cla12_pg_logic1_or0[0], h_s_cla12_and3);
  and_gate and_gate_h_s_cla12_and4(h_s_cla12_pg_logic1_and0[0], h_s_cla12_pg_logic2_or0[0], h_s_cla12_and4);
  or_gate or_gate_h_s_cla12_or1(h_s_cla12_and3[0], h_s_cla12_and4[0], h_s_cla12_or1);
  or_gate or_gate_h_s_cla12_or2(h_s_cla12_pg_logic2_and0[0], h_s_cla12_or1[0], h_s_cla12_or2);
  pg_logic pg_logic_h_s_cla12_pg_logic3_out(a[3], b[3], h_s_cla12_pg_logic3_or0, h_s_cla12_pg_logic3_and0, h_s_cla12_pg_logic3_xor0);
  xor_gate xor_gate_h_s_cla12_xor3(h_s_cla12_pg_logic3_xor0[0], h_s_cla12_or2[0], h_s_cla12_xor3);
  and_gate and_gate_h_s_cla12_and5(h_s_cla12_pg_logic3_or0[0], h_s_cla12_pg_logic1_or0[0], h_s_cla12_and5);
  and_gate and_gate_h_s_cla12_and6(h_s_cla12_pg_logic0_and0[0], h_s_cla12_pg_logic2_or0[0], h_s_cla12_and6);
  and_gate and_gate_h_s_cla12_and7(h_s_cla12_pg_logic3_or0[0], h_s_cla12_pg_logic1_or0[0], h_s_cla12_and7);
  and_gate and_gate_h_s_cla12_and8(h_s_cla12_and6[0], h_s_cla12_and7[0], h_s_cla12_and8);
  and_gate and_gate_h_s_cla12_and9(h_s_cla12_pg_logic1_and0[0], h_s_cla12_pg_logic3_or0[0], h_s_cla12_and9);
  and_gate and_gate_h_s_cla12_and10(h_s_cla12_and9[0], h_s_cla12_pg_logic2_or0[0], h_s_cla12_and10);
  and_gate and_gate_h_s_cla12_and11(h_s_cla12_pg_logic2_and0[0], h_s_cla12_pg_logic3_or0[0], h_s_cla12_and11);
  or_gate or_gate_h_s_cla12_or3(h_s_cla12_and8[0], h_s_cla12_and11[0], h_s_cla12_or3);
  or_gate or_gate_h_s_cla12_or4(h_s_cla12_and10[0], h_s_cla12_or3[0], h_s_cla12_or4);
  or_gate or_gate_h_s_cla12_or5(h_s_cla12_pg_logic3_and0[0], h_s_cla12_or4[0], h_s_cla12_or5);
  pg_logic pg_logic_h_s_cla12_pg_logic4_out(a[4], b[4], h_s_cla12_pg_logic4_or0, h_s_cla12_pg_logic4_and0, h_s_cla12_pg_logic4_xor0);
  xor_gate xor_gate_h_s_cla12_xor4(h_s_cla12_pg_logic4_xor0[0], h_s_cla12_or5[0], h_s_cla12_xor4);
  and_gate and_gate_h_s_cla12_and12(h_s_cla12_or5[0], h_s_cla12_pg_logic4_or0[0], h_s_cla12_and12);
  or_gate or_gate_h_s_cla12_or6(h_s_cla12_pg_logic4_and0[0], h_s_cla12_and12[0], h_s_cla12_or6);
  pg_logic pg_logic_h_s_cla12_pg_logic5_out(a[5], b[5], h_s_cla12_pg_logic5_or0, h_s_cla12_pg_logic5_and0, h_s_cla12_pg_logic5_xor0);
  xor_gate xor_gate_h_s_cla12_xor5(h_s_cla12_pg_logic5_xor0[0], h_s_cla12_or6[0], h_s_cla12_xor5);
  and_gate and_gate_h_s_cla12_and13(h_s_cla12_or5[0], h_s_cla12_pg_logic5_or0[0], h_s_cla12_and13);
  and_gate and_gate_h_s_cla12_and14(h_s_cla12_and13[0], h_s_cla12_pg_logic4_or0[0], h_s_cla12_and14);
  and_gate and_gate_h_s_cla12_and15(h_s_cla12_pg_logic4_and0[0], h_s_cla12_pg_logic5_or0[0], h_s_cla12_and15);
  or_gate or_gate_h_s_cla12_or7(h_s_cla12_and14[0], h_s_cla12_and15[0], h_s_cla12_or7);
  or_gate or_gate_h_s_cla12_or8(h_s_cla12_pg_logic5_and0[0], h_s_cla12_or7[0], h_s_cla12_or8);
  pg_logic pg_logic_h_s_cla12_pg_logic6_out(a[6], b[6], h_s_cla12_pg_logic6_or0, h_s_cla12_pg_logic6_and0, h_s_cla12_pg_logic6_xor0);
  xor_gate xor_gate_h_s_cla12_xor6(h_s_cla12_pg_logic6_xor0[0], h_s_cla12_or8[0], h_s_cla12_xor6);
  and_gate and_gate_h_s_cla12_and16(h_s_cla12_or5[0], h_s_cla12_pg_logic5_or0[0], h_s_cla12_and16);
  and_gate and_gate_h_s_cla12_and17(h_s_cla12_pg_logic6_or0[0], h_s_cla12_pg_logic4_or0[0], h_s_cla12_and17);
  and_gate and_gate_h_s_cla12_and18(h_s_cla12_and16[0], h_s_cla12_and17[0], h_s_cla12_and18);
  and_gate and_gate_h_s_cla12_and19(h_s_cla12_pg_logic4_and0[0], h_s_cla12_pg_logic6_or0[0], h_s_cla12_and19);
  and_gate and_gate_h_s_cla12_and20(h_s_cla12_and19[0], h_s_cla12_pg_logic5_or0[0], h_s_cla12_and20);
  and_gate and_gate_h_s_cla12_and21(h_s_cla12_pg_logic5_and0[0], h_s_cla12_pg_logic6_or0[0], h_s_cla12_and21);
  or_gate or_gate_h_s_cla12_or9(h_s_cla12_and18[0], h_s_cla12_and20[0], h_s_cla12_or9);
  or_gate or_gate_h_s_cla12_or10(h_s_cla12_or9[0], h_s_cla12_and21[0], h_s_cla12_or10);
  or_gate or_gate_h_s_cla12_or11(h_s_cla12_pg_logic6_and0[0], h_s_cla12_or10[0], h_s_cla12_or11);
  pg_logic pg_logic_h_s_cla12_pg_logic7_out(a[7], b[7], h_s_cla12_pg_logic7_or0, h_s_cla12_pg_logic7_and0, h_s_cla12_pg_logic7_xor0);
  xor_gate xor_gate_h_s_cla12_xor7(h_s_cla12_pg_logic7_xor0[0], h_s_cla12_or11[0], h_s_cla12_xor7);
  and_gate and_gate_h_s_cla12_and22(h_s_cla12_or5[0], h_s_cla12_pg_logic6_or0[0], h_s_cla12_and22);
  and_gate and_gate_h_s_cla12_and23(h_s_cla12_pg_logic7_or0[0], h_s_cla12_pg_logic5_or0[0], h_s_cla12_and23);
  and_gate and_gate_h_s_cla12_and24(h_s_cla12_and22[0], h_s_cla12_and23[0], h_s_cla12_and24);
  and_gate and_gate_h_s_cla12_and25(h_s_cla12_and24[0], h_s_cla12_pg_logic4_or0[0], h_s_cla12_and25);
  and_gate and_gate_h_s_cla12_and26(h_s_cla12_pg_logic4_and0[0], h_s_cla12_pg_logic6_or0[0], h_s_cla12_and26);
  and_gate and_gate_h_s_cla12_and27(h_s_cla12_pg_logic7_or0[0], h_s_cla12_pg_logic5_or0[0], h_s_cla12_and27);
  and_gate and_gate_h_s_cla12_and28(h_s_cla12_and26[0], h_s_cla12_and27[0], h_s_cla12_and28);
  and_gate and_gate_h_s_cla12_and29(h_s_cla12_pg_logic5_and0[0], h_s_cla12_pg_logic7_or0[0], h_s_cla12_and29);
  and_gate and_gate_h_s_cla12_and30(h_s_cla12_and29[0], h_s_cla12_pg_logic6_or0[0], h_s_cla12_and30);
  and_gate and_gate_h_s_cla12_and31(h_s_cla12_pg_logic6_and0[0], h_s_cla12_pg_logic7_or0[0], h_s_cla12_and31);
  or_gate or_gate_h_s_cla12_or12(h_s_cla12_and25[0], h_s_cla12_and30[0], h_s_cla12_or12);
  or_gate or_gate_h_s_cla12_or13(h_s_cla12_and28[0], h_s_cla12_and31[0], h_s_cla12_or13);
  or_gate or_gate_h_s_cla12_or14(h_s_cla12_or12[0], h_s_cla12_or13[0], h_s_cla12_or14);
  or_gate or_gate_h_s_cla12_or15(h_s_cla12_pg_logic7_and0[0], h_s_cla12_or14[0], h_s_cla12_or15);
  pg_logic pg_logic_h_s_cla12_pg_logic8_out(a[8], b[8], h_s_cla12_pg_logic8_or0, h_s_cla12_pg_logic8_and0, h_s_cla12_pg_logic8_xor0);
  xor_gate xor_gate_h_s_cla12_xor8(h_s_cla12_pg_logic8_xor0[0], h_s_cla12_or15[0], h_s_cla12_xor8);
  and_gate and_gate_h_s_cla12_and32(h_s_cla12_or15[0], h_s_cla12_pg_logic8_or0[0], h_s_cla12_and32);
  or_gate or_gate_h_s_cla12_or16(h_s_cla12_pg_logic8_and0[0], h_s_cla12_and32[0], h_s_cla12_or16);
  pg_logic pg_logic_h_s_cla12_pg_logic9_out(a[9], b[9], h_s_cla12_pg_logic9_or0, h_s_cla12_pg_logic9_and0, h_s_cla12_pg_logic9_xor0);
  xor_gate xor_gate_h_s_cla12_xor9(h_s_cla12_pg_logic9_xor0[0], h_s_cla12_or16[0], h_s_cla12_xor9);
  and_gate and_gate_h_s_cla12_and33(h_s_cla12_or15[0], h_s_cla12_pg_logic9_or0[0], h_s_cla12_and33);
  and_gate and_gate_h_s_cla12_and34(h_s_cla12_and33[0], h_s_cla12_pg_logic8_or0[0], h_s_cla12_and34);
  and_gate and_gate_h_s_cla12_and35(h_s_cla12_pg_logic8_and0[0], h_s_cla12_pg_logic9_or0[0], h_s_cla12_and35);
  or_gate or_gate_h_s_cla12_or17(h_s_cla12_and34[0], h_s_cla12_and35[0], h_s_cla12_or17);
  or_gate or_gate_h_s_cla12_or18(h_s_cla12_pg_logic9_and0[0], h_s_cla12_or17[0], h_s_cla12_or18);
  pg_logic pg_logic_h_s_cla12_pg_logic10_out(a[10], b[10], h_s_cla12_pg_logic10_or0, h_s_cla12_pg_logic10_and0, h_s_cla12_pg_logic10_xor0);
  xor_gate xor_gate_h_s_cla12_xor10(h_s_cla12_pg_logic10_xor0[0], h_s_cla12_or18[0], h_s_cla12_xor10);
  and_gate and_gate_h_s_cla12_and36(h_s_cla12_or15[0], h_s_cla12_pg_logic9_or0[0], h_s_cla12_and36);
  and_gate and_gate_h_s_cla12_and37(h_s_cla12_pg_logic10_or0[0], h_s_cla12_pg_logic8_or0[0], h_s_cla12_and37);
  and_gate and_gate_h_s_cla12_and38(h_s_cla12_and36[0], h_s_cla12_and37[0], h_s_cla12_and38);
  and_gate and_gate_h_s_cla12_and39(h_s_cla12_pg_logic8_and0[0], h_s_cla12_pg_logic10_or0[0], h_s_cla12_and39);
  and_gate and_gate_h_s_cla12_and40(h_s_cla12_and39[0], h_s_cla12_pg_logic9_or0[0], h_s_cla12_and40);
  and_gate and_gate_h_s_cla12_and41(h_s_cla12_pg_logic9_and0[0], h_s_cla12_pg_logic10_or0[0], h_s_cla12_and41);
  or_gate or_gate_h_s_cla12_or19(h_s_cla12_and38[0], h_s_cla12_and40[0], h_s_cla12_or19);
  or_gate or_gate_h_s_cla12_or20(h_s_cla12_or19[0], h_s_cla12_and41[0], h_s_cla12_or20);
  or_gate or_gate_h_s_cla12_or21(h_s_cla12_pg_logic10_and0[0], h_s_cla12_or20[0], h_s_cla12_or21);
  pg_logic pg_logic_h_s_cla12_pg_logic11_out(a[11], b[11], h_s_cla12_pg_logic11_or0, h_s_cla12_pg_logic11_and0, h_s_cla12_pg_logic11_xor0);
  xor_gate xor_gate_h_s_cla12_xor11(h_s_cla12_pg_logic11_xor0[0], h_s_cla12_or21[0], h_s_cla12_xor11);
  and_gate and_gate_h_s_cla12_and42(h_s_cla12_or15[0], h_s_cla12_pg_logic10_or0[0], h_s_cla12_and42);
  and_gate and_gate_h_s_cla12_and43(h_s_cla12_pg_logic11_or0[0], h_s_cla12_pg_logic9_or0[0], h_s_cla12_and43);
  and_gate and_gate_h_s_cla12_and44(h_s_cla12_and42[0], h_s_cla12_and43[0], h_s_cla12_and44);
  and_gate and_gate_h_s_cla12_and45(h_s_cla12_and44[0], h_s_cla12_pg_logic8_or0[0], h_s_cla12_and45);
  and_gate and_gate_h_s_cla12_and46(h_s_cla12_pg_logic8_and0[0], h_s_cla12_pg_logic10_or0[0], h_s_cla12_and46);
  and_gate and_gate_h_s_cla12_and47(h_s_cla12_pg_logic11_or0[0], h_s_cla12_pg_logic9_or0[0], h_s_cla12_and47);
  and_gate and_gate_h_s_cla12_and48(h_s_cla12_and46[0], h_s_cla12_and47[0], h_s_cla12_and48);
  and_gate and_gate_h_s_cla12_and49(h_s_cla12_pg_logic9_and0[0], h_s_cla12_pg_logic11_or0[0], h_s_cla12_and49);
  and_gate and_gate_h_s_cla12_and50(h_s_cla12_and49[0], h_s_cla12_pg_logic10_or0[0], h_s_cla12_and50);
  and_gate and_gate_h_s_cla12_and51(h_s_cla12_pg_logic10_and0[0], h_s_cla12_pg_logic11_or0[0], h_s_cla12_and51);
  or_gate or_gate_h_s_cla12_or22(h_s_cla12_and45[0], h_s_cla12_and50[0], h_s_cla12_or22);
  or_gate or_gate_h_s_cla12_or23(h_s_cla12_and48[0], h_s_cla12_and51[0], h_s_cla12_or23);
  or_gate or_gate_h_s_cla12_or24(h_s_cla12_or22[0], h_s_cla12_or23[0], h_s_cla12_or24);
  or_gate or_gate_h_s_cla12_or25(h_s_cla12_pg_logic11_and0[0], h_s_cla12_or24[0], h_s_cla12_or25);
  xor_gate xor_gate_h_s_cla12_xor12(a[11], b[11], h_s_cla12_xor12);
  xor_gate xor_gate_h_s_cla12_xor13(h_s_cla12_xor12[0], h_s_cla12_or25[0], h_s_cla12_xor13);

  assign h_s_cla12_out[0] = h_s_cla12_pg_logic0_xor0[0];
  assign h_s_cla12_out[1] = h_s_cla12_xor1[0];
  assign h_s_cla12_out[2] = h_s_cla12_xor2[0];
  assign h_s_cla12_out[3] = h_s_cla12_xor3[0];
  assign h_s_cla12_out[4] = h_s_cla12_xor4[0];
  assign h_s_cla12_out[5] = h_s_cla12_xor5[0];
  assign h_s_cla12_out[6] = h_s_cla12_xor6[0];
  assign h_s_cla12_out[7] = h_s_cla12_xor7[0];
  assign h_s_cla12_out[8] = h_s_cla12_xor8[0];
  assign h_s_cla12_out[9] = h_s_cla12_xor9[0];
  assign h_s_cla12_out[10] = h_s_cla12_xor10[0];
  assign h_s_cla12_out[11] = h_s_cla12_xor11[0];
  assign h_s_cla12_out[12] = h_s_cla12_xor13[0];
endmodule