module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module csa_component10(input [9:0] a, input [9:0] b, input [9:0] c, output [21:0] csa_component10_out);
  wire [0:0] csa_component10_fa0_xor1;
  wire [0:0] csa_component10_fa0_or0;
  wire [0:0] csa_component10_fa1_xor1;
  wire [0:0] csa_component10_fa1_or0;
  wire [0:0] csa_component10_fa2_xor1;
  wire [0:0] csa_component10_fa2_or0;
  wire [0:0] csa_component10_fa3_xor1;
  wire [0:0] csa_component10_fa3_or0;
  wire [0:0] csa_component10_fa4_xor1;
  wire [0:0] csa_component10_fa4_or0;
  wire [0:0] csa_component10_fa5_xor1;
  wire [0:0] csa_component10_fa5_or0;
  wire [0:0] csa_component10_fa6_xor1;
  wire [0:0] csa_component10_fa6_or0;
  wire [0:0] csa_component10_fa7_xor1;
  wire [0:0] csa_component10_fa7_or0;
  wire [0:0] csa_component10_fa8_xor1;
  wire [0:0] csa_component10_fa8_or0;
  wire [0:0] csa_component10_fa9_xor1;
  wire [0:0] csa_component10_fa9_or0;

  fa fa_csa_component10_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component10_fa0_xor1), .fa_or0(csa_component10_fa0_or0));
  fa fa_csa_component10_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component10_fa1_xor1), .fa_or0(csa_component10_fa1_or0));
  fa fa_csa_component10_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component10_fa2_xor1), .fa_or0(csa_component10_fa2_or0));
  fa fa_csa_component10_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component10_fa3_xor1), .fa_or0(csa_component10_fa3_or0));
  fa fa_csa_component10_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component10_fa4_xor1), .fa_or0(csa_component10_fa4_or0));
  fa fa_csa_component10_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component10_fa5_xor1), .fa_or0(csa_component10_fa5_or0));
  fa fa_csa_component10_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component10_fa6_xor1), .fa_or0(csa_component10_fa6_or0));
  fa fa_csa_component10_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component10_fa7_xor1), .fa_or0(csa_component10_fa7_or0));
  fa fa_csa_component10_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component10_fa8_xor1), .fa_or0(csa_component10_fa8_or0));
  fa fa_csa_component10_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component10_fa9_xor1), .fa_or0(csa_component10_fa9_or0));

  assign csa_component10_out[0] = csa_component10_fa0_xor1[0];
  assign csa_component10_out[1] = csa_component10_fa1_xor1[0];
  assign csa_component10_out[2] = csa_component10_fa2_xor1[0];
  assign csa_component10_out[3] = csa_component10_fa3_xor1[0];
  assign csa_component10_out[4] = csa_component10_fa4_xor1[0];
  assign csa_component10_out[5] = csa_component10_fa5_xor1[0];
  assign csa_component10_out[6] = csa_component10_fa6_xor1[0];
  assign csa_component10_out[7] = csa_component10_fa7_xor1[0];
  assign csa_component10_out[8] = csa_component10_fa8_xor1[0];
  assign csa_component10_out[9] = csa_component10_fa9_xor1[0];
  assign csa_component10_out[10] = 1'b0;
  assign csa_component10_out[11] = 1'b0;
  assign csa_component10_out[12] = csa_component10_fa0_or0[0];
  assign csa_component10_out[13] = csa_component10_fa1_or0[0];
  assign csa_component10_out[14] = csa_component10_fa2_or0[0];
  assign csa_component10_out[15] = csa_component10_fa3_or0[0];
  assign csa_component10_out[16] = csa_component10_fa4_or0[0];
  assign csa_component10_out[17] = csa_component10_fa5_or0[0];
  assign csa_component10_out[18] = csa_component10_fa6_or0[0];
  assign csa_component10_out[19] = csa_component10_fa7_or0[0];
  assign csa_component10_out[20] = csa_component10_fa8_or0[0];
  assign csa_component10_out[21] = csa_component10_fa9_or0[0];
endmodule

module csa_component13(input [12:0] a, input [12:0] b, input [12:0] c, output [27:0] csa_component13_out);
  wire [0:0] csa_component13_fa0_xor1;
  wire [0:0] csa_component13_fa0_or0;
  wire [0:0] csa_component13_fa1_xor1;
  wire [0:0] csa_component13_fa1_or0;
  wire [0:0] csa_component13_fa2_xor1;
  wire [0:0] csa_component13_fa2_or0;
  wire [0:0] csa_component13_fa3_xor1;
  wire [0:0] csa_component13_fa3_or0;
  wire [0:0] csa_component13_fa4_xor1;
  wire [0:0] csa_component13_fa4_or0;
  wire [0:0] csa_component13_fa5_xor1;
  wire [0:0] csa_component13_fa5_or0;
  wire [0:0] csa_component13_fa6_xor1;
  wire [0:0] csa_component13_fa6_or0;
  wire [0:0] csa_component13_fa7_xor1;
  wire [0:0] csa_component13_fa7_or0;
  wire [0:0] csa_component13_fa8_xor1;
  wire [0:0] csa_component13_fa8_or0;
  wire [0:0] csa_component13_fa9_xor1;
  wire [0:0] csa_component13_fa9_or0;
  wire [0:0] csa_component13_fa10_xor1;
  wire [0:0] csa_component13_fa10_or0;
  wire [0:0] csa_component13_fa11_xor1;
  wire [0:0] csa_component13_fa11_or0;
  wire [0:0] csa_component13_fa12_xor1;
  wire [0:0] csa_component13_fa12_or0;

  fa fa_csa_component13_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component13_fa0_xor1), .fa_or0(csa_component13_fa0_or0));
  fa fa_csa_component13_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component13_fa1_xor1), .fa_or0(csa_component13_fa1_or0));
  fa fa_csa_component13_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component13_fa2_xor1), .fa_or0(csa_component13_fa2_or0));
  fa fa_csa_component13_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component13_fa3_xor1), .fa_or0(csa_component13_fa3_or0));
  fa fa_csa_component13_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component13_fa4_xor1), .fa_or0(csa_component13_fa4_or0));
  fa fa_csa_component13_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component13_fa5_xor1), .fa_or0(csa_component13_fa5_or0));
  fa fa_csa_component13_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component13_fa6_xor1), .fa_or0(csa_component13_fa6_or0));
  fa fa_csa_component13_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component13_fa7_xor1), .fa_or0(csa_component13_fa7_or0));
  fa fa_csa_component13_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component13_fa8_xor1), .fa_or0(csa_component13_fa8_or0));
  fa fa_csa_component13_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component13_fa9_xor1), .fa_or0(csa_component13_fa9_or0));
  fa fa_csa_component13_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component13_fa10_xor1), .fa_or0(csa_component13_fa10_or0));
  fa fa_csa_component13_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component13_fa11_xor1), .fa_or0(csa_component13_fa11_or0));
  fa fa_csa_component13_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component13_fa12_xor1), .fa_or0(csa_component13_fa12_or0));

  assign csa_component13_out[0] = csa_component13_fa0_xor1[0];
  assign csa_component13_out[1] = csa_component13_fa1_xor1[0];
  assign csa_component13_out[2] = csa_component13_fa2_xor1[0];
  assign csa_component13_out[3] = csa_component13_fa3_xor1[0];
  assign csa_component13_out[4] = csa_component13_fa4_xor1[0];
  assign csa_component13_out[5] = csa_component13_fa5_xor1[0];
  assign csa_component13_out[6] = csa_component13_fa6_xor1[0];
  assign csa_component13_out[7] = csa_component13_fa7_xor1[0];
  assign csa_component13_out[8] = csa_component13_fa8_xor1[0];
  assign csa_component13_out[9] = csa_component13_fa9_xor1[0];
  assign csa_component13_out[10] = csa_component13_fa10_xor1[0];
  assign csa_component13_out[11] = csa_component13_fa11_xor1[0];
  assign csa_component13_out[12] = csa_component13_fa12_xor1[0];
  assign csa_component13_out[13] = 1'b0;
  assign csa_component13_out[14] = 1'b0;
  assign csa_component13_out[15] = csa_component13_fa0_or0[0];
  assign csa_component13_out[16] = csa_component13_fa1_or0[0];
  assign csa_component13_out[17] = csa_component13_fa2_or0[0];
  assign csa_component13_out[18] = csa_component13_fa3_or0[0];
  assign csa_component13_out[19] = csa_component13_fa4_or0[0];
  assign csa_component13_out[20] = csa_component13_fa5_or0[0];
  assign csa_component13_out[21] = csa_component13_fa6_or0[0];
  assign csa_component13_out[22] = csa_component13_fa7_or0[0];
  assign csa_component13_out[23] = csa_component13_fa8_or0[0];
  assign csa_component13_out[24] = csa_component13_fa9_or0[0];
  assign csa_component13_out[25] = csa_component13_fa10_or0[0];
  assign csa_component13_out[26] = csa_component13_fa11_or0[0];
  assign csa_component13_out[27] = csa_component13_fa12_or0[0];
endmodule

module csa_component14(input [13:0] a, input [13:0] b, input [13:0] c, output [29:0] csa_component14_out);
  wire [0:0] csa_component14_fa0_xor1;
  wire [0:0] csa_component14_fa0_or0;
  wire [0:0] csa_component14_fa1_xor1;
  wire [0:0] csa_component14_fa1_or0;
  wire [0:0] csa_component14_fa2_xor1;
  wire [0:0] csa_component14_fa2_or0;
  wire [0:0] csa_component14_fa3_xor1;
  wire [0:0] csa_component14_fa3_or0;
  wire [0:0] csa_component14_fa4_xor1;
  wire [0:0] csa_component14_fa4_or0;
  wire [0:0] csa_component14_fa5_xor1;
  wire [0:0] csa_component14_fa5_or0;
  wire [0:0] csa_component14_fa6_xor1;
  wire [0:0] csa_component14_fa6_or0;
  wire [0:0] csa_component14_fa7_xor1;
  wire [0:0] csa_component14_fa7_or0;
  wire [0:0] csa_component14_fa8_xor1;
  wire [0:0] csa_component14_fa8_or0;
  wire [0:0] csa_component14_fa9_xor1;
  wire [0:0] csa_component14_fa9_or0;
  wire [0:0] csa_component14_fa10_xor1;
  wire [0:0] csa_component14_fa10_or0;
  wire [0:0] csa_component14_fa11_xor1;
  wire [0:0] csa_component14_fa11_or0;
  wire [0:0] csa_component14_fa12_xor1;
  wire [0:0] csa_component14_fa12_or0;
  wire [0:0] csa_component14_fa13_xor1;
  wire [0:0] csa_component14_fa13_or0;

  fa fa_csa_component14_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component14_fa0_xor1), .fa_or0(csa_component14_fa0_or0));
  fa fa_csa_component14_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component14_fa1_xor1), .fa_or0(csa_component14_fa1_or0));
  fa fa_csa_component14_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component14_fa2_xor1), .fa_or0(csa_component14_fa2_or0));
  fa fa_csa_component14_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component14_fa3_xor1), .fa_or0(csa_component14_fa3_or0));
  fa fa_csa_component14_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component14_fa4_xor1), .fa_or0(csa_component14_fa4_or0));
  fa fa_csa_component14_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component14_fa5_xor1), .fa_or0(csa_component14_fa5_or0));
  fa fa_csa_component14_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component14_fa6_xor1), .fa_or0(csa_component14_fa6_or0));
  fa fa_csa_component14_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component14_fa7_xor1), .fa_or0(csa_component14_fa7_or0));
  fa fa_csa_component14_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component14_fa8_xor1), .fa_or0(csa_component14_fa8_or0));
  fa fa_csa_component14_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component14_fa9_xor1), .fa_or0(csa_component14_fa9_or0));
  fa fa_csa_component14_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component14_fa10_xor1), .fa_or0(csa_component14_fa10_or0));
  fa fa_csa_component14_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component14_fa11_xor1), .fa_or0(csa_component14_fa11_or0));
  fa fa_csa_component14_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component14_fa12_xor1), .fa_or0(csa_component14_fa12_or0));
  fa fa_csa_component14_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component14_fa13_xor1), .fa_or0(csa_component14_fa13_or0));

  assign csa_component14_out[0] = csa_component14_fa0_xor1[0];
  assign csa_component14_out[1] = csa_component14_fa1_xor1[0];
  assign csa_component14_out[2] = csa_component14_fa2_xor1[0];
  assign csa_component14_out[3] = csa_component14_fa3_xor1[0];
  assign csa_component14_out[4] = csa_component14_fa4_xor1[0];
  assign csa_component14_out[5] = csa_component14_fa5_xor1[0];
  assign csa_component14_out[6] = csa_component14_fa6_xor1[0];
  assign csa_component14_out[7] = csa_component14_fa7_xor1[0];
  assign csa_component14_out[8] = csa_component14_fa8_xor1[0];
  assign csa_component14_out[9] = csa_component14_fa9_xor1[0];
  assign csa_component14_out[10] = csa_component14_fa10_xor1[0];
  assign csa_component14_out[11] = csa_component14_fa11_xor1[0];
  assign csa_component14_out[12] = csa_component14_fa12_xor1[0];
  assign csa_component14_out[13] = csa_component14_fa13_xor1[0];
  assign csa_component14_out[14] = 1'b0;
  assign csa_component14_out[15] = 1'b0;
  assign csa_component14_out[16] = csa_component14_fa0_or0[0];
  assign csa_component14_out[17] = csa_component14_fa1_or0[0];
  assign csa_component14_out[18] = csa_component14_fa2_or0[0];
  assign csa_component14_out[19] = csa_component14_fa3_or0[0];
  assign csa_component14_out[20] = csa_component14_fa4_or0[0];
  assign csa_component14_out[21] = csa_component14_fa5_or0[0];
  assign csa_component14_out[22] = csa_component14_fa6_or0[0];
  assign csa_component14_out[23] = csa_component14_fa7_or0[0];
  assign csa_component14_out[24] = csa_component14_fa8_or0[0];
  assign csa_component14_out[25] = csa_component14_fa9_or0[0];
  assign csa_component14_out[26] = csa_component14_fa10_or0[0];
  assign csa_component14_out[27] = csa_component14_fa11_or0[0];
  assign csa_component14_out[28] = csa_component14_fa12_or0[0];
  assign csa_component14_out[29] = csa_component14_fa13_or0[0];
endmodule

module csa_component15(input [14:0] a, input [14:0] b, input [14:0] c, output [31:0] csa_component15_out);
  wire [0:0] csa_component15_fa0_xor1;
  wire [0:0] csa_component15_fa0_or0;
  wire [0:0] csa_component15_fa1_xor1;
  wire [0:0] csa_component15_fa1_or0;
  wire [0:0] csa_component15_fa2_xor1;
  wire [0:0] csa_component15_fa2_or0;
  wire [0:0] csa_component15_fa3_xor1;
  wire [0:0] csa_component15_fa3_or0;
  wire [0:0] csa_component15_fa4_xor1;
  wire [0:0] csa_component15_fa4_or0;
  wire [0:0] csa_component15_fa5_xor1;
  wire [0:0] csa_component15_fa5_or0;
  wire [0:0] csa_component15_fa6_xor1;
  wire [0:0] csa_component15_fa6_or0;
  wire [0:0] csa_component15_fa7_xor1;
  wire [0:0] csa_component15_fa7_or0;
  wire [0:0] csa_component15_fa8_xor1;
  wire [0:0] csa_component15_fa8_or0;
  wire [0:0] csa_component15_fa9_xor1;
  wire [0:0] csa_component15_fa9_or0;
  wire [0:0] csa_component15_fa10_xor1;
  wire [0:0] csa_component15_fa10_or0;
  wire [0:0] csa_component15_fa11_xor1;
  wire [0:0] csa_component15_fa11_or0;
  wire [0:0] csa_component15_fa12_xor1;
  wire [0:0] csa_component15_fa12_or0;
  wire [0:0] csa_component15_fa13_xor1;
  wire [0:0] csa_component15_fa13_or0;
  wire [0:0] csa_component15_fa14_xor1;
  wire [0:0] csa_component15_fa14_or0;

  fa fa_csa_component15_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component15_fa0_xor1), .fa_or0(csa_component15_fa0_or0));
  fa fa_csa_component15_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component15_fa1_xor1), .fa_or0(csa_component15_fa1_or0));
  fa fa_csa_component15_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component15_fa2_xor1), .fa_or0(csa_component15_fa2_or0));
  fa fa_csa_component15_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component15_fa3_xor1), .fa_or0(csa_component15_fa3_or0));
  fa fa_csa_component15_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component15_fa4_xor1), .fa_or0(csa_component15_fa4_or0));
  fa fa_csa_component15_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component15_fa5_xor1), .fa_or0(csa_component15_fa5_or0));
  fa fa_csa_component15_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component15_fa6_xor1), .fa_or0(csa_component15_fa6_or0));
  fa fa_csa_component15_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component15_fa7_xor1), .fa_or0(csa_component15_fa7_or0));
  fa fa_csa_component15_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component15_fa8_xor1), .fa_or0(csa_component15_fa8_or0));
  fa fa_csa_component15_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component15_fa9_xor1), .fa_or0(csa_component15_fa9_or0));
  fa fa_csa_component15_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component15_fa10_xor1), .fa_or0(csa_component15_fa10_or0));
  fa fa_csa_component15_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component15_fa11_xor1), .fa_or0(csa_component15_fa11_or0));
  fa fa_csa_component15_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component15_fa12_xor1), .fa_or0(csa_component15_fa12_or0));
  fa fa_csa_component15_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component15_fa13_xor1), .fa_or0(csa_component15_fa13_or0));
  fa fa_csa_component15_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component15_fa14_xor1), .fa_or0(csa_component15_fa14_or0));

  assign csa_component15_out[0] = csa_component15_fa0_xor1[0];
  assign csa_component15_out[1] = csa_component15_fa1_xor1[0];
  assign csa_component15_out[2] = csa_component15_fa2_xor1[0];
  assign csa_component15_out[3] = csa_component15_fa3_xor1[0];
  assign csa_component15_out[4] = csa_component15_fa4_xor1[0];
  assign csa_component15_out[5] = csa_component15_fa5_xor1[0];
  assign csa_component15_out[6] = csa_component15_fa6_xor1[0];
  assign csa_component15_out[7] = csa_component15_fa7_xor1[0];
  assign csa_component15_out[8] = csa_component15_fa8_xor1[0];
  assign csa_component15_out[9] = csa_component15_fa9_xor1[0];
  assign csa_component15_out[10] = csa_component15_fa10_xor1[0];
  assign csa_component15_out[11] = csa_component15_fa11_xor1[0];
  assign csa_component15_out[12] = csa_component15_fa12_xor1[0];
  assign csa_component15_out[13] = csa_component15_fa13_xor1[0];
  assign csa_component15_out[14] = csa_component15_fa14_xor1[0];
  assign csa_component15_out[15] = 1'b0;
  assign csa_component15_out[16] = 1'b0;
  assign csa_component15_out[17] = csa_component15_fa0_or0[0];
  assign csa_component15_out[18] = csa_component15_fa1_or0[0];
  assign csa_component15_out[19] = csa_component15_fa2_or0[0];
  assign csa_component15_out[20] = csa_component15_fa3_or0[0];
  assign csa_component15_out[21] = csa_component15_fa4_or0[0];
  assign csa_component15_out[22] = csa_component15_fa5_or0[0];
  assign csa_component15_out[23] = csa_component15_fa6_or0[0];
  assign csa_component15_out[24] = csa_component15_fa7_or0[0];
  assign csa_component15_out[25] = csa_component15_fa8_or0[0];
  assign csa_component15_out[26] = csa_component15_fa9_or0[0];
  assign csa_component15_out[27] = csa_component15_fa10_or0[0];
  assign csa_component15_out[28] = csa_component15_fa11_or0[0];
  assign csa_component15_out[29] = csa_component15_fa12_or0[0];
  assign csa_component15_out[30] = csa_component15_fa13_or0[0];
  assign csa_component15_out[31] = csa_component15_fa14_or0[0];
endmodule

module csa_component16(input [15:0] a, input [15:0] b, input [15:0] c, output [33:0] csa_component16_out);
  wire [0:0] csa_component16_fa0_xor1;
  wire [0:0] csa_component16_fa0_or0;
  wire [0:0] csa_component16_fa1_xor1;
  wire [0:0] csa_component16_fa1_or0;
  wire [0:0] csa_component16_fa2_xor1;
  wire [0:0] csa_component16_fa2_or0;
  wire [0:0] csa_component16_fa3_xor1;
  wire [0:0] csa_component16_fa3_or0;
  wire [0:0] csa_component16_fa4_xor1;
  wire [0:0] csa_component16_fa4_or0;
  wire [0:0] csa_component16_fa5_xor1;
  wire [0:0] csa_component16_fa5_or0;
  wire [0:0] csa_component16_fa6_xor1;
  wire [0:0] csa_component16_fa6_or0;
  wire [0:0] csa_component16_fa7_xor1;
  wire [0:0] csa_component16_fa7_or0;
  wire [0:0] csa_component16_fa8_xor1;
  wire [0:0] csa_component16_fa8_or0;
  wire [0:0] csa_component16_fa9_xor1;
  wire [0:0] csa_component16_fa9_or0;
  wire [0:0] csa_component16_fa10_xor1;
  wire [0:0] csa_component16_fa10_or0;
  wire [0:0] csa_component16_fa11_xor1;
  wire [0:0] csa_component16_fa11_or0;
  wire [0:0] csa_component16_fa12_xor1;
  wire [0:0] csa_component16_fa12_or0;
  wire [0:0] csa_component16_fa13_xor1;
  wire [0:0] csa_component16_fa13_or0;
  wire [0:0] csa_component16_fa14_xor1;
  wire [0:0] csa_component16_fa14_or0;
  wire [0:0] csa_component16_fa15_xor1;
  wire [0:0] csa_component16_fa15_or0;

  fa fa_csa_component16_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component16_fa0_xor1), .fa_or0(csa_component16_fa0_or0));
  fa fa_csa_component16_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component16_fa1_xor1), .fa_or0(csa_component16_fa1_or0));
  fa fa_csa_component16_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component16_fa2_xor1), .fa_or0(csa_component16_fa2_or0));
  fa fa_csa_component16_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component16_fa3_xor1), .fa_or0(csa_component16_fa3_or0));
  fa fa_csa_component16_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component16_fa4_xor1), .fa_or0(csa_component16_fa4_or0));
  fa fa_csa_component16_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component16_fa5_xor1), .fa_or0(csa_component16_fa5_or0));
  fa fa_csa_component16_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component16_fa6_xor1), .fa_or0(csa_component16_fa6_or0));
  fa fa_csa_component16_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component16_fa7_xor1), .fa_or0(csa_component16_fa7_or0));
  fa fa_csa_component16_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component16_fa8_xor1), .fa_or0(csa_component16_fa8_or0));
  fa fa_csa_component16_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component16_fa9_xor1), .fa_or0(csa_component16_fa9_or0));
  fa fa_csa_component16_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component16_fa10_xor1), .fa_or0(csa_component16_fa10_or0));
  fa fa_csa_component16_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component16_fa11_xor1), .fa_or0(csa_component16_fa11_or0));
  fa fa_csa_component16_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component16_fa12_xor1), .fa_or0(csa_component16_fa12_or0));
  fa fa_csa_component16_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component16_fa13_xor1), .fa_or0(csa_component16_fa13_or0));
  fa fa_csa_component16_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component16_fa14_xor1), .fa_or0(csa_component16_fa14_or0));
  fa fa_csa_component16_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component16_fa15_xor1), .fa_or0(csa_component16_fa15_or0));

  assign csa_component16_out[0] = csa_component16_fa0_xor1[0];
  assign csa_component16_out[1] = csa_component16_fa1_xor1[0];
  assign csa_component16_out[2] = csa_component16_fa2_xor1[0];
  assign csa_component16_out[3] = csa_component16_fa3_xor1[0];
  assign csa_component16_out[4] = csa_component16_fa4_xor1[0];
  assign csa_component16_out[5] = csa_component16_fa5_xor1[0];
  assign csa_component16_out[6] = csa_component16_fa6_xor1[0];
  assign csa_component16_out[7] = csa_component16_fa7_xor1[0];
  assign csa_component16_out[8] = csa_component16_fa8_xor1[0];
  assign csa_component16_out[9] = csa_component16_fa9_xor1[0];
  assign csa_component16_out[10] = csa_component16_fa10_xor1[0];
  assign csa_component16_out[11] = csa_component16_fa11_xor1[0];
  assign csa_component16_out[12] = csa_component16_fa12_xor1[0];
  assign csa_component16_out[13] = csa_component16_fa13_xor1[0];
  assign csa_component16_out[14] = csa_component16_fa14_xor1[0];
  assign csa_component16_out[15] = csa_component16_fa15_xor1[0];
  assign csa_component16_out[16] = 1'b0;
  assign csa_component16_out[17] = 1'b0;
  assign csa_component16_out[18] = csa_component16_fa0_or0[0];
  assign csa_component16_out[19] = csa_component16_fa1_or0[0];
  assign csa_component16_out[20] = csa_component16_fa2_or0[0];
  assign csa_component16_out[21] = csa_component16_fa3_or0[0];
  assign csa_component16_out[22] = csa_component16_fa4_or0[0];
  assign csa_component16_out[23] = csa_component16_fa5_or0[0];
  assign csa_component16_out[24] = csa_component16_fa6_or0[0];
  assign csa_component16_out[25] = csa_component16_fa7_or0[0];
  assign csa_component16_out[26] = csa_component16_fa8_or0[0];
  assign csa_component16_out[27] = csa_component16_fa9_or0[0];
  assign csa_component16_out[28] = csa_component16_fa10_or0[0];
  assign csa_component16_out[29] = csa_component16_fa11_or0[0];
  assign csa_component16_out[30] = csa_component16_fa12_or0[0];
  assign csa_component16_out[31] = csa_component16_fa13_or0[0];
  assign csa_component16_out[32] = csa_component16_fa14_or0[0];
  assign csa_component16_out[33] = csa_component16_fa15_or0[0];
endmodule

module u_cska16(input [15:0] a, input [15:0] b, output [16:0] u_cska16_out);
  wire [0:0] u_cska16_xor0;
  wire [0:0] u_cska16_ha0_xor0;
  wire [0:0] u_cska16_ha0_and0;
  wire [0:0] u_cska16_xor1;
  wire [0:0] u_cska16_fa0_xor1;
  wire [0:0] u_cska16_fa0_or0;
  wire [0:0] u_cska16_xor2;
  wire [0:0] u_cska16_fa1_xor1;
  wire [0:0] u_cska16_fa1_or0;
  wire [0:0] u_cska16_xor3;
  wire [0:0] u_cska16_fa2_xor1;
  wire [0:0] u_cska16_fa2_or0;
  wire [0:0] u_cska16_and_propagate00;
  wire [0:0] u_cska16_and_propagate01;
  wire [0:0] u_cska16_and_propagate02;
  wire [0:0] u_cska16_mux2to10_and1;
  wire [0:0] u_cska16_xor4;
  wire [0:0] u_cska16_fa3_xor1;
  wire [0:0] u_cska16_fa3_or0;
  wire [0:0] u_cska16_xor5;
  wire [0:0] u_cska16_fa4_xor1;
  wire [0:0] u_cska16_fa4_or0;
  wire [0:0] u_cska16_xor6;
  wire [0:0] u_cska16_fa5_xor1;
  wire [0:0] u_cska16_fa5_or0;
  wire [0:0] u_cska16_xor7;
  wire [0:0] u_cska16_fa6_xor1;
  wire [0:0] u_cska16_fa6_or0;
  wire [0:0] u_cska16_and_propagate13;
  wire [0:0] u_cska16_and_propagate14;
  wire [0:0] u_cska16_and_propagate15;
  wire [0:0] u_cska16_mux2to11_xor0;
  wire [0:0] u_cska16_xor8;
  wire [0:0] u_cska16_fa7_xor1;
  wire [0:0] u_cska16_fa7_or0;
  wire [0:0] u_cska16_xor9;
  wire [0:0] u_cska16_fa8_xor1;
  wire [0:0] u_cska16_fa8_or0;
  wire [0:0] u_cska16_xor10;
  wire [0:0] u_cska16_fa9_xor1;
  wire [0:0] u_cska16_fa9_or0;
  wire [0:0] u_cska16_xor11;
  wire [0:0] u_cska16_fa10_xor1;
  wire [0:0] u_cska16_fa10_or0;
  wire [0:0] u_cska16_and_propagate26;
  wire [0:0] u_cska16_and_propagate27;
  wire [0:0] u_cska16_and_propagate28;
  wire [0:0] u_cska16_mux2to12_xor0;
  wire [0:0] u_cska16_xor12;
  wire [0:0] u_cska16_fa11_xor1;
  wire [0:0] u_cska16_fa11_or0;
  wire [0:0] u_cska16_xor13;
  wire [0:0] u_cska16_fa12_xor1;
  wire [0:0] u_cska16_fa12_or0;
  wire [0:0] u_cska16_xor14;
  wire [0:0] u_cska16_fa13_xor1;
  wire [0:0] u_cska16_fa13_or0;
  wire [0:0] u_cska16_xor15;
  wire [0:0] u_cska16_fa14_xor1;
  wire [0:0] u_cska16_fa14_or0;
  wire [0:0] u_cska16_and_propagate39;
  wire [0:0] u_cska16_and_propagate310;
  wire [0:0] u_cska16_and_propagate311;
  wire [0:0] u_cska16_mux2to13_xor0;

  xor_gate xor_gate_u_cska16_xor0(.a(a[0]), .b(b[0]), .out(u_cska16_xor0));
  ha ha_u_cska16_ha0_out(.a(a[0]), .b(b[0]), .ha_xor0(u_cska16_ha0_xor0), .ha_and0(u_cska16_ha0_and0));
  xor_gate xor_gate_u_cska16_xor1(.a(a[1]), .b(b[1]), .out(u_cska16_xor1));
  fa fa_u_cska16_fa0_out(.a(a[1]), .b(b[1]), .cin(u_cska16_ha0_and0[0]), .fa_xor1(u_cska16_fa0_xor1), .fa_or0(u_cska16_fa0_or0));
  xor_gate xor_gate_u_cska16_xor2(.a(a[2]), .b(b[2]), .out(u_cska16_xor2));
  fa fa_u_cska16_fa1_out(.a(a[2]), .b(b[2]), .cin(u_cska16_fa0_or0[0]), .fa_xor1(u_cska16_fa1_xor1), .fa_or0(u_cska16_fa1_or0));
  xor_gate xor_gate_u_cska16_xor3(.a(a[3]), .b(b[3]), .out(u_cska16_xor3));
  fa fa_u_cska16_fa2_out(.a(a[3]), .b(b[3]), .cin(u_cska16_fa1_or0[0]), .fa_xor1(u_cska16_fa2_xor1), .fa_or0(u_cska16_fa2_or0));
  and_gate and_gate_u_cska16_and_propagate00(.a(u_cska16_xor0[0]), .b(u_cska16_xor2[0]), .out(u_cska16_and_propagate00));
  and_gate and_gate_u_cska16_and_propagate01(.a(u_cska16_xor1[0]), .b(u_cska16_xor3[0]), .out(u_cska16_and_propagate01));
  and_gate and_gate_u_cska16_and_propagate02(.a(u_cska16_and_propagate00[0]), .b(u_cska16_and_propagate01[0]), .out(u_cska16_and_propagate02));
  mux2to1 mux2to1_u_cska16_mux2to10_out(.d0(u_cska16_fa2_or0[0]), .d1(1'b0), .sel(u_cska16_and_propagate02[0]), .mux2to1_xor0(u_cska16_mux2to10_and1));
  xor_gate xor_gate_u_cska16_xor4(.a(a[4]), .b(b[4]), .out(u_cska16_xor4));
  fa fa_u_cska16_fa3_out(.a(a[4]), .b(b[4]), .cin(u_cska16_mux2to10_and1[0]), .fa_xor1(u_cska16_fa3_xor1), .fa_or0(u_cska16_fa3_or0));
  xor_gate xor_gate_u_cska16_xor5(.a(a[5]), .b(b[5]), .out(u_cska16_xor5));
  fa fa_u_cska16_fa4_out(.a(a[5]), .b(b[5]), .cin(u_cska16_fa3_or0[0]), .fa_xor1(u_cska16_fa4_xor1), .fa_or0(u_cska16_fa4_or0));
  xor_gate xor_gate_u_cska16_xor6(.a(a[6]), .b(b[6]), .out(u_cska16_xor6));
  fa fa_u_cska16_fa5_out(.a(a[6]), .b(b[6]), .cin(u_cska16_fa4_or0[0]), .fa_xor1(u_cska16_fa5_xor1), .fa_or0(u_cska16_fa5_or0));
  xor_gate xor_gate_u_cska16_xor7(.a(a[7]), .b(b[7]), .out(u_cska16_xor7));
  fa fa_u_cska16_fa6_out(.a(a[7]), .b(b[7]), .cin(u_cska16_fa5_or0[0]), .fa_xor1(u_cska16_fa6_xor1), .fa_or0(u_cska16_fa6_or0));
  and_gate and_gate_u_cska16_and_propagate13(.a(u_cska16_xor4[0]), .b(u_cska16_xor6[0]), .out(u_cska16_and_propagate13));
  and_gate and_gate_u_cska16_and_propagate14(.a(u_cska16_xor5[0]), .b(u_cska16_xor7[0]), .out(u_cska16_and_propagate14));
  and_gate and_gate_u_cska16_and_propagate15(.a(u_cska16_and_propagate13[0]), .b(u_cska16_and_propagate14[0]), .out(u_cska16_and_propagate15));
  mux2to1 mux2to1_u_cska16_mux2to11_out(.d0(u_cska16_fa6_or0[0]), .d1(u_cska16_mux2to10_and1[0]), .sel(u_cska16_and_propagate15[0]), .mux2to1_xor0(u_cska16_mux2to11_xor0));
  xor_gate xor_gate_u_cska16_xor8(.a(a[8]), .b(b[8]), .out(u_cska16_xor8));
  fa fa_u_cska16_fa7_out(.a(a[8]), .b(b[8]), .cin(u_cska16_mux2to11_xor0[0]), .fa_xor1(u_cska16_fa7_xor1), .fa_or0(u_cska16_fa7_or0));
  xor_gate xor_gate_u_cska16_xor9(.a(a[9]), .b(b[9]), .out(u_cska16_xor9));
  fa fa_u_cska16_fa8_out(.a(a[9]), .b(b[9]), .cin(u_cska16_fa7_or0[0]), .fa_xor1(u_cska16_fa8_xor1), .fa_or0(u_cska16_fa8_or0));
  xor_gate xor_gate_u_cska16_xor10(.a(a[10]), .b(b[10]), .out(u_cska16_xor10));
  fa fa_u_cska16_fa9_out(.a(a[10]), .b(b[10]), .cin(u_cska16_fa8_or0[0]), .fa_xor1(u_cska16_fa9_xor1), .fa_or0(u_cska16_fa9_or0));
  xor_gate xor_gate_u_cska16_xor11(.a(a[11]), .b(b[11]), .out(u_cska16_xor11));
  fa fa_u_cska16_fa10_out(.a(a[11]), .b(b[11]), .cin(u_cska16_fa9_or0[0]), .fa_xor1(u_cska16_fa10_xor1), .fa_or0(u_cska16_fa10_or0));
  and_gate and_gate_u_cska16_and_propagate26(.a(u_cska16_xor8[0]), .b(u_cska16_xor10[0]), .out(u_cska16_and_propagate26));
  and_gate and_gate_u_cska16_and_propagate27(.a(u_cska16_xor9[0]), .b(u_cska16_xor11[0]), .out(u_cska16_and_propagate27));
  and_gate and_gate_u_cska16_and_propagate28(.a(u_cska16_and_propagate26[0]), .b(u_cska16_and_propagate27[0]), .out(u_cska16_and_propagate28));
  mux2to1 mux2to1_u_cska16_mux2to12_out(.d0(u_cska16_fa10_or0[0]), .d1(u_cska16_mux2to11_xor0[0]), .sel(u_cska16_and_propagate28[0]), .mux2to1_xor0(u_cska16_mux2to12_xor0));
  xor_gate xor_gate_u_cska16_xor12(.a(a[12]), .b(b[12]), .out(u_cska16_xor12));
  fa fa_u_cska16_fa11_out(.a(a[12]), .b(b[12]), .cin(u_cska16_mux2to12_xor0[0]), .fa_xor1(u_cska16_fa11_xor1), .fa_or0(u_cska16_fa11_or0));
  xor_gate xor_gate_u_cska16_xor13(.a(a[13]), .b(b[13]), .out(u_cska16_xor13));
  fa fa_u_cska16_fa12_out(.a(a[13]), .b(b[13]), .cin(u_cska16_fa11_or0[0]), .fa_xor1(u_cska16_fa12_xor1), .fa_or0(u_cska16_fa12_or0));
  xor_gate xor_gate_u_cska16_xor14(.a(a[14]), .b(b[14]), .out(u_cska16_xor14));
  fa fa_u_cska16_fa13_out(.a(a[14]), .b(b[14]), .cin(u_cska16_fa12_or0[0]), .fa_xor1(u_cska16_fa13_xor1), .fa_or0(u_cska16_fa13_or0));
  xor_gate xor_gate_u_cska16_xor15(.a(a[15]), .b(b[15]), .out(u_cska16_xor15));
  fa fa_u_cska16_fa14_out(.a(a[15]), .b(b[15]), .cin(u_cska16_fa13_or0[0]), .fa_xor1(u_cska16_fa14_xor1), .fa_or0(u_cska16_fa14_or0));
  and_gate and_gate_u_cska16_and_propagate39(.a(u_cska16_xor12[0]), .b(u_cska16_xor14[0]), .out(u_cska16_and_propagate39));
  and_gate and_gate_u_cska16_and_propagate310(.a(u_cska16_xor13[0]), .b(u_cska16_xor15[0]), .out(u_cska16_and_propagate310));
  and_gate and_gate_u_cska16_and_propagate311(.a(u_cska16_and_propagate39[0]), .b(u_cska16_and_propagate310[0]), .out(u_cska16_and_propagate311));
  mux2to1 mux2to1_u_cska16_mux2to13_out(.d0(u_cska16_fa14_or0[0]), .d1(u_cska16_mux2to12_xor0[0]), .sel(u_cska16_and_propagate311[0]), .mux2to1_xor0(u_cska16_mux2to13_xor0));

  assign u_cska16_out[0] = u_cska16_ha0_xor0[0];
  assign u_cska16_out[1] = u_cska16_fa0_xor1[0];
  assign u_cska16_out[2] = u_cska16_fa1_xor1[0];
  assign u_cska16_out[3] = u_cska16_fa2_xor1[0];
  assign u_cska16_out[4] = u_cska16_fa3_xor1[0];
  assign u_cska16_out[5] = u_cska16_fa4_xor1[0];
  assign u_cska16_out[6] = u_cska16_fa5_xor1[0];
  assign u_cska16_out[7] = u_cska16_fa6_xor1[0];
  assign u_cska16_out[8] = u_cska16_fa7_xor1[0];
  assign u_cska16_out[9] = u_cska16_fa8_xor1[0];
  assign u_cska16_out[10] = u_cska16_fa9_xor1[0];
  assign u_cska16_out[11] = u_cska16_fa10_xor1[0];
  assign u_cska16_out[12] = u_cska16_fa11_xor1[0];
  assign u_cska16_out[13] = u_cska16_fa12_xor1[0];
  assign u_cska16_out[14] = u_cska16_fa13_xor1[0];
  assign u_cska16_out[15] = u_cska16_fa14_xor1[0];
  assign u_cska16_out[16] = u_cska16_mux2to13_xor0[0];
endmodule

module u_CSAwallace_cska8(input [7:0] a, input [7:0] b, output [15:0] u_CSAwallace_cska8_out);
  wire [0:0] u_CSAwallace_cska8_and_0_0;
  wire [0:0] u_CSAwallace_cska8_and_1_0;
  wire [0:0] u_CSAwallace_cska8_and_2_0;
  wire [0:0] u_CSAwallace_cska8_and_3_0;
  wire [0:0] u_CSAwallace_cska8_and_4_0;
  wire [0:0] u_CSAwallace_cska8_and_5_0;
  wire [0:0] u_CSAwallace_cska8_and_6_0;
  wire [0:0] u_CSAwallace_cska8_and_7_0;
  wire [0:0] u_CSAwallace_cska8_and_0_1;
  wire [0:0] u_CSAwallace_cska8_and_1_1;
  wire [0:0] u_CSAwallace_cska8_and_2_1;
  wire [0:0] u_CSAwallace_cska8_and_3_1;
  wire [0:0] u_CSAwallace_cska8_and_4_1;
  wire [0:0] u_CSAwallace_cska8_and_5_1;
  wire [0:0] u_CSAwallace_cska8_and_6_1;
  wire [0:0] u_CSAwallace_cska8_and_7_1;
  wire [0:0] u_CSAwallace_cska8_and_0_2;
  wire [0:0] u_CSAwallace_cska8_and_1_2;
  wire [0:0] u_CSAwallace_cska8_and_2_2;
  wire [0:0] u_CSAwallace_cska8_and_3_2;
  wire [0:0] u_CSAwallace_cska8_and_4_2;
  wire [0:0] u_CSAwallace_cska8_and_5_2;
  wire [0:0] u_CSAwallace_cska8_and_6_2;
  wire [0:0] u_CSAwallace_cska8_and_7_2;
  wire [0:0] u_CSAwallace_cska8_and_0_3;
  wire [0:0] u_CSAwallace_cska8_and_1_3;
  wire [0:0] u_CSAwallace_cska8_and_2_3;
  wire [0:0] u_CSAwallace_cska8_and_3_3;
  wire [0:0] u_CSAwallace_cska8_and_4_3;
  wire [0:0] u_CSAwallace_cska8_and_5_3;
  wire [0:0] u_CSAwallace_cska8_and_6_3;
  wire [0:0] u_CSAwallace_cska8_and_7_3;
  wire [0:0] u_CSAwallace_cska8_and_0_4;
  wire [0:0] u_CSAwallace_cska8_and_1_4;
  wire [0:0] u_CSAwallace_cska8_and_2_4;
  wire [0:0] u_CSAwallace_cska8_and_3_4;
  wire [0:0] u_CSAwallace_cska8_and_4_4;
  wire [0:0] u_CSAwallace_cska8_and_5_4;
  wire [0:0] u_CSAwallace_cska8_and_6_4;
  wire [0:0] u_CSAwallace_cska8_and_7_4;
  wire [0:0] u_CSAwallace_cska8_and_0_5;
  wire [0:0] u_CSAwallace_cska8_and_1_5;
  wire [0:0] u_CSAwallace_cska8_and_2_5;
  wire [0:0] u_CSAwallace_cska8_and_3_5;
  wire [0:0] u_CSAwallace_cska8_and_4_5;
  wire [0:0] u_CSAwallace_cska8_and_5_5;
  wire [0:0] u_CSAwallace_cska8_and_6_5;
  wire [0:0] u_CSAwallace_cska8_and_7_5;
  wire [0:0] u_CSAwallace_cska8_and_0_6;
  wire [0:0] u_CSAwallace_cska8_and_1_6;
  wire [0:0] u_CSAwallace_cska8_and_2_6;
  wire [0:0] u_CSAwallace_cska8_and_3_6;
  wire [0:0] u_CSAwallace_cska8_and_4_6;
  wire [0:0] u_CSAwallace_cska8_and_5_6;
  wire [0:0] u_CSAwallace_cska8_and_6_6;
  wire [0:0] u_CSAwallace_cska8_and_7_6;
  wire [0:0] u_CSAwallace_cska8_and_0_7;
  wire [0:0] u_CSAwallace_cska8_and_1_7;
  wire [0:0] u_CSAwallace_cska8_and_2_7;
  wire [0:0] u_CSAwallace_cska8_and_3_7;
  wire [0:0] u_CSAwallace_cska8_and_4_7;
  wire [0:0] u_CSAwallace_cska8_and_5_7;
  wire [0:0] u_CSAwallace_cska8_and_6_7;
  wire [0:0] u_CSAwallace_cska8_and_7_7;
  wire [9:0] u_CSAwallace_cska8_csa0_csa_component_pp_row0;
  wire [9:0] u_CSAwallace_cska8_csa0_csa_component_pp_row1;
  wire [9:0] u_CSAwallace_cska8_csa0_csa_component_pp_row2;
  wire [21:0] u_CSAwallace_cska8_csa0_csa_component_out;
  wire [12:0] u_CSAwallace_cska8_csa1_csa_component_pp_row3;
  wire [12:0] u_CSAwallace_cska8_csa1_csa_component_pp_row4;
  wire [12:0] u_CSAwallace_cska8_csa1_csa_component_pp_row5;
  wire [27:0] u_CSAwallace_cska8_csa1_csa_component_out;
  wire [13:0] u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1;
  wire [13:0] u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1;
  wire [13:0] u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2;
  wire [29:0] u_CSAwallace_cska8_csa2_csa_component_out;
  wire [14:0] u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2;
  wire [14:0] u_CSAwallace_cska8_csa3_csa_component_pp_row6;
  wire [14:0] u_CSAwallace_cska8_csa3_csa_component_pp_row7;
  wire [31:0] u_CSAwallace_cska8_csa3_csa_component_out;
  wire [15:0] u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3;
  wire [15:0] u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3;
  wire [15:0] u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4;
  wire [33:0] u_CSAwallace_cska8_csa4_csa_component_out;
  wire [15:0] u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5;
  wire [15:0] u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5;
  wire [15:0] u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4;
  wire [33:0] u_CSAwallace_cska8_csa5_csa_component_out;
  wire [15:0] u_CSAwallace_cska8_u_cska16_a;
  wire [15:0] u_CSAwallace_cska8_u_cska16_b;
  wire [16:0] u_CSAwallace_cska8_u_cska16_out;

  and_gate and_gate_u_CSAwallace_cska8_and_0_0(.a(a[0]), .b(b[0]), .out(u_CSAwallace_cska8_and_0_0));
  and_gate and_gate_u_CSAwallace_cska8_and_1_0(.a(a[1]), .b(b[0]), .out(u_CSAwallace_cska8_and_1_0));
  and_gate and_gate_u_CSAwallace_cska8_and_2_0(.a(a[2]), .b(b[0]), .out(u_CSAwallace_cska8_and_2_0));
  and_gate and_gate_u_CSAwallace_cska8_and_3_0(.a(a[3]), .b(b[0]), .out(u_CSAwallace_cska8_and_3_0));
  and_gate and_gate_u_CSAwallace_cska8_and_4_0(.a(a[4]), .b(b[0]), .out(u_CSAwallace_cska8_and_4_0));
  and_gate and_gate_u_CSAwallace_cska8_and_5_0(.a(a[5]), .b(b[0]), .out(u_CSAwallace_cska8_and_5_0));
  and_gate and_gate_u_CSAwallace_cska8_and_6_0(.a(a[6]), .b(b[0]), .out(u_CSAwallace_cska8_and_6_0));
  and_gate and_gate_u_CSAwallace_cska8_and_7_0(.a(a[7]), .b(b[0]), .out(u_CSAwallace_cska8_and_7_0));
  and_gate and_gate_u_CSAwallace_cska8_and_0_1(.a(a[0]), .b(b[1]), .out(u_CSAwallace_cska8_and_0_1));
  and_gate and_gate_u_CSAwallace_cska8_and_1_1(.a(a[1]), .b(b[1]), .out(u_CSAwallace_cska8_and_1_1));
  and_gate and_gate_u_CSAwallace_cska8_and_2_1(.a(a[2]), .b(b[1]), .out(u_CSAwallace_cska8_and_2_1));
  and_gate and_gate_u_CSAwallace_cska8_and_3_1(.a(a[3]), .b(b[1]), .out(u_CSAwallace_cska8_and_3_1));
  and_gate and_gate_u_CSAwallace_cska8_and_4_1(.a(a[4]), .b(b[1]), .out(u_CSAwallace_cska8_and_4_1));
  and_gate and_gate_u_CSAwallace_cska8_and_5_1(.a(a[5]), .b(b[1]), .out(u_CSAwallace_cska8_and_5_1));
  and_gate and_gate_u_CSAwallace_cska8_and_6_1(.a(a[6]), .b(b[1]), .out(u_CSAwallace_cska8_and_6_1));
  and_gate and_gate_u_CSAwallace_cska8_and_7_1(.a(a[7]), .b(b[1]), .out(u_CSAwallace_cska8_and_7_1));
  and_gate and_gate_u_CSAwallace_cska8_and_0_2(.a(a[0]), .b(b[2]), .out(u_CSAwallace_cska8_and_0_2));
  and_gate and_gate_u_CSAwallace_cska8_and_1_2(.a(a[1]), .b(b[2]), .out(u_CSAwallace_cska8_and_1_2));
  and_gate and_gate_u_CSAwallace_cska8_and_2_2(.a(a[2]), .b(b[2]), .out(u_CSAwallace_cska8_and_2_2));
  and_gate and_gate_u_CSAwallace_cska8_and_3_2(.a(a[3]), .b(b[2]), .out(u_CSAwallace_cska8_and_3_2));
  and_gate and_gate_u_CSAwallace_cska8_and_4_2(.a(a[4]), .b(b[2]), .out(u_CSAwallace_cska8_and_4_2));
  and_gate and_gate_u_CSAwallace_cska8_and_5_2(.a(a[5]), .b(b[2]), .out(u_CSAwallace_cska8_and_5_2));
  and_gate and_gate_u_CSAwallace_cska8_and_6_2(.a(a[6]), .b(b[2]), .out(u_CSAwallace_cska8_and_6_2));
  and_gate and_gate_u_CSAwallace_cska8_and_7_2(.a(a[7]), .b(b[2]), .out(u_CSAwallace_cska8_and_7_2));
  and_gate and_gate_u_CSAwallace_cska8_and_0_3(.a(a[0]), .b(b[3]), .out(u_CSAwallace_cska8_and_0_3));
  and_gate and_gate_u_CSAwallace_cska8_and_1_3(.a(a[1]), .b(b[3]), .out(u_CSAwallace_cska8_and_1_3));
  and_gate and_gate_u_CSAwallace_cska8_and_2_3(.a(a[2]), .b(b[3]), .out(u_CSAwallace_cska8_and_2_3));
  and_gate and_gate_u_CSAwallace_cska8_and_3_3(.a(a[3]), .b(b[3]), .out(u_CSAwallace_cska8_and_3_3));
  and_gate and_gate_u_CSAwallace_cska8_and_4_3(.a(a[4]), .b(b[3]), .out(u_CSAwallace_cska8_and_4_3));
  and_gate and_gate_u_CSAwallace_cska8_and_5_3(.a(a[5]), .b(b[3]), .out(u_CSAwallace_cska8_and_5_3));
  and_gate and_gate_u_CSAwallace_cska8_and_6_3(.a(a[6]), .b(b[3]), .out(u_CSAwallace_cska8_and_6_3));
  and_gate and_gate_u_CSAwallace_cska8_and_7_3(.a(a[7]), .b(b[3]), .out(u_CSAwallace_cska8_and_7_3));
  and_gate and_gate_u_CSAwallace_cska8_and_0_4(.a(a[0]), .b(b[4]), .out(u_CSAwallace_cska8_and_0_4));
  and_gate and_gate_u_CSAwallace_cska8_and_1_4(.a(a[1]), .b(b[4]), .out(u_CSAwallace_cska8_and_1_4));
  and_gate and_gate_u_CSAwallace_cska8_and_2_4(.a(a[2]), .b(b[4]), .out(u_CSAwallace_cska8_and_2_4));
  and_gate and_gate_u_CSAwallace_cska8_and_3_4(.a(a[3]), .b(b[4]), .out(u_CSAwallace_cska8_and_3_4));
  and_gate and_gate_u_CSAwallace_cska8_and_4_4(.a(a[4]), .b(b[4]), .out(u_CSAwallace_cska8_and_4_4));
  and_gate and_gate_u_CSAwallace_cska8_and_5_4(.a(a[5]), .b(b[4]), .out(u_CSAwallace_cska8_and_5_4));
  and_gate and_gate_u_CSAwallace_cska8_and_6_4(.a(a[6]), .b(b[4]), .out(u_CSAwallace_cska8_and_6_4));
  and_gate and_gate_u_CSAwallace_cska8_and_7_4(.a(a[7]), .b(b[4]), .out(u_CSAwallace_cska8_and_7_4));
  and_gate and_gate_u_CSAwallace_cska8_and_0_5(.a(a[0]), .b(b[5]), .out(u_CSAwallace_cska8_and_0_5));
  and_gate and_gate_u_CSAwallace_cska8_and_1_5(.a(a[1]), .b(b[5]), .out(u_CSAwallace_cska8_and_1_5));
  and_gate and_gate_u_CSAwallace_cska8_and_2_5(.a(a[2]), .b(b[5]), .out(u_CSAwallace_cska8_and_2_5));
  and_gate and_gate_u_CSAwallace_cska8_and_3_5(.a(a[3]), .b(b[5]), .out(u_CSAwallace_cska8_and_3_5));
  and_gate and_gate_u_CSAwallace_cska8_and_4_5(.a(a[4]), .b(b[5]), .out(u_CSAwallace_cska8_and_4_5));
  and_gate and_gate_u_CSAwallace_cska8_and_5_5(.a(a[5]), .b(b[5]), .out(u_CSAwallace_cska8_and_5_5));
  and_gate and_gate_u_CSAwallace_cska8_and_6_5(.a(a[6]), .b(b[5]), .out(u_CSAwallace_cska8_and_6_5));
  and_gate and_gate_u_CSAwallace_cska8_and_7_5(.a(a[7]), .b(b[5]), .out(u_CSAwallace_cska8_and_7_5));
  and_gate and_gate_u_CSAwallace_cska8_and_0_6(.a(a[0]), .b(b[6]), .out(u_CSAwallace_cska8_and_0_6));
  and_gate and_gate_u_CSAwallace_cska8_and_1_6(.a(a[1]), .b(b[6]), .out(u_CSAwallace_cska8_and_1_6));
  and_gate and_gate_u_CSAwallace_cska8_and_2_6(.a(a[2]), .b(b[6]), .out(u_CSAwallace_cska8_and_2_6));
  and_gate and_gate_u_CSAwallace_cska8_and_3_6(.a(a[3]), .b(b[6]), .out(u_CSAwallace_cska8_and_3_6));
  and_gate and_gate_u_CSAwallace_cska8_and_4_6(.a(a[4]), .b(b[6]), .out(u_CSAwallace_cska8_and_4_6));
  and_gate and_gate_u_CSAwallace_cska8_and_5_6(.a(a[5]), .b(b[6]), .out(u_CSAwallace_cska8_and_5_6));
  and_gate and_gate_u_CSAwallace_cska8_and_6_6(.a(a[6]), .b(b[6]), .out(u_CSAwallace_cska8_and_6_6));
  and_gate and_gate_u_CSAwallace_cska8_and_7_6(.a(a[7]), .b(b[6]), .out(u_CSAwallace_cska8_and_7_6));
  and_gate and_gate_u_CSAwallace_cska8_and_0_7(.a(a[0]), .b(b[7]), .out(u_CSAwallace_cska8_and_0_7));
  and_gate and_gate_u_CSAwallace_cska8_and_1_7(.a(a[1]), .b(b[7]), .out(u_CSAwallace_cska8_and_1_7));
  and_gate and_gate_u_CSAwallace_cska8_and_2_7(.a(a[2]), .b(b[7]), .out(u_CSAwallace_cska8_and_2_7));
  and_gate and_gate_u_CSAwallace_cska8_and_3_7(.a(a[3]), .b(b[7]), .out(u_CSAwallace_cska8_and_3_7));
  and_gate and_gate_u_CSAwallace_cska8_and_4_7(.a(a[4]), .b(b[7]), .out(u_CSAwallace_cska8_and_4_7));
  and_gate and_gate_u_CSAwallace_cska8_and_5_7(.a(a[5]), .b(b[7]), .out(u_CSAwallace_cska8_and_5_7));
  and_gate and_gate_u_CSAwallace_cska8_and_6_7(.a(a[6]), .b(b[7]), .out(u_CSAwallace_cska8_and_6_7));
  and_gate and_gate_u_CSAwallace_cska8_and_7_7(.a(a[7]), .b(b[7]), .out(u_CSAwallace_cska8_and_7_7));
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[0] = u_CSAwallace_cska8_and_0_0[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[1] = u_CSAwallace_cska8_and_1_0[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[2] = u_CSAwallace_cska8_and_2_0[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[3] = u_CSAwallace_cska8_and_3_0[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[4] = u_CSAwallace_cska8_and_4_0[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[5] = u_CSAwallace_cska8_and_5_0[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[6] = u_CSAwallace_cska8_and_6_0[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[7] = u_CSAwallace_cska8_and_7_0[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[8] = 1'b0;
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row0[9] = 1'b0;
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[0] = 1'b0;
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[1] = u_CSAwallace_cska8_and_0_1[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[2] = u_CSAwallace_cska8_and_1_1[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[3] = u_CSAwallace_cska8_and_2_1[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[4] = u_CSAwallace_cska8_and_3_1[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[5] = u_CSAwallace_cska8_and_4_1[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[6] = u_CSAwallace_cska8_and_5_1[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[7] = u_CSAwallace_cska8_and_6_1[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[8] = u_CSAwallace_cska8_and_7_1[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row1[9] = 1'b0;
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[0] = 1'b0;
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[1] = 1'b0;
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[2] = u_CSAwallace_cska8_and_0_2[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[3] = u_CSAwallace_cska8_and_1_2[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[4] = u_CSAwallace_cska8_and_2_2[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[5] = u_CSAwallace_cska8_and_3_2[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[6] = u_CSAwallace_cska8_and_4_2[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[7] = u_CSAwallace_cska8_and_5_2[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[8] = u_CSAwallace_cska8_and_6_2[0];
  assign u_CSAwallace_cska8_csa0_csa_component_pp_row2[9] = u_CSAwallace_cska8_and_7_2[0];
  csa_component10 csa_component10_u_CSAwallace_cska8_csa0_csa_component_out(.a(u_CSAwallace_cska8_csa0_csa_component_pp_row0), .b(u_CSAwallace_cska8_csa0_csa_component_pp_row1), .c(u_CSAwallace_cska8_csa0_csa_component_pp_row2), .csa_component10_out(u_CSAwallace_cska8_csa0_csa_component_out));
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[0] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[1] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[2] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[3] = u_CSAwallace_cska8_and_0_3[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[4] = u_CSAwallace_cska8_and_1_3[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[5] = u_CSAwallace_cska8_and_2_3[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[6] = u_CSAwallace_cska8_and_3_3[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[7] = u_CSAwallace_cska8_and_4_3[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[8] = u_CSAwallace_cska8_and_5_3[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[9] = u_CSAwallace_cska8_and_6_3[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[10] = u_CSAwallace_cska8_and_7_3[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[11] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row3[12] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[0] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[1] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[2] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[3] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[4] = u_CSAwallace_cska8_and_0_4[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[5] = u_CSAwallace_cska8_and_1_4[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[6] = u_CSAwallace_cska8_and_2_4[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[7] = u_CSAwallace_cska8_and_3_4[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[8] = u_CSAwallace_cska8_and_4_4[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[9] = u_CSAwallace_cska8_and_5_4[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[10] = u_CSAwallace_cska8_and_6_4[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[11] = u_CSAwallace_cska8_and_7_4[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row4[12] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[0] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[1] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[2] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[3] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[4] = 1'b0;
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[5] = u_CSAwallace_cska8_and_0_5[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[6] = u_CSAwallace_cska8_and_1_5[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[7] = u_CSAwallace_cska8_and_2_5[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[8] = u_CSAwallace_cska8_and_3_5[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[9] = u_CSAwallace_cska8_and_4_5[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[10] = u_CSAwallace_cska8_and_5_5[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[11] = u_CSAwallace_cska8_and_6_5[0];
  assign u_CSAwallace_cska8_csa1_csa_component_pp_row5[12] = u_CSAwallace_cska8_and_7_5[0];
  csa_component13 csa_component13_u_CSAwallace_cska8_csa1_csa_component_out(.a(u_CSAwallace_cska8_csa1_csa_component_pp_row3), .b(u_CSAwallace_cska8_csa1_csa_component_pp_row4), .c(u_CSAwallace_cska8_csa1_csa_component_pp_row5), .csa_component13_out(u_CSAwallace_cska8_csa1_csa_component_out));
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[0] = u_CSAwallace_cska8_csa0_csa_component_out[0];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[1] = u_CSAwallace_cska8_csa0_csa_component_out[1];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[2] = u_CSAwallace_cska8_csa0_csa_component_out[2];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[3] = u_CSAwallace_cska8_csa0_csa_component_out[3];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[4] = u_CSAwallace_cska8_csa0_csa_component_out[4];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[5] = u_CSAwallace_cska8_csa0_csa_component_out[5];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[6] = u_CSAwallace_cska8_csa0_csa_component_out[6];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[7] = u_CSAwallace_cska8_csa0_csa_component_out[7];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[8] = u_CSAwallace_cska8_csa0_csa_component_out[8];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[9] = u_CSAwallace_cska8_csa0_csa_component_out[9];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[10] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[11] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[12] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1[13] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[0] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[1] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[2] = u_CSAwallace_cska8_csa0_csa_component_out[13];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[3] = u_CSAwallace_cska8_csa0_csa_component_out[14];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[4] = u_CSAwallace_cska8_csa0_csa_component_out[15];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[5] = u_CSAwallace_cska8_csa0_csa_component_out[16];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[6] = u_CSAwallace_cska8_csa0_csa_component_out[17];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[7] = u_CSAwallace_cska8_csa0_csa_component_out[18];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[8] = u_CSAwallace_cska8_csa0_csa_component_out[19];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[9] = u_CSAwallace_cska8_csa0_csa_component_out[20];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[10] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[11] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[12] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1[13] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[0] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[1] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[2] = 1'b0;
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[3] = u_CSAwallace_cska8_csa1_csa_component_out[3];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[4] = u_CSAwallace_cska8_csa1_csa_component_out[4];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[5] = u_CSAwallace_cska8_csa1_csa_component_out[5];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[6] = u_CSAwallace_cska8_csa1_csa_component_out[6];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[7] = u_CSAwallace_cska8_csa1_csa_component_out[7];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[8] = u_CSAwallace_cska8_csa1_csa_component_out[8];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[9] = u_CSAwallace_cska8_csa1_csa_component_out[9];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[10] = u_CSAwallace_cska8_csa1_csa_component_out[10];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[11] = u_CSAwallace_cska8_csa1_csa_component_out[11];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[12] = u_CSAwallace_cska8_csa1_csa_component_out[12];
  assign u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2[13] = 1'b0;
  csa_component14 csa_component14_u_CSAwallace_cska8_csa2_csa_component_out(.a(u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s1), .b(u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_c1), .c(u_CSAwallace_cska8_csa2_csa_component_u_CSAwallace_cska8_csa_s2), .csa_component14_out(u_CSAwallace_cska8_csa2_csa_component_out));
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[0] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[1] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[2] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[3] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[4] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[5] = u_CSAwallace_cska8_csa1_csa_component_out[19];
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[6] = u_CSAwallace_cska8_csa1_csa_component_out[20];
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[7] = u_CSAwallace_cska8_csa1_csa_component_out[21];
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[8] = u_CSAwallace_cska8_csa1_csa_component_out[22];
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[9] = u_CSAwallace_cska8_csa1_csa_component_out[23];
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[10] = u_CSAwallace_cska8_csa1_csa_component_out[24];
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[11] = u_CSAwallace_cska8_csa1_csa_component_out[25];
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[12] = u_CSAwallace_cska8_csa1_csa_component_out[26];
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[13] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2[14] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[0] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[1] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[2] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[3] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[4] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[5] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[6] = u_CSAwallace_cska8_and_0_6[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[7] = u_CSAwallace_cska8_and_1_6[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[8] = u_CSAwallace_cska8_and_2_6[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[9] = u_CSAwallace_cska8_and_3_6[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[10] = u_CSAwallace_cska8_and_4_6[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[11] = u_CSAwallace_cska8_and_5_6[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[12] = u_CSAwallace_cska8_and_6_6[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[13] = u_CSAwallace_cska8_and_7_6[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row6[14] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[0] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[1] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[2] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[3] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[4] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[5] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[6] = 1'b0;
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[7] = u_CSAwallace_cska8_and_0_7[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[8] = u_CSAwallace_cska8_and_1_7[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[9] = u_CSAwallace_cska8_and_2_7[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[10] = u_CSAwallace_cska8_and_3_7[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[11] = u_CSAwallace_cska8_and_4_7[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[12] = u_CSAwallace_cska8_and_5_7[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[13] = u_CSAwallace_cska8_and_6_7[0];
  assign u_CSAwallace_cska8_csa3_csa_component_pp_row7[14] = u_CSAwallace_cska8_and_7_7[0];
  csa_component15 csa_component15_u_CSAwallace_cska8_csa3_csa_component_out(.a(u_CSAwallace_cska8_csa3_csa_component_u_CSAwallace_cska8_csa_c2), .b(u_CSAwallace_cska8_csa3_csa_component_pp_row6), .c(u_CSAwallace_cska8_csa3_csa_component_pp_row7), .csa_component15_out(u_CSAwallace_cska8_csa3_csa_component_out));
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[0] = u_CSAwallace_cska8_csa2_csa_component_out[0];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[1] = u_CSAwallace_cska8_csa2_csa_component_out[1];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[2] = u_CSAwallace_cska8_csa2_csa_component_out[2];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[3] = u_CSAwallace_cska8_csa2_csa_component_out[3];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[4] = u_CSAwallace_cska8_csa2_csa_component_out[4];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[5] = u_CSAwallace_cska8_csa2_csa_component_out[5];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[6] = u_CSAwallace_cska8_csa2_csa_component_out[6];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[7] = u_CSAwallace_cska8_csa2_csa_component_out[7];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[8] = u_CSAwallace_cska8_csa2_csa_component_out[8];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[9] = u_CSAwallace_cska8_csa2_csa_component_out[9];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[10] = u_CSAwallace_cska8_csa2_csa_component_out[10];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[11] = u_CSAwallace_cska8_csa2_csa_component_out[11];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[12] = u_CSAwallace_cska8_csa2_csa_component_out[12];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[13] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[14] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3[15] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[0] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[1] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[2] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[3] = u_CSAwallace_cska8_csa2_csa_component_out[18];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[4] = u_CSAwallace_cska8_csa2_csa_component_out[19];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[5] = u_CSAwallace_cska8_csa2_csa_component_out[20];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[6] = u_CSAwallace_cska8_csa2_csa_component_out[21];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[7] = u_CSAwallace_cska8_csa2_csa_component_out[22];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[8] = u_CSAwallace_cska8_csa2_csa_component_out[23];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[9] = u_CSAwallace_cska8_csa2_csa_component_out[24];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[10] = u_CSAwallace_cska8_csa2_csa_component_out[25];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[11] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[12] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[13] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[14] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3[15] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[0] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[1] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[2] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[3] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[4] = 1'b0;
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[5] = u_CSAwallace_cska8_csa3_csa_component_out[5];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[6] = u_CSAwallace_cska8_csa3_csa_component_out[6];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[7] = u_CSAwallace_cska8_csa3_csa_component_out[7];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[8] = u_CSAwallace_cska8_csa3_csa_component_out[8];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[9] = u_CSAwallace_cska8_csa3_csa_component_out[9];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[10] = u_CSAwallace_cska8_csa3_csa_component_out[10];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[11] = u_CSAwallace_cska8_csa3_csa_component_out[11];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[12] = u_CSAwallace_cska8_csa3_csa_component_out[12];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[13] = u_CSAwallace_cska8_csa3_csa_component_out[13];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[14] = u_CSAwallace_cska8_csa3_csa_component_out[14];
  assign u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4[15] = 1'b0;
  csa_component16 csa_component16_u_CSAwallace_cska8_csa4_csa_component_out(.a(u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s3), .b(u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_c3), .c(u_CSAwallace_cska8_csa4_csa_component_u_CSAwallace_cska8_csa_s4), .csa_component16_out(u_CSAwallace_cska8_csa4_csa_component_out));
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[0] = u_CSAwallace_cska8_csa4_csa_component_out[0];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[1] = u_CSAwallace_cska8_csa4_csa_component_out[1];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[2] = u_CSAwallace_cska8_csa4_csa_component_out[2];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[3] = u_CSAwallace_cska8_csa4_csa_component_out[3];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[4] = u_CSAwallace_cska8_csa4_csa_component_out[4];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[5] = u_CSAwallace_cska8_csa4_csa_component_out[5];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[6] = u_CSAwallace_cska8_csa4_csa_component_out[6];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[7] = u_CSAwallace_cska8_csa4_csa_component_out[7];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[8] = u_CSAwallace_cska8_csa4_csa_component_out[8];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[9] = u_CSAwallace_cska8_csa4_csa_component_out[9];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[10] = u_CSAwallace_cska8_csa4_csa_component_out[10];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[11] = u_CSAwallace_cska8_csa4_csa_component_out[11];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[12] = u_CSAwallace_cska8_csa4_csa_component_out[12];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[13] = u_CSAwallace_cska8_csa4_csa_component_out[13];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[14] = u_CSAwallace_cska8_csa4_csa_component_out[14];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5[15] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[0] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[1] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[2] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[3] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[4] = u_CSAwallace_cska8_csa4_csa_component_out[21];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[5] = u_CSAwallace_cska8_csa4_csa_component_out[22];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[6] = u_CSAwallace_cska8_csa4_csa_component_out[23];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[7] = u_CSAwallace_cska8_csa4_csa_component_out[24];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[8] = u_CSAwallace_cska8_csa4_csa_component_out[25];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[9] = u_CSAwallace_cska8_csa4_csa_component_out[26];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[10] = u_CSAwallace_cska8_csa4_csa_component_out[27];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[11] = u_CSAwallace_cska8_csa4_csa_component_out[28];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[12] = u_CSAwallace_cska8_csa4_csa_component_out[29];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[13] = u_CSAwallace_cska8_csa4_csa_component_out[30];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[14] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5[15] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[0] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[1] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[2] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[3] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[4] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[5] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[6] = 1'b0;
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[7] = u_CSAwallace_cska8_csa3_csa_component_out[23];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[8] = u_CSAwallace_cska8_csa3_csa_component_out[24];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[9] = u_CSAwallace_cska8_csa3_csa_component_out[25];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[10] = u_CSAwallace_cska8_csa3_csa_component_out[26];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[11] = u_CSAwallace_cska8_csa3_csa_component_out[27];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[12] = u_CSAwallace_cska8_csa3_csa_component_out[28];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[13] = u_CSAwallace_cska8_csa3_csa_component_out[29];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[14] = u_CSAwallace_cska8_csa3_csa_component_out[30];
  assign u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4[15] = 1'b0;
  csa_component16 csa_component16_u_CSAwallace_cska8_csa5_csa_component_out(.a(u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_s5), .b(u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c5), .c(u_CSAwallace_cska8_csa5_csa_component_u_CSAwallace_cska8_csa_c4), .csa_component16_out(u_CSAwallace_cska8_csa5_csa_component_out));
  assign u_CSAwallace_cska8_u_cska16_a[0] = u_CSAwallace_cska8_csa5_csa_component_out[0];
  assign u_CSAwallace_cska8_u_cska16_a[1] = u_CSAwallace_cska8_csa5_csa_component_out[1];
  assign u_CSAwallace_cska8_u_cska16_a[2] = u_CSAwallace_cska8_csa5_csa_component_out[2];
  assign u_CSAwallace_cska8_u_cska16_a[3] = u_CSAwallace_cska8_csa5_csa_component_out[3];
  assign u_CSAwallace_cska8_u_cska16_a[4] = u_CSAwallace_cska8_csa5_csa_component_out[4];
  assign u_CSAwallace_cska8_u_cska16_a[5] = u_CSAwallace_cska8_csa5_csa_component_out[5];
  assign u_CSAwallace_cska8_u_cska16_a[6] = u_CSAwallace_cska8_csa5_csa_component_out[6];
  assign u_CSAwallace_cska8_u_cska16_a[7] = u_CSAwallace_cska8_csa5_csa_component_out[7];
  assign u_CSAwallace_cska8_u_cska16_a[8] = u_CSAwallace_cska8_csa5_csa_component_out[8];
  assign u_CSAwallace_cska8_u_cska16_a[9] = u_CSAwallace_cska8_csa5_csa_component_out[9];
  assign u_CSAwallace_cska8_u_cska16_a[10] = u_CSAwallace_cska8_csa5_csa_component_out[10];
  assign u_CSAwallace_cska8_u_cska16_a[11] = u_CSAwallace_cska8_csa5_csa_component_out[11];
  assign u_CSAwallace_cska8_u_cska16_a[12] = u_CSAwallace_cska8_csa5_csa_component_out[12];
  assign u_CSAwallace_cska8_u_cska16_a[13] = u_CSAwallace_cska8_csa5_csa_component_out[13];
  assign u_CSAwallace_cska8_u_cska16_a[14] = u_CSAwallace_cska8_csa5_csa_component_out[14];
  assign u_CSAwallace_cska8_u_cska16_a[15] = 1'b0;
  assign u_CSAwallace_cska8_u_cska16_b[0] = 1'b0;
  assign u_CSAwallace_cska8_u_cska16_b[1] = 1'b0;
  assign u_CSAwallace_cska8_u_cska16_b[2] = 1'b0;
  assign u_CSAwallace_cska8_u_cska16_b[3] = 1'b0;
  assign u_CSAwallace_cska8_u_cska16_b[4] = 1'b0;
  assign u_CSAwallace_cska8_u_cska16_b[5] = u_CSAwallace_cska8_csa5_csa_component_out[22];
  assign u_CSAwallace_cska8_u_cska16_b[6] = u_CSAwallace_cska8_csa5_csa_component_out[23];
  assign u_CSAwallace_cska8_u_cska16_b[7] = u_CSAwallace_cska8_csa5_csa_component_out[24];
  assign u_CSAwallace_cska8_u_cska16_b[8] = u_CSAwallace_cska8_csa5_csa_component_out[25];
  assign u_CSAwallace_cska8_u_cska16_b[9] = u_CSAwallace_cska8_csa5_csa_component_out[26];
  assign u_CSAwallace_cska8_u_cska16_b[10] = u_CSAwallace_cska8_csa5_csa_component_out[27];
  assign u_CSAwallace_cska8_u_cska16_b[11] = u_CSAwallace_cska8_csa5_csa_component_out[28];
  assign u_CSAwallace_cska8_u_cska16_b[12] = u_CSAwallace_cska8_csa5_csa_component_out[29];
  assign u_CSAwallace_cska8_u_cska16_b[13] = u_CSAwallace_cska8_csa5_csa_component_out[30];
  assign u_CSAwallace_cska8_u_cska16_b[14] = u_CSAwallace_cska8_csa5_csa_component_out[31];
  assign u_CSAwallace_cska8_u_cska16_b[15] = u_CSAwallace_cska8_csa5_csa_component_out[32];
  u_cska16 u_cska16_u_CSAwallace_cska8_u_cska16_out(.a(u_CSAwallace_cska8_u_cska16_a), .b(u_CSAwallace_cska8_u_cska16_b), .u_cska16_out(u_CSAwallace_cska8_u_cska16_out));

  assign u_CSAwallace_cska8_out[0] = u_CSAwallace_cska8_u_cska16_out[0];
  assign u_CSAwallace_cska8_out[1] = u_CSAwallace_cska8_u_cska16_out[1];
  assign u_CSAwallace_cska8_out[2] = u_CSAwallace_cska8_u_cska16_out[2];
  assign u_CSAwallace_cska8_out[3] = u_CSAwallace_cska8_u_cska16_out[3];
  assign u_CSAwallace_cska8_out[4] = u_CSAwallace_cska8_u_cska16_out[4];
  assign u_CSAwallace_cska8_out[5] = u_CSAwallace_cska8_u_cska16_out[5];
  assign u_CSAwallace_cska8_out[6] = u_CSAwallace_cska8_u_cska16_out[6];
  assign u_CSAwallace_cska8_out[7] = u_CSAwallace_cska8_u_cska16_out[7];
  assign u_CSAwallace_cska8_out[8] = u_CSAwallace_cska8_u_cska16_out[8];
  assign u_CSAwallace_cska8_out[9] = u_CSAwallace_cska8_u_cska16_out[9];
  assign u_CSAwallace_cska8_out[10] = u_CSAwallace_cska8_u_cska16_out[10];
  assign u_CSAwallace_cska8_out[11] = u_CSAwallace_cska8_u_cska16_out[11];
  assign u_CSAwallace_cska8_out[12] = u_CSAwallace_cska8_u_cska16_out[12];
  assign u_CSAwallace_cska8_out[13] = u_CSAwallace_cska8_u_cska16_out[13];
  assign u_CSAwallace_cska8_out[14] = u_CSAwallace_cska8_u_cska16_out[14];
  assign u_CSAwallace_cska8_out[15] = u_CSAwallace_cska8_u_cska16_out[15];
endmodule