module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module u_rca30(input [29:0] a, input [29:0] b, output [30:0] u_rca30_out);
  wire [0:0] u_rca30_ha_xor0;
  wire [0:0] u_rca30_ha_and0;
  wire [0:0] u_rca30_fa1_xor1;
  wire [0:0] u_rca30_fa1_or0;
  wire [0:0] u_rca30_fa2_xor1;
  wire [0:0] u_rca30_fa2_or0;
  wire [0:0] u_rca30_fa3_xor1;
  wire [0:0] u_rca30_fa3_or0;
  wire [0:0] u_rca30_fa4_xor1;
  wire [0:0] u_rca30_fa4_or0;
  wire [0:0] u_rca30_fa5_xor1;
  wire [0:0] u_rca30_fa5_or0;
  wire [0:0] u_rca30_fa6_xor1;
  wire [0:0] u_rca30_fa6_or0;
  wire [0:0] u_rca30_fa7_xor1;
  wire [0:0] u_rca30_fa7_or0;
  wire [0:0] u_rca30_fa8_xor1;
  wire [0:0] u_rca30_fa8_or0;
  wire [0:0] u_rca30_fa9_xor1;
  wire [0:0] u_rca30_fa9_or0;
  wire [0:0] u_rca30_fa10_xor1;
  wire [0:0] u_rca30_fa10_or0;
  wire [0:0] u_rca30_fa11_xor1;
  wire [0:0] u_rca30_fa11_or0;
  wire [0:0] u_rca30_fa12_xor1;
  wire [0:0] u_rca30_fa12_or0;
  wire [0:0] u_rca30_fa13_xor1;
  wire [0:0] u_rca30_fa13_or0;
  wire [0:0] u_rca30_fa14_xor1;
  wire [0:0] u_rca30_fa14_or0;
  wire [0:0] u_rca30_fa15_xor1;
  wire [0:0] u_rca30_fa15_or0;
  wire [0:0] u_rca30_fa16_xor1;
  wire [0:0] u_rca30_fa16_or0;
  wire [0:0] u_rca30_fa17_xor1;
  wire [0:0] u_rca30_fa17_or0;
  wire [0:0] u_rca30_fa18_xor1;
  wire [0:0] u_rca30_fa18_or0;
  wire [0:0] u_rca30_fa19_xor1;
  wire [0:0] u_rca30_fa19_or0;
  wire [0:0] u_rca30_fa20_xor1;
  wire [0:0] u_rca30_fa20_or0;
  wire [0:0] u_rca30_fa21_xor1;
  wire [0:0] u_rca30_fa21_or0;
  wire [0:0] u_rca30_fa22_xor1;
  wire [0:0] u_rca30_fa22_or0;
  wire [0:0] u_rca30_fa23_xor1;
  wire [0:0] u_rca30_fa23_or0;
  wire [0:0] u_rca30_fa24_xor1;
  wire [0:0] u_rca30_fa24_or0;
  wire [0:0] u_rca30_fa25_xor1;
  wire [0:0] u_rca30_fa25_or0;
  wire [0:0] u_rca30_fa26_xor1;
  wire [0:0] u_rca30_fa26_or0;
  wire [0:0] u_rca30_fa27_xor1;
  wire [0:0] u_rca30_fa27_or0;
  wire [0:0] u_rca30_fa28_xor1;
  wire [0:0] u_rca30_fa28_or0;
  wire [0:0] u_rca30_fa29_xor1;
  wire [0:0] u_rca30_fa29_or0;

  ha ha_u_rca30_ha_out(.a(a[0]), .b(b[0]), .ha_xor0(u_rca30_ha_xor0), .ha_and0(u_rca30_ha_and0));
  fa fa_u_rca30_fa1_out(.a(a[1]), .b(b[1]), .cin(u_rca30_ha_and0[0]), .fa_xor1(u_rca30_fa1_xor1), .fa_or0(u_rca30_fa1_or0));
  fa fa_u_rca30_fa2_out(.a(a[2]), .b(b[2]), .cin(u_rca30_fa1_or0[0]), .fa_xor1(u_rca30_fa2_xor1), .fa_or0(u_rca30_fa2_or0));
  fa fa_u_rca30_fa3_out(.a(a[3]), .b(b[3]), .cin(u_rca30_fa2_or0[0]), .fa_xor1(u_rca30_fa3_xor1), .fa_or0(u_rca30_fa3_or0));
  fa fa_u_rca30_fa4_out(.a(a[4]), .b(b[4]), .cin(u_rca30_fa3_or0[0]), .fa_xor1(u_rca30_fa4_xor1), .fa_or0(u_rca30_fa4_or0));
  fa fa_u_rca30_fa5_out(.a(a[5]), .b(b[5]), .cin(u_rca30_fa4_or0[0]), .fa_xor1(u_rca30_fa5_xor1), .fa_or0(u_rca30_fa5_or0));
  fa fa_u_rca30_fa6_out(.a(a[6]), .b(b[6]), .cin(u_rca30_fa5_or0[0]), .fa_xor1(u_rca30_fa6_xor1), .fa_or0(u_rca30_fa6_or0));
  fa fa_u_rca30_fa7_out(.a(a[7]), .b(b[7]), .cin(u_rca30_fa6_or0[0]), .fa_xor1(u_rca30_fa7_xor1), .fa_or0(u_rca30_fa7_or0));
  fa fa_u_rca30_fa8_out(.a(a[8]), .b(b[8]), .cin(u_rca30_fa7_or0[0]), .fa_xor1(u_rca30_fa8_xor1), .fa_or0(u_rca30_fa8_or0));
  fa fa_u_rca30_fa9_out(.a(a[9]), .b(b[9]), .cin(u_rca30_fa8_or0[0]), .fa_xor1(u_rca30_fa9_xor1), .fa_or0(u_rca30_fa9_or0));
  fa fa_u_rca30_fa10_out(.a(a[10]), .b(b[10]), .cin(u_rca30_fa9_or0[0]), .fa_xor1(u_rca30_fa10_xor1), .fa_or0(u_rca30_fa10_or0));
  fa fa_u_rca30_fa11_out(.a(a[11]), .b(b[11]), .cin(u_rca30_fa10_or0[0]), .fa_xor1(u_rca30_fa11_xor1), .fa_or0(u_rca30_fa11_or0));
  fa fa_u_rca30_fa12_out(.a(a[12]), .b(b[12]), .cin(u_rca30_fa11_or0[0]), .fa_xor1(u_rca30_fa12_xor1), .fa_or0(u_rca30_fa12_or0));
  fa fa_u_rca30_fa13_out(.a(a[13]), .b(b[13]), .cin(u_rca30_fa12_or0[0]), .fa_xor1(u_rca30_fa13_xor1), .fa_or0(u_rca30_fa13_or0));
  fa fa_u_rca30_fa14_out(.a(a[14]), .b(b[14]), .cin(u_rca30_fa13_or0[0]), .fa_xor1(u_rca30_fa14_xor1), .fa_or0(u_rca30_fa14_or0));
  fa fa_u_rca30_fa15_out(.a(a[15]), .b(b[15]), .cin(u_rca30_fa14_or0[0]), .fa_xor1(u_rca30_fa15_xor1), .fa_or0(u_rca30_fa15_or0));
  fa fa_u_rca30_fa16_out(.a(a[16]), .b(b[16]), .cin(u_rca30_fa15_or0[0]), .fa_xor1(u_rca30_fa16_xor1), .fa_or0(u_rca30_fa16_or0));
  fa fa_u_rca30_fa17_out(.a(a[17]), .b(b[17]), .cin(u_rca30_fa16_or0[0]), .fa_xor1(u_rca30_fa17_xor1), .fa_or0(u_rca30_fa17_or0));
  fa fa_u_rca30_fa18_out(.a(a[18]), .b(b[18]), .cin(u_rca30_fa17_or0[0]), .fa_xor1(u_rca30_fa18_xor1), .fa_or0(u_rca30_fa18_or0));
  fa fa_u_rca30_fa19_out(.a(a[19]), .b(b[19]), .cin(u_rca30_fa18_or0[0]), .fa_xor1(u_rca30_fa19_xor1), .fa_or0(u_rca30_fa19_or0));
  fa fa_u_rca30_fa20_out(.a(a[20]), .b(b[20]), .cin(u_rca30_fa19_or0[0]), .fa_xor1(u_rca30_fa20_xor1), .fa_or0(u_rca30_fa20_or0));
  fa fa_u_rca30_fa21_out(.a(a[21]), .b(b[21]), .cin(u_rca30_fa20_or0[0]), .fa_xor1(u_rca30_fa21_xor1), .fa_or0(u_rca30_fa21_or0));
  fa fa_u_rca30_fa22_out(.a(a[22]), .b(b[22]), .cin(u_rca30_fa21_or0[0]), .fa_xor1(u_rca30_fa22_xor1), .fa_or0(u_rca30_fa22_or0));
  fa fa_u_rca30_fa23_out(.a(a[23]), .b(b[23]), .cin(u_rca30_fa22_or0[0]), .fa_xor1(u_rca30_fa23_xor1), .fa_or0(u_rca30_fa23_or0));
  fa fa_u_rca30_fa24_out(.a(a[24]), .b(b[24]), .cin(u_rca30_fa23_or0[0]), .fa_xor1(u_rca30_fa24_xor1), .fa_or0(u_rca30_fa24_or0));
  fa fa_u_rca30_fa25_out(.a(a[25]), .b(b[25]), .cin(u_rca30_fa24_or0[0]), .fa_xor1(u_rca30_fa25_xor1), .fa_or0(u_rca30_fa25_or0));
  fa fa_u_rca30_fa26_out(.a(a[26]), .b(b[26]), .cin(u_rca30_fa25_or0[0]), .fa_xor1(u_rca30_fa26_xor1), .fa_or0(u_rca30_fa26_or0));
  fa fa_u_rca30_fa27_out(.a(a[27]), .b(b[27]), .cin(u_rca30_fa26_or0[0]), .fa_xor1(u_rca30_fa27_xor1), .fa_or0(u_rca30_fa27_or0));
  fa fa_u_rca30_fa28_out(.a(a[28]), .b(b[28]), .cin(u_rca30_fa27_or0[0]), .fa_xor1(u_rca30_fa28_xor1), .fa_or0(u_rca30_fa28_or0));
  fa fa_u_rca30_fa29_out(.a(a[29]), .b(b[29]), .cin(u_rca30_fa28_or0[0]), .fa_xor1(u_rca30_fa29_xor1), .fa_or0(u_rca30_fa29_or0));

  assign u_rca30_out[0] = u_rca30_ha_xor0[0];
  assign u_rca30_out[1] = u_rca30_fa1_xor1[0];
  assign u_rca30_out[2] = u_rca30_fa2_xor1[0];
  assign u_rca30_out[3] = u_rca30_fa3_xor1[0];
  assign u_rca30_out[4] = u_rca30_fa4_xor1[0];
  assign u_rca30_out[5] = u_rca30_fa5_xor1[0];
  assign u_rca30_out[6] = u_rca30_fa6_xor1[0];
  assign u_rca30_out[7] = u_rca30_fa7_xor1[0];
  assign u_rca30_out[8] = u_rca30_fa8_xor1[0];
  assign u_rca30_out[9] = u_rca30_fa9_xor1[0];
  assign u_rca30_out[10] = u_rca30_fa10_xor1[0];
  assign u_rca30_out[11] = u_rca30_fa11_xor1[0];
  assign u_rca30_out[12] = u_rca30_fa12_xor1[0];
  assign u_rca30_out[13] = u_rca30_fa13_xor1[0];
  assign u_rca30_out[14] = u_rca30_fa14_xor1[0];
  assign u_rca30_out[15] = u_rca30_fa15_xor1[0];
  assign u_rca30_out[16] = u_rca30_fa16_xor1[0];
  assign u_rca30_out[17] = u_rca30_fa17_xor1[0];
  assign u_rca30_out[18] = u_rca30_fa18_xor1[0];
  assign u_rca30_out[19] = u_rca30_fa19_xor1[0];
  assign u_rca30_out[20] = u_rca30_fa20_xor1[0];
  assign u_rca30_out[21] = u_rca30_fa21_xor1[0];
  assign u_rca30_out[22] = u_rca30_fa22_xor1[0];
  assign u_rca30_out[23] = u_rca30_fa23_xor1[0];
  assign u_rca30_out[24] = u_rca30_fa24_xor1[0];
  assign u_rca30_out[25] = u_rca30_fa25_xor1[0];
  assign u_rca30_out[26] = u_rca30_fa26_xor1[0];
  assign u_rca30_out[27] = u_rca30_fa27_xor1[0];
  assign u_rca30_out[28] = u_rca30_fa28_xor1[0];
  assign u_rca30_out[29] = u_rca30_fa29_xor1[0];
  assign u_rca30_out[30] = u_rca30_fa29_or0[0];
endmodule

module h_u_dadda_rca16(input [15:0] a, input [15:0] b, output [31:0] h_u_dadda_rca16_out);
  wire [0:0] h_u_dadda_rca16_and_13_0;
  wire [0:0] h_u_dadda_rca16_and_12_1;
  wire [0:0] h_u_dadda_rca16_ha0_xor0;
  wire [0:0] h_u_dadda_rca16_ha0_and0;
  wire [0:0] h_u_dadda_rca16_and_14_0;
  wire [0:0] h_u_dadda_rca16_and_13_1;
  wire [0:0] h_u_dadda_rca16_fa0_xor1;
  wire [0:0] h_u_dadda_rca16_fa0_or0;
  wire [0:0] h_u_dadda_rca16_and_12_2;
  wire [0:0] h_u_dadda_rca16_and_11_3;
  wire [0:0] h_u_dadda_rca16_ha1_xor0;
  wire [0:0] h_u_dadda_rca16_ha1_and0;
  wire [0:0] h_u_dadda_rca16_and_15_0;
  wire [0:0] h_u_dadda_rca16_fa1_xor1;
  wire [0:0] h_u_dadda_rca16_fa1_or0;
  wire [0:0] h_u_dadda_rca16_and_14_1;
  wire [0:0] h_u_dadda_rca16_and_13_2;
  wire [0:0] h_u_dadda_rca16_and_12_3;
  wire [0:0] h_u_dadda_rca16_fa2_xor1;
  wire [0:0] h_u_dadda_rca16_fa2_or0;
  wire [0:0] h_u_dadda_rca16_and_11_4;
  wire [0:0] h_u_dadda_rca16_and_10_5;
  wire [0:0] h_u_dadda_rca16_ha2_xor0;
  wire [0:0] h_u_dadda_rca16_ha2_and0;
  wire [0:0] h_u_dadda_rca16_fa3_xor1;
  wire [0:0] h_u_dadda_rca16_fa3_or0;
  wire [0:0] h_u_dadda_rca16_and_15_1;
  wire [0:0] h_u_dadda_rca16_and_14_2;
  wire [0:0] h_u_dadda_rca16_and_13_3;
  wire [0:0] h_u_dadda_rca16_fa4_xor1;
  wire [0:0] h_u_dadda_rca16_fa4_or0;
  wire [0:0] h_u_dadda_rca16_and_12_4;
  wire [0:0] h_u_dadda_rca16_and_11_5;
  wire [0:0] h_u_dadda_rca16_ha3_xor0;
  wire [0:0] h_u_dadda_rca16_ha3_and0;
  wire [0:0] h_u_dadda_rca16_fa5_xor1;
  wire [0:0] h_u_dadda_rca16_fa5_or0;
  wire [0:0] h_u_dadda_rca16_and_15_2;
  wire [0:0] h_u_dadda_rca16_and_14_3;
  wire [0:0] h_u_dadda_rca16_and_13_4;
  wire [0:0] h_u_dadda_rca16_fa6_xor1;
  wire [0:0] h_u_dadda_rca16_fa6_or0;
  wire [0:0] h_u_dadda_rca16_and_15_3;
  wire [0:0] h_u_dadda_rca16_fa7_xor1;
  wire [0:0] h_u_dadda_rca16_fa7_or0;
  wire [0:0] h_u_dadda_rca16_and_4_0;
  wire [0:0] h_u_dadda_rca16_and_3_1;
  wire [0:0] h_u_dadda_rca16_ha4_xor0;
  wire [0:0] h_u_dadda_rca16_ha4_and0;
  wire [0:0] h_u_dadda_rca16_and_5_0;
  wire [0:0] h_u_dadda_rca16_and_4_1;
  wire [0:0] h_u_dadda_rca16_fa8_xor1;
  wire [0:0] h_u_dadda_rca16_fa8_or0;
  wire [0:0] h_u_dadda_rca16_and_3_2;
  wire [0:0] h_u_dadda_rca16_and_2_3;
  wire [0:0] h_u_dadda_rca16_ha5_xor0;
  wire [0:0] h_u_dadda_rca16_ha5_and0;
  wire [0:0] h_u_dadda_rca16_and_6_0;
  wire [0:0] h_u_dadda_rca16_fa9_xor1;
  wire [0:0] h_u_dadda_rca16_fa9_or0;
  wire [0:0] h_u_dadda_rca16_and_5_1;
  wire [0:0] h_u_dadda_rca16_and_4_2;
  wire [0:0] h_u_dadda_rca16_and_3_3;
  wire [0:0] h_u_dadda_rca16_fa10_xor1;
  wire [0:0] h_u_dadda_rca16_fa10_or0;
  wire [0:0] h_u_dadda_rca16_and_2_4;
  wire [0:0] h_u_dadda_rca16_and_1_5;
  wire [0:0] h_u_dadda_rca16_ha6_xor0;
  wire [0:0] h_u_dadda_rca16_ha6_and0;
  wire [0:0] h_u_dadda_rca16_fa11_xor1;
  wire [0:0] h_u_dadda_rca16_fa11_or0;
  wire [0:0] h_u_dadda_rca16_and_7_0;
  wire [0:0] h_u_dadda_rca16_and_6_1;
  wire [0:0] h_u_dadda_rca16_and_5_2;
  wire [0:0] h_u_dadda_rca16_fa12_xor1;
  wire [0:0] h_u_dadda_rca16_fa12_or0;
  wire [0:0] h_u_dadda_rca16_and_4_3;
  wire [0:0] h_u_dadda_rca16_and_3_4;
  wire [0:0] h_u_dadda_rca16_and_2_5;
  wire [0:0] h_u_dadda_rca16_fa13_xor1;
  wire [0:0] h_u_dadda_rca16_fa13_or0;
  wire [0:0] h_u_dadda_rca16_and_1_6;
  wire [0:0] h_u_dadda_rca16_and_0_7;
  wire [0:0] h_u_dadda_rca16_ha7_xor0;
  wire [0:0] h_u_dadda_rca16_ha7_and0;
  wire [0:0] h_u_dadda_rca16_fa14_xor1;
  wire [0:0] h_u_dadda_rca16_fa14_or0;
  wire [0:0] h_u_dadda_rca16_and_8_0;
  wire [0:0] h_u_dadda_rca16_and_7_1;
  wire [0:0] h_u_dadda_rca16_fa15_xor1;
  wire [0:0] h_u_dadda_rca16_fa15_or0;
  wire [0:0] h_u_dadda_rca16_and_6_2;
  wire [0:0] h_u_dadda_rca16_and_5_3;
  wire [0:0] h_u_dadda_rca16_and_4_4;
  wire [0:0] h_u_dadda_rca16_fa16_xor1;
  wire [0:0] h_u_dadda_rca16_fa16_or0;
  wire [0:0] h_u_dadda_rca16_and_3_5;
  wire [0:0] h_u_dadda_rca16_and_2_6;
  wire [0:0] h_u_dadda_rca16_and_1_7;
  wire [0:0] h_u_dadda_rca16_fa17_xor1;
  wire [0:0] h_u_dadda_rca16_fa17_or0;
  wire [0:0] h_u_dadda_rca16_and_0_8;
  wire [0:0] h_u_dadda_rca16_ha8_xor0;
  wire [0:0] h_u_dadda_rca16_ha8_and0;
  wire [0:0] h_u_dadda_rca16_fa18_xor1;
  wire [0:0] h_u_dadda_rca16_fa18_or0;
  wire [0:0] h_u_dadda_rca16_and_9_0;
  wire [0:0] h_u_dadda_rca16_fa19_xor1;
  wire [0:0] h_u_dadda_rca16_fa19_or0;
  wire [0:0] h_u_dadda_rca16_and_8_1;
  wire [0:0] h_u_dadda_rca16_and_7_2;
  wire [0:0] h_u_dadda_rca16_and_6_3;
  wire [0:0] h_u_dadda_rca16_fa20_xor1;
  wire [0:0] h_u_dadda_rca16_fa20_or0;
  wire [0:0] h_u_dadda_rca16_and_5_4;
  wire [0:0] h_u_dadda_rca16_and_4_5;
  wire [0:0] h_u_dadda_rca16_and_3_6;
  wire [0:0] h_u_dadda_rca16_fa21_xor1;
  wire [0:0] h_u_dadda_rca16_fa21_or0;
  wire [0:0] h_u_dadda_rca16_and_2_7;
  wire [0:0] h_u_dadda_rca16_and_1_8;
  wire [0:0] h_u_dadda_rca16_and_0_9;
  wire [0:0] h_u_dadda_rca16_fa22_xor1;
  wire [0:0] h_u_dadda_rca16_fa22_or0;
  wire [0:0] h_u_dadda_rca16_ha9_xor0;
  wire [0:0] h_u_dadda_rca16_ha9_and0;
  wire [0:0] h_u_dadda_rca16_fa23_xor1;
  wire [0:0] h_u_dadda_rca16_fa23_or0;
  wire [0:0] h_u_dadda_rca16_fa24_xor1;
  wire [0:0] h_u_dadda_rca16_fa24_or0;
  wire [0:0] h_u_dadda_rca16_and_10_0;
  wire [0:0] h_u_dadda_rca16_and_9_1;
  wire [0:0] h_u_dadda_rca16_and_8_2;
  wire [0:0] h_u_dadda_rca16_fa25_xor1;
  wire [0:0] h_u_dadda_rca16_fa25_or0;
  wire [0:0] h_u_dadda_rca16_and_7_3;
  wire [0:0] h_u_dadda_rca16_and_6_4;
  wire [0:0] h_u_dadda_rca16_and_5_5;
  wire [0:0] h_u_dadda_rca16_fa26_xor1;
  wire [0:0] h_u_dadda_rca16_fa26_or0;
  wire [0:0] h_u_dadda_rca16_and_4_6;
  wire [0:0] h_u_dadda_rca16_and_3_7;
  wire [0:0] h_u_dadda_rca16_and_2_8;
  wire [0:0] h_u_dadda_rca16_fa27_xor1;
  wire [0:0] h_u_dadda_rca16_fa27_or0;
  wire [0:0] h_u_dadda_rca16_and_1_9;
  wire [0:0] h_u_dadda_rca16_and_0_10;
  wire [0:0] h_u_dadda_rca16_fa28_xor1;
  wire [0:0] h_u_dadda_rca16_fa28_or0;
  wire [0:0] h_u_dadda_rca16_ha10_xor0;
  wire [0:0] h_u_dadda_rca16_ha10_and0;
  wire [0:0] h_u_dadda_rca16_fa29_xor1;
  wire [0:0] h_u_dadda_rca16_fa29_or0;
  wire [0:0] h_u_dadda_rca16_fa30_xor1;
  wire [0:0] h_u_dadda_rca16_fa30_or0;
  wire [0:0] h_u_dadda_rca16_and_11_0;
  wire [0:0] h_u_dadda_rca16_and_10_1;
  wire [0:0] h_u_dadda_rca16_fa31_xor1;
  wire [0:0] h_u_dadda_rca16_fa31_or0;
  wire [0:0] h_u_dadda_rca16_and_9_2;
  wire [0:0] h_u_dadda_rca16_and_8_3;
  wire [0:0] h_u_dadda_rca16_and_7_4;
  wire [0:0] h_u_dadda_rca16_fa32_xor1;
  wire [0:0] h_u_dadda_rca16_fa32_or0;
  wire [0:0] h_u_dadda_rca16_and_6_5;
  wire [0:0] h_u_dadda_rca16_and_5_6;
  wire [0:0] h_u_dadda_rca16_and_4_7;
  wire [0:0] h_u_dadda_rca16_fa33_xor1;
  wire [0:0] h_u_dadda_rca16_fa33_or0;
  wire [0:0] h_u_dadda_rca16_and_3_8;
  wire [0:0] h_u_dadda_rca16_and_2_9;
  wire [0:0] h_u_dadda_rca16_and_1_10;
  wire [0:0] h_u_dadda_rca16_fa34_xor1;
  wire [0:0] h_u_dadda_rca16_fa34_or0;
  wire [0:0] h_u_dadda_rca16_and_0_11;
  wire [0:0] h_u_dadda_rca16_fa35_xor1;
  wire [0:0] h_u_dadda_rca16_fa35_or0;
  wire [0:0] h_u_dadda_rca16_ha11_xor0;
  wire [0:0] h_u_dadda_rca16_ha11_and0;
  wire [0:0] h_u_dadda_rca16_fa36_xor1;
  wire [0:0] h_u_dadda_rca16_fa36_or0;
  wire [0:0] h_u_dadda_rca16_fa37_xor1;
  wire [0:0] h_u_dadda_rca16_fa37_or0;
  wire [0:0] h_u_dadda_rca16_and_12_0;
  wire [0:0] h_u_dadda_rca16_fa38_xor1;
  wire [0:0] h_u_dadda_rca16_fa38_or0;
  wire [0:0] h_u_dadda_rca16_and_11_1;
  wire [0:0] h_u_dadda_rca16_and_10_2;
  wire [0:0] h_u_dadda_rca16_and_9_3;
  wire [0:0] h_u_dadda_rca16_fa39_xor1;
  wire [0:0] h_u_dadda_rca16_fa39_or0;
  wire [0:0] h_u_dadda_rca16_and_8_4;
  wire [0:0] h_u_dadda_rca16_and_7_5;
  wire [0:0] h_u_dadda_rca16_and_6_6;
  wire [0:0] h_u_dadda_rca16_fa40_xor1;
  wire [0:0] h_u_dadda_rca16_fa40_or0;
  wire [0:0] h_u_dadda_rca16_and_5_7;
  wire [0:0] h_u_dadda_rca16_and_4_8;
  wire [0:0] h_u_dadda_rca16_and_3_9;
  wire [0:0] h_u_dadda_rca16_fa41_xor1;
  wire [0:0] h_u_dadda_rca16_fa41_or0;
  wire [0:0] h_u_dadda_rca16_and_2_10;
  wire [0:0] h_u_dadda_rca16_and_1_11;
  wire [0:0] h_u_dadda_rca16_and_0_12;
  wire [0:0] h_u_dadda_rca16_fa42_xor1;
  wire [0:0] h_u_dadda_rca16_fa42_or0;
  wire [0:0] h_u_dadda_rca16_fa43_xor1;
  wire [0:0] h_u_dadda_rca16_fa43_or0;
  wire [0:0] h_u_dadda_rca16_ha12_xor0;
  wire [0:0] h_u_dadda_rca16_ha12_and0;
  wire [0:0] h_u_dadda_rca16_fa44_xor1;
  wire [0:0] h_u_dadda_rca16_fa44_or0;
  wire [0:0] h_u_dadda_rca16_fa45_xor1;
  wire [0:0] h_u_dadda_rca16_fa45_or0;
  wire [0:0] h_u_dadda_rca16_fa46_xor1;
  wire [0:0] h_u_dadda_rca16_fa46_or0;
  wire [0:0] h_u_dadda_rca16_and_11_2;
  wire [0:0] h_u_dadda_rca16_and_10_3;
  wire [0:0] h_u_dadda_rca16_and_9_4;
  wire [0:0] h_u_dadda_rca16_fa47_xor1;
  wire [0:0] h_u_dadda_rca16_fa47_or0;
  wire [0:0] h_u_dadda_rca16_and_8_5;
  wire [0:0] h_u_dadda_rca16_and_7_6;
  wire [0:0] h_u_dadda_rca16_and_6_7;
  wire [0:0] h_u_dadda_rca16_fa48_xor1;
  wire [0:0] h_u_dadda_rca16_fa48_or0;
  wire [0:0] h_u_dadda_rca16_and_5_8;
  wire [0:0] h_u_dadda_rca16_and_4_9;
  wire [0:0] h_u_dadda_rca16_and_3_10;
  wire [0:0] h_u_dadda_rca16_fa49_xor1;
  wire [0:0] h_u_dadda_rca16_fa49_or0;
  wire [0:0] h_u_dadda_rca16_and_2_11;
  wire [0:0] h_u_dadda_rca16_and_1_12;
  wire [0:0] h_u_dadda_rca16_and_0_13;
  wire [0:0] h_u_dadda_rca16_fa50_xor1;
  wire [0:0] h_u_dadda_rca16_fa50_or0;
  wire [0:0] h_u_dadda_rca16_fa51_xor1;
  wire [0:0] h_u_dadda_rca16_fa51_or0;
  wire [0:0] h_u_dadda_rca16_fa52_xor1;
  wire [0:0] h_u_dadda_rca16_fa52_or0;
  wire [0:0] h_u_dadda_rca16_fa53_xor1;
  wire [0:0] h_u_dadda_rca16_fa53_or0;
  wire [0:0] h_u_dadda_rca16_fa54_xor1;
  wire [0:0] h_u_dadda_rca16_fa54_or0;
  wire [0:0] h_u_dadda_rca16_fa55_xor1;
  wire [0:0] h_u_dadda_rca16_fa55_or0;
  wire [0:0] h_u_dadda_rca16_and_10_4;
  wire [0:0] h_u_dadda_rca16_and_9_5;
  wire [0:0] h_u_dadda_rca16_and_8_6;
  wire [0:0] h_u_dadda_rca16_fa56_xor1;
  wire [0:0] h_u_dadda_rca16_fa56_or0;
  wire [0:0] h_u_dadda_rca16_and_7_7;
  wire [0:0] h_u_dadda_rca16_and_6_8;
  wire [0:0] h_u_dadda_rca16_and_5_9;
  wire [0:0] h_u_dadda_rca16_fa57_xor1;
  wire [0:0] h_u_dadda_rca16_fa57_or0;
  wire [0:0] h_u_dadda_rca16_and_4_10;
  wire [0:0] h_u_dadda_rca16_and_3_11;
  wire [0:0] h_u_dadda_rca16_and_2_12;
  wire [0:0] h_u_dadda_rca16_fa58_xor1;
  wire [0:0] h_u_dadda_rca16_fa58_or0;
  wire [0:0] h_u_dadda_rca16_and_1_13;
  wire [0:0] h_u_dadda_rca16_and_0_14;
  wire [0:0] h_u_dadda_rca16_fa59_xor1;
  wire [0:0] h_u_dadda_rca16_fa59_or0;
  wire [0:0] h_u_dadda_rca16_fa60_xor1;
  wire [0:0] h_u_dadda_rca16_fa60_or0;
  wire [0:0] h_u_dadda_rca16_fa61_xor1;
  wire [0:0] h_u_dadda_rca16_fa61_or0;
  wire [0:0] h_u_dadda_rca16_fa62_xor1;
  wire [0:0] h_u_dadda_rca16_fa62_or0;
  wire [0:0] h_u_dadda_rca16_fa63_xor1;
  wire [0:0] h_u_dadda_rca16_fa63_or0;
  wire [0:0] h_u_dadda_rca16_fa64_xor1;
  wire [0:0] h_u_dadda_rca16_fa64_or0;
  wire [0:0] h_u_dadda_rca16_and_9_6;
  wire [0:0] h_u_dadda_rca16_and_8_7;
  wire [0:0] h_u_dadda_rca16_and_7_8;
  wire [0:0] h_u_dadda_rca16_fa65_xor1;
  wire [0:0] h_u_dadda_rca16_fa65_or0;
  wire [0:0] h_u_dadda_rca16_and_6_9;
  wire [0:0] h_u_dadda_rca16_and_5_10;
  wire [0:0] h_u_dadda_rca16_and_4_11;
  wire [0:0] h_u_dadda_rca16_fa66_xor1;
  wire [0:0] h_u_dadda_rca16_fa66_or0;
  wire [0:0] h_u_dadda_rca16_and_3_12;
  wire [0:0] h_u_dadda_rca16_and_2_13;
  wire [0:0] h_u_dadda_rca16_and_1_14;
  wire [0:0] h_u_dadda_rca16_fa67_xor1;
  wire [0:0] h_u_dadda_rca16_fa67_or0;
  wire [0:0] h_u_dadda_rca16_and_0_15;
  wire [0:0] h_u_dadda_rca16_fa68_xor1;
  wire [0:0] h_u_dadda_rca16_fa68_or0;
  wire [0:0] h_u_dadda_rca16_fa69_xor1;
  wire [0:0] h_u_dadda_rca16_fa69_or0;
  wire [0:0] h_u_dadda_rca16_fa70_xor1;
  wire [0:0] h_u_dadda_rca16_fa70_or0;
  wire [0:0] h_u_dadda_rca16_fa71_xor1;
  wire [0:0] h_u_dadda_rca16_fa71_or0;
  wire [0:0] h_u_dadda_rca16_fa72_xor1;
  wire [0:0] h_u_dadda_rca16_fa72_or0;
  wire [0:0] h_u_dadda_rca16_fa73_xor1;
  wire [0:0] h_u_dadda_rca16_fa73_or0;
  wire [0:0] h_u_dadda_rca16_and_10_6;
  wire [0:0] h_u_dadda_rca16_and_9_7;
  wire [0:0] h_u_dadda_rca16_and_8_8;
  wire [0:0] h_u_dadda_rca16_fa74_xor1;
  wire [0:0] h_u_dadda_rca16_fa74_or0;
  wire [0:0] h_u_dadda_rca16_and_7_9;
  wire [0:0] h_u_dadda_rca16_and_6_10;
  wire [0:0] h_u_dadda_rca16_and_5_11;
  wire [0:0] h_u_dadda_rca16_fa75_xor1;
  wire [0:0] h_u_dadda_rca16_fa75_or0;
  wire [0:0] h_u_dadda_rca16_and_4_12;
  wire [0:0] h_u_dadda_rca16_and_3_13;
  wire [0:0] h_u_dadda_rca16_and_2_14;
  wire [0:0] h_u_dadda_rca16_fa76_xor1;
  wire [0:0] h_u_dadda_rca16_fa76_or0;
  wire [0:0] h_u_dadda_rca16_and_1_15;
  wire [0:0] h_u_dadda_rca16_fa77_xor1;
  wire [0:0] h_u_dadda_rca16_fa77_or0;
  wire [0:0] h_u_dadda_rca16_fa78_xor1;
  wire [0:0] h_u_dadda_rca16_fa78_or0;
  wire [0:0] h_u_dadda_rca16_fa79_xor1;
  wire [0:0] h_u_dadda_rca16_fa79_or0;
  wire [0:0] h_u_dadda_rca16_fa80_xor1;
  wire [0:0] h_u_dadda_rca16_fa80_or0;
  wire [0:0] h_u_dadda_rca16_fa81_xor1;
  wire [0:0] h_u_dadda_rca16_fa81_or0;
  wire [0:0] h_u_dadda_rca16_fa82_xor1;
  wire [0:0] h_u_dadda_rca16_fa82_or0;
  wire [0:0] h_u_dadda_rca16_and_12_5;
  wire [0:0] h_u_dadda_rca16_and_11_6;
  wire [0:0] h_u_dadda_rca16_and_10_7;
  wire [0:0] h_u_dadda_rca16_fa83_xor1;
  wire [0:0] h_u_dadda_rca16_fa83_or0;
  wire [0:0] h_u_dadda_rca16_and_9_8;
  wire [0:0] h_u_dadda_rca16_and_8_9;
  wire [0:0] h_u_dadda_rca16_and_7_10;
  wire [0:0] h_u_dadda_rca16_fa84_xor1;
  wire [0:0] h_u_dadda_rca16_fa84_or0;
  wire [0:0] h_u_dadda_rca16_and_6_11;
  wire [0:0] h_u_dadda_rca16_and_5_12;
  wire [0:0] h_u_dadda_rca16_and_4_13;
  wire [0:0] h_u_dadda_rca16_fa85_xor1;
  wire [0:0] h_u_dadda_rca16_fa85_or0;
  wire [0:0] h_u_dadda_rca16_and_3_14;
  wire [0:0] h_u_dadda_rca16_and_2_15;
  wire [0:0] h_u_dadda_rca16_fa86_xor1;
  wire [0:0] h_u_dadda_rca16_fa86_or0;
  wire [0:0] h_u_dadda_rca16_fa87_xor1;
  wire [0:0] h_u_dadda_rca16_fa87_or0;
  wire [0:0] h_u_dadda_rca16_fa88_xor1;
  wire [0:0] h_u_dadda_rca16_fa88_or0;
  wire [0:0] h_u_dadda_rca16_fa89_xor1;
  wire [0:0] h_u_dadda_rca16_fa89_or0;
  wire [0:0] h_u_dadda_rca16_fa90_xor1;
  wire [0:0] h_u_dadda_rca16_fa90_or0;
  wire [0:0] h_u_dadda_rca16_fa91_xor1;
  wire [0:0] h_u_dadda_rca16_fa91_or0;
  wire [0:0] h_u_dadda_rca16_and_14_4;
  wire [0:0] h_u_dadda_rca16_and_13_5;
  wire [0:0] h_u_dadda_rca16_and_12_6;
  wire [0:0] h_u_dadda_rca16_fa92_xor1;
  wire [0:0] h_u_dadda_rca16_fa92_or0;
  wire [0:0] h_u_dadda_rca16_and_11_7;
  wire [0:0] h_u_dadda_rca16_and_10_8;
  wire [0:0] h_u_dadda_rca16_and_9_9;
  wire [0:0] h_u_dadda_rca16_fa93_xor1;
  wire [0:0] h_u_dadda_rca16_fa93_or0;
  wire [0:0] h_u_dadda_rca16_and_8_10;
  wire [0:0] h_u_dadda_rca16_and_7_11;
  wire [0:0] h_u_dadda_rca16_and_6_12;
  wire [0:0] h_u_dadda_rca16_fa94_xor1;
  wire [0:0] h_u_dadda_rca16_fa94_or0;
  wire [0:0] h_u_dadda_rca16_and_5_13;
  wire [0:0] h_u_dadda_rca16_and_4_14;
  wire [0:0] h_u_dadda_rca16_and_3_15;
  wire [0:0] h_u_dadda_rca16_fa95_xor1;
  wire [0:0] h_u_dadda_rca16_fa95_or0;
  wire [0:0] h_u_dadda_rca16_fa96_xor1;
  wire [0:0] h_u_dadda_rca16_fa96_or0;
  wire [0:0] h_u_dadda_rca16_fa97_xor1;
  wire [0:0] h_u_dadda_rca16_fa97_or0;
  wire [0:0] h_u_dadda_rca16_fa98_xor1;
  wire [0:0] h_u_dadda_rca16_fa98_or0;
  wire [0:0] h_u_dadda_rca16_fa99_xor1;
  wire [0:0] h_u_dadda_rca16_fa99_or0;
  wire [0:0] h_u_dadda_rca16_fa100_xor1;
  wire [0:0] h_u_dadda_rca16_fa100_or0;
  wire [0:0] h_u_dadda_rca16_and_15_4;
  wire [0:0] h_u_dadda_rca16_and_14_5;
  wire [0:0] h_u_dadda_rca16_fa101_xor1;
  wire [0:0] h_u_dadda_rca16_fa101_or0;
  wire [0:0] h_u_dadda_rca16_and_13_6;
  wire [0:0] h_u_dadda_rca16_and_12_7;
  wire [0:0] h_u_dadda_rca16_and_11_8;
  wire [0:0] h_u_dadda_rca16_fa102_xor1;
  wire [0:0] h_u_dadda_rca16_fa102_or0;
  wire [0:0] h_u_dadda_rca16_and_10_9;
  wire [0:0] h_u_dadda_rca16_and_9_10;
  wire [0:0] h_u_dadda_rca16_and_8_11;
  wire [0:0] h_u_dadda_rca16_fa103_xor1;
  wire [0:0] h_u_dadda_rca16_fa103_or0;
  wire [0:0] h_u_dadda_rca16_and_7_12;
  wire [0:0] h_u_dadda_rca16_and_6_13;
  wire [0:0] h_u_dadda_rca16_and_5_14;
  wire [0:0] h_u_dadda_rca16_fa104_xor1;
  wire [0:0] h_u_dadda_rca16_fa104_or0;
  wire [0:0] h_u_dadda_rca16_and_4_15;
  wire [0:0] h_u_dadda_rca16_fa105_xor1;
  wire [0:0] h_u_dadda_rca16_fa105_or0;
  wire [0:0] h_u_dadda_rca16_fa106_xor1;
  wire [0:0] h_u_dadda_rca16_fa106_or0;
  wire [0:0] h_u_dadda_rca16_fa107_xor1;
  wire [0:0] h_u_dadda_rca16_fa107_or0;
  wire [0:0] h_u_dadda_rca16_fa108_xor1;
  wire [0:0] h_u_dadda_rca16_fa108_or0;
  wire [0:0] h_u_dadda_rca16_fa109_xor1;
  wire [0:0] h_u_dadda_rca16_fa109_or0;
  wire [0:0] h_u_dadda_rca16_and_15_5;
  wire [0:0] h_u_dadda_rca16_and_14_6;
  wire [0:0] h_u_dadda_rca16_and_13_7;
  wire [0:0] h_u_dadda_rca16_fa110_xor1;
  wire [0:0] h_u_dadda_rca16_fa110_or0;
  wire [0:0] h_u_dadda_rca16_and_12_8;
  wire [0:0] h_u_dadda_rca16_and_11_9;
  wire [0:0] h_u_dadda_rca16_and_10_10;
  wire [0:0] h_u_dadda_rca16_fa111_xor1;
  wire [0:0] h_u_dadda_rca16_fa111_or0;
  wire [0:0] h_u_dadda_rca16_and_9_11;
  wire [0:0] h_u_dadda_rca16_and_8_12;
  wire [0:0] h_u_dadda_rca16_and_7_13;
  wire [0:0] h_u_dadda_rca16_fa112_xor1;
  wire [0:0] h_u_dadda_rca16_fa112_or0;
  wire [0:0] h_u_dadda_rca16_and_6_14;
  wire [0:0] h_u_dadda_rca16_and_5_15;
  wire [0:0] h_u_dadda_rca16_fa113_xor1;
  wire [0:0] h_u_dadda_rca16_fa113_or0;
  wire [0:0] h_u_dadda_rca16_fa114_xor1;
  wire [0:0] h_u_dadda_rca16_fa114_or0;
  wire [0:0] h_u_dadda_rca16_fa115_xor1;
  wire [0:0] h_u_dadda_rca16_fa115_or0;
  wire [0:0] h_u_dadda_rca16_fa116_xor1;
  wire [0:0] h_u_dadda_rca16_fa116_or0;
  wire [0:0] h_u_dadda_rca16_and_15_6;
  wire [0:0] h_u_dadda_rca16_fa117_xor1;
  wire [0:0] h_u_dadda_rca16_fa117_or0;
  wire [0:0] h_u_dadda_rca16_and_14_7;
  wire [0:0] h_u_dadda_rca16_and_13_8;
  wire [0:0] h_u_dadda_rca16_and_12_9;
  wire [0:0] h_u_dadda_rca16_fa118_xor1;
  wire [0:0] h_u_dadda_rca16_fa118_or0;
  wire [0:0] h_u_dadda_rca16_and_11_10;
  wire [0:0] h_u_dadda_rca16_and_10_11;
  wire [0:0] h_u_dadda_rca16_and_9_12;
  wire [0:0] h_u_dadda_rca16_fa119_xor1;
  wire [0:0] h_u_dadda_rca16_fa119_or0;
  wire [0:0] h_u_dadda_rca16_and_8_13;
  wire [0:0] h_u_dadda_rca16_and_7_14;
  wire [0:0] h_u_dadda_rca16_and_6_15;
  wire [0:0] h_u_dadda_rca16_fa120_xor1;
  wire [0:0] h_u_dadda_rca16_fa120_or0;
  wire [0:0] h_u_dadda_rca16_fa121_xor1;
  wire [0:0] h_u_dadda_rca16_fa121_or0;
  wire [0:0] h_u_dadda_rca16_fa122_xor1;
  wire [0:0] h_u_dadda_rca16_fa122_or0;
  wire [0:0] h_u_dadda_rca16_fa123_xor1;
  wire [0:0] h_u_dadda_rca16_fa123_or0;
  wire [0:0] h_u_dadda_rca16_and_15_7;
  wire [0:0] h_u_dadda_rca16_and_14_8;
  wire [0:0] h_u_dadda_rca16_fa124_xor1;
  wire [0:0] h_u_dadda_rca16_fa124_or0;
  wire [0:0] h_u_dadda_rca16_and_13_9;
  wire [0:0] h_u_dadda_rca16_and_12_10;
  wire [0:0] h_u_dadda_rca16_and_11_11;
  wire [0:0] h_u_dadda_rca16_fa125_xor1;
  wire [0:0] h_u_dadda_rca16_fa125_or0;
  wire [0:0] h_u_dadda_rca16_and_10_12;
  wire [0:0] h_u_dadda_rca16_and_9_13;
  wire [0:0] h_u_dadda_rca16_and_8_14;
  wire [0:0] h_u_dadda_rca16_fa126_xor1;
  wire [0:0] h_u_dadda_rca16_fa126_or0;
  wire [0:0] h_u_dadda_rca16_and_7_15;
  wire [0:0] h_u_dadda_rca16_fa127_xor1;
  wire [0:0] h_u_dadda_rca16_fa127_or0;
  wire [0:0] h_u_dadda_rca16_fa128_xor1;
  wire [0:0] h_u_dadda_rca16_fa128_or0;
  wire [0:0] h_u_dadda_rca16_fa129_xor1;
  wire [0:0] h_u_dadda_rca16_fa129_or0;
  wire [0:0] h_u_dadda_rca16_and_15_8;
  wire [0:0] h_u_dadda_rca16_and_14_9;
  wire [0:0] h_u_dadda_rca16_and_13_10;
  wire [0:0] h_u_dadda_rca16_fa130_xor1;
  wire [0:0] h_u_dadda_rca16_fa130_or0;
  wire [0:0] h_u_dadda_rca16_and_12_11;
  wire [0:0] h_u_dadda_rca16_and_11_12;
  wire [0:0] h_u_dadda_rca16_and_10_13;
  wire [0:0] h_u_dadda_rca16_fa131_xor1;
  wire [0:0] h_u_dadda_rca16_fa131_or0;
  wire [0:0] h_u_dadda_rca16_and_9_14;
  wire [0:0] h_u_dadda_rca16_and_8_15;
  wire [0:0] h_u_dadda_rca16_fa132_xor1;
  wire [0:0] h_u_dadda_rca16_fa132_or0;
  wire [0:0] h_u_dadda_rca16_fa133_xor1;
  wire [0:0] h_u_dadda_rca16_fa133_or0;
  wire [0:0] h_u_dadda_rca16_and_15_9;
  wire [0:0] h_u_dadda_rca16_fa134_xor1;
  wire [0:0] h_u_dadda_rca16_fa134_or0;
  wire [0:0] h_u_dadda_rca16_and_14_10;
  wire [0:0] h_u_dadda_rca16_and_13_11;
  wire [0:0] h_u_dadda_rca16_and_12_12;
  wire [0:0] h_u_dadda_rca16_fa135_xor1;
  wire [0:0] h_u_dadda_rca16_fa135_or0;
  wire [0:0] h_u_dadda_rca16_and_11_13;
  wire [0:0] h_u_dadda_rca16_and_10_14;
  wire [0:0] h_u_dadda_rca16_and_9_15;
  wire [0:0] h_u_dadda_rca16_fa136_xor1;
  wire [0:0] h_u_dadda_rca16_fa136_or0;
  wire [0:0] h_u_dadda_rca16_fa137_xor1;
  wire [0:0] h_u_dadda_rca16_fa137_or0;
  wire [0:0] h_u_dadda_rca16_and_15_10;
  wire [0:0] h_u_dadda_rca16_and_14_11;
  wire [0:0] h_u_dadda_rca16_fa138_xor1;
  wire [0:0] h_u_dadda_rca16_fa138_or0;
  wire [0:0] h_u_dadda_rca16_and_13_12;
  wire [0:0] h_u_dadda_rca16_and_12_13;
  wire [0:0] h_u_dadda_rca16_and_11_14;
  wire [0:0] h_u_dadda_rca16_fa139_xor1;
  wire [0:0] h_u_dadda_rca16_fa139_or0;
  wire [0:0] h_u_dadda_rca16_fa140_xor1;
  wire [0:0] h_u_dadda_rca16_fa140_or0;
  wire [0:0] h_u_dadda_rca16_and_15_11;
  wire [0:0] h_u_dadda_rca16_and_14_12;
  wire [0:0] h_u_dadda_rca16_and_13_13;
  wire [0:0] h_u_dadda_rca16_fa141_xor1;
  wire [0:0] h_u_dadda_rca16_fa141_or0;
  wire [0:0] h_u_dadda_rca16_and_15_12;
  wire [0:0] h_u_dadda_rca16_fa142_xor1;
  wire [0:0] h_u_dadda_rca16_fa142_or0;
  wire [0:0] h_u_dadda_rca16_and_3_0;
  wire [0:0] h_u_dadda_rca16_and_2_1;
  wire [0:0] h_u_dadda_rca16_ha13_xor0;
  wire [0:0] h_u_dadda_rca16_ha13_and0;
  wire [0:0] h_u_dadda_rca16_and_2_2;
  wire [0:0] h_u_dadda_rca16_and_1_3;
  wire [0:0] h_u_dadda_rca16_fa143_xor1;
  wire [0:0] h_u_dadda_rca16_fa143_or0;
  wire [0:0] h_u_dadda_rca16_and_1_4;
  wire [0:0] h_u_dadda_rca16_and_0_5;
  wire [0:0] h_u_dadda_rca16_fa144_xor1;
  wire [0:0] h_u_dadda_rca16_fa144_or0;
  wire [0:0] h_u_dadda_rca16_and_0_6;
  wire [0:0] h_u_dadda_rca16_fa145_xor1;
  wire [0:0] h_u_dadda_rca16_fa145_or0;
  wire [0:0] h_u_dadda_rca16_fa146_xor1;
  wire [0:0] h_u_dadda_rca16_fa146_or0;
  wire [0:0] h_u_dadda_rca16_fa147_xor1;
  wire [0:0] h_u_dadda_rca16_fa147_or0;
  wire [0:0] h_u_dadda_rca16_fa148_xor1;
  wire [0:0] h_u_dadda_rca16_fa148_or0;
  wire [0:0] h_u_dadda_rca16_fa149_xor1;
  wire [0:0] h_u_dadda_rca16_fa149_or0;
  wire [0:0] h_u_dadda_rca16_fa150_xor1;
  wire [0:0] h_u_dadda_rca16_fa150_or0;
  wire [0:0] h_u_dadda_rca16_fa151_xor1;
  wire [0:0] h_u_dadda_rca16_fa151_or0;
  wire [0:0] h_u_dadda_rca16_fa152_xor1;
  wire [0:0] h_u_dadda_rca16_fa152_or0;
  wire [0:0] h_u_dadda_rca16_fa153_xor1;
  wire [0:0] h_u_dadda_rca16_fa153_or0;
  wire [0:0] h_u_dadda_rca16_fa154_xor1;
  wire [0:0] h_u_dadda_rca16_fa154_or0;
  wire [0:0] h_u_dadda_rca16_fa155_xor1;
  wire [0:0] h_u_dadda_rca16_fa155_or0;
  wire [0:0] h_u_dadda_rca16_fa156_xor1;
  wire [0:0] h_u_dadda_rca16_fa156_or0;
  wire [0:0] h_u_dadda_rca16_fa157_xor1;
  wire [0:0] h_u_dadda_rca16_fa157_or0;
  wire [0:0] h_u_dadda_rca16_fa158_xor1;
  wire [0:0] h_u_dadda_rca16_fa158_or0;
  wire [0:0] h_u_dadda_rca16_fa159_xor1;
  wire [0:0] h_u_dadda_rca16_fa159_or0;
  wire [0:0] h_u_dadda_rca16_fa160_xor1;
  wire [0:0] h_u_dadda_rca16_fa160_or0;
  wire [0:0] h_u_dadda_rca16_fa161_xor1;
  wire [0:0] h_u_dadda_rca16_fa161_or0;
  wire [0:0] h_u_dadda_rca16_fa162_xor1;
  wire [0:0] h_u_dadda_rca16_fa162_or0;
  wire [0:0] h_u_dadda_rca16_fa163_xor1;
  wire [0:0] h_u_dadda_rca16_fa163_or0;
  wire [0:0] h_u_dadda_rca16_and_10_15;
  wire [0:0] h_u_dadda_rca16_fa164_xor1;
  wire [0:0] h_u_dadda_rca16_fa164_or0;
  wire [0:0] h_u_dadda_rca16_and_12_14;
  wire [0:0] h_u_dadda_rca16_and_11_15;
  wire [0:0] h_u_dadda_rca16_fa165_xor1;
  wire [0:0] h_u_dadda_rca16_fa165_or0;
  wire [0:0] h_u_dadda_rca16_and_14_13;
  wire [0:0] h_u_dadda_rca16_and_13_14;
  wire [0:0] h_u_dadda_rca16_fa166_xor1;
  wire [0:0] h_u_dadda_rca16_fa166_or0;
  wire [0:0] h_u_dadda_rca16_and_15_13;
  wire [0:0] h_u_dadda_rca16_fa167_xor1;
  wire [0:0] h_u_dadda_rca16_fa167_or0;
  wire [0:0] h_u_dadda_rca16_and_2_0;
  wire [0:0] h_u_dadda_rca16_and_1_1;
  wire [0:0] h_u_dadda_rca16_ha14_xor0;
  wire [0:0] h_u_dadda_rca16_ha14_and0;
  wire [0:0] h_u_dadda_rca16_and_1_2;
  wire [0:0] h_u_dadda_rca16_and_0_3;
  wire [0:0] h_u_dadda_rca16_fa168_xor1;
  wire [0:0] h_u_dadda_rca16_fa168_or0;
  wire [0:0] h_u_dadda_rca16_and_0_4;
  wire [0:0] h_u_dadda_rca16_fa169_xor1;
  wire [0:0] h_u_dadda_rca16_fa169_or0;
  wire [0:0] h_u_dadda_rca16_fa170_xor1;
  wire [0:0] h_u_dadda_rca16_fa170_or0;
  wire [0:0] h_u_dadda_rca16_fa171_xor1;
  wire [0:0] h_u_dadda_rca16_fa171_or0;
  wire [0:0] h_u_dadda_rca16_fa172_xor1;
  wire [0:0] h_u_dadda_rca16_fa172_or0;
  wire [0:0] h_u_dadda_rca16_fa173_xor1;
  wire [0:0] h_u_dadda_rca16_fa173_or0;
  wire [0:0] h_u_dadda_rca16_fa174_xor1;
  wire [0:0] h_u_dadda_rca16_fa174_or0;
  wire [0:0] h_u_dadda_rca16_fa175_xor1;
  wire [0:0] h_u_dadda_rca16_fa175_or0;
  wire [0:0] h_u_dadda_rca16_fa176_xor1;
  wire [0:0] h_u_dadda_rca16_fa176_or0;
  wire [0:0] h_u_dadda_rca16_fa177_xor1;
  wire [0:0] h_u_dadda_rca16_fa177_or0;
  wire [0:0] h_u_dadda_rca16_fa178_xor1;
  wire [0:0] h_u_dadda_rca16_fa178_or0;
  wire [0:0] h_u_dadda_rca16_fa179_xor1;
  wire [0:0] h_u_dadda_rca16_fa179_or0;
  wire [0:0] h_u_dadda_rca16_fa180_xor1;
  wire [0:0] h_u_dadda_rca16_fa180_or0;
  wire [0:0] h_u_dadda_rca16_fa181_xor1;
  wire [0:0] h_u_dadda_rca16_fa181_or0;
  wire [0:0] h_u_dadda_rca16_fa182_xor1;
  wire [0:0] h_u_dadda_rca16_fa182_or0;
  wire [0:0] h_u_dadda_rca16_fa183_xor1;
  wire [0:0] h_u_dadda_rca16_fa183_or0;
  wire [0:0] h_u_dadda_rca16_fa184_xor1;
  wire [0:0] h_u_dadda_rca16_fa184_or0;
  wire [0:0] h_u_dadda_rca16_fa185_xor1;
  wire [0:0] h_u_dadda_rca16_fa185_or0;
  wire [0:0] h_u_dadda_rca16_fa186_xor1;
  wire [0:0] h_u_dadda_rca16_fa186_or0;
  wire [0:0] h_u_dadda_rca16_fa187_xor1;
  wire [0:0] h_u_dadda_rca16_fa187_or0;
  wire [0:0] h_u_dadda_rca16_fa188_xor1;
  wire [0:0] h_u_dadda_rca16_fa188_or0;
  wire [0:0] h_u_dadda_rca16_fa189_xor1;
  wire [0:0] h_u_dadda_rca16_fa189_or0;
  wire [0:0] h_u_dadda_rca16_fa190_xor1;
  wire [0:0] h_u_dadda_rca16_fa190_or0;
  wire [0:0] h_u_dadda_rca16_fa191_xor1;
  wire [0:0] h_u_dadda_rca16_fa191_or0;
  wire [0:0] h_u_dadda_rca16_and_12_15;
  wire [0:0] h_u_dadda_rca16_fa192_xor1;
  wire [0:0] h_u_dadda_rca16_fa192_or0;
  wire [0:0] h_u_dadda_rca16_and_14_14;
  wire [0:0] h_u_dadda_rca16_and_13_15;
  wire [0:0] h_u_dadda_rca16_fa193_xor1;
  wire [0:0] h_u_dadda_rca16_fa193_or0;
  wire [0:0] h_u_dadda_rca16_and_15_14;
  wire [0:0] h_u_dadda_rca16_fa194_xor1;
  wire [0:0] h_u_dadda_rca16_fa194_or0;
  wire [0:0] h_u_dadda_rca16_and_0_0;
  wire [0:0] h_u_dadda_rca16_and_1_0;
  wire [0:0] h_u_dadda_rca16_and_0_2;
  wire [0:0] h_u_dadda_rca16_and_14_15;
  wire [0:0] h_u_dadda_rca16_and_0_1;
  wire [0:0] h_u_dadda_rca16_and_15_15;
  wire [29:0] h_u_dadda_rca16_u_rca30_a;
  wire [29:0] h_u_dadda_rca16_u_rca30_b;
  wire [30:0] h_u_dadda_rca16_u_rca30_out;

  and_gate and_gate_h_u_dadda_rca16_and_13_0(.a(a[13]), .b(b[0]), .out(h_u_dadda_rca16_and_13_0));
  and_gate and_gate_h_u_dadda_rca16_and_12_1(.a(a[12]), .b(b[1]), .out(h_u_dadda_rca16_and_12_1));
  ha ha_h_u_dadda_rca16_ha0_out(.a(h_u_dadda_rca16_and_13_0[0]), .b(h_u_dadda_rca16_and_12_1[0]), .ha_xor0(h_u_dadda_rca16_ha0_xor0), .ha_and0(h_u_dadda_rca16_ha0_and0));
  and_gate and_gate_h_u_dadda_rca16_and_14_0(.a(a[14]), .b(b[0]), .out(h_u_dadda_rca16_and_14_0));
  and_gate and_gate_h_u_dadda_rca16_and_13_1(.a(a[13]), .b(b[1]), .out(h_u_dadda_rca16_and_13_1));
  fa fa_h_u_dadda_rca16_fa0_out(.a(h_u_dadda_rca16_ha0_and0[0]), .b(h_u_dadda_rca16_and_14_0[0]), .cin(h_u_dadda_rca16_and_13_1[0]), .fa_xor1(h_u_dadda_rca16_fa0_xor1), .fa_or0(h_u_dadda_rca16_fa0_or0));
  and_gate and_gate_h_u_dadda_rca16_and_12_2(.a(a[12]), .b(b[2]), .out(h_u_dadda_rca16_and_12_2));
  and_gate and_gate_h_u_dadda_rca16_and_11_3(.a(a[11]), .b(b[3]), .out(h_u_dadda_rca16_and_11_3));
  ha ha_h_u_dadda_rca16_ha1_out(.a(h_u_dadda_rca16_and_12_2[0]), .b(h_u_dadda_rca16_and_11_3[0]), .ha_xor0(h_u_dadda_rca16_ha1_xor0), .ha_and0(h_u_dadda_rca16_ha1_and0));
  and_gate and_gate_h_u_dadda_rca16_and_15_0(.a(a[15]), .b(b[0]), .out(h_u_dadda_rca16_and_15_0));
  fa fa_h_u_dadda_rca16_fa1_out(.a(h_u_dadda_rca16_ha1_and0[0]), .b(h_u_dadda_rca16_fa0_or0[0]), .cin(h_u_dadda_rca16_and_15_0[0]), .fa_xor1(h_u_dadda_rca16_fa1_xor1), .fa_or0(h_u_dadda_rca16_fa1_or0));
  and_gate and_gate_h_u_dadda_rca16_and_14_1(.a(a[14]), .b(b[1]), .out(h_u_dadda_rca16_and_14_1));
  and_gate and_gate_h_u_dadda_rca16_and_13_2(.a(a[13]), .b(b[2]), .out(h_u_dadda_rca16_and_13_2));
  and_gate and_gate_h_u_dadda_rca16_and_12_3(.a(a[12]), .b(b[3]), .out(h_u_dadda_rca16_and_12_3));
  fa fa_h_u_dadda_rca16_fa2_out(.a(h_u_dadda_rca16_and_14_1[0]), .b(h_u_dadda_rca16_and_13_2[0]), .cin(h_u_dadda_rca16_and_12_3[0]), .fa_xor1(h_u_dadda_rca16_fa2_xor1), .fa_or0(h_u_dadda_rca16_fa2_or0));
  and_gate and_gate_h_u_dadda_rca16_and_11_4(.a(a[11]), .b(b[4]), .out(h_u_dadda_rca16_and_11_4));
  and_gate and_gate_h_u_dadda_rca16_and_10_5(.a(a[10]), .b(b[5]), .out(h_u_dadda_rca16_and_10_5));
  ha ha_h_u_dadda_rca16_ha2_out(.a(h_u_dadda_rca16_and_11_4[0]), .b(h_u_dadda_rca16_and_10_5[0]), .ha_xor0(h_u_dadda_rca16_ha2_xor0), .ha_and0(h_u_dadda_rca16_ha2_and0));
  fa fa_h_u_dadda_rca16_fa3_out(.a(h_u_dadda_rca16_ha2_and0[0]), .b(h_u_dadda_rca16_fa2_or0[0]), .cin(h_u_dadda_rca16_fa1_or0[0]), .fa_xor1(h_u_dadda_rca16_fa3_xor1), .fa_or0(h_u_dadda_rca16_fa3_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_1(.a(a[15]), .b(b[1]), .out(h_u_dadda_rca16_and_15_1));
  and_gate and_gate_h_u_dadda_rca16_and_14_2(.a(a[14]), .b(b[2]), .out(h_u_dadda_rca16_and_14_2));
  and_gate and_gate_h_u_dadda_rca16_and_13_3(.a(a[13]), .b(b[3]), .out(h_u_dadda_rca16_and_13_3));
  fa fa_h_u_dadda_rca16_fa4_out(.a(h_u_dadda_rca16_and_15_1[0]), .b(h_u_dadda_rca16_and_14_2[0]), .cin(h_u_dadda_rca16_and_13_3[0]), .fa_xor1(h_u_dadda_rca16_fa4_xor1), .fa_or0(h_u_dadda_rca16_fa4_or0));
  and_gate and_gate_h_u_dadda_rca16_and_12_4(.a(a[12]), .b(b[4]), .out(h_u_dadda_rca16_and_12_4));
  and_gate and_gate_h_u_dadda_rca16_and_11_5(.a(a[11]), .b(b[5]), .out(h_u_dadda_rca16_and_11_5));
  ha ha_h_u_dadda_rca16_ha3_out(.a(h_u_dadda_rca16_and_12_4[0]), .b(h_u_dadda_rca16_and_11_5[0]), .ha_xor0(h_u_dadda_rca16_ha3_xor0), .ha_and0(h_u_dadda_rca16_ha3_and0));
  fa fa_h_u_dadda_rca16_fa5_out(.a(h_u_dadda_rca16_ha3_and0[0]), .b(h_u_dadda_rca16_fa4_or0[0]), .cin(h_u_dadda_rca16_fa3_or0[0]), .fa_xor1(h_u_dadda_rca16_fa5_xor1), .fa_or0(h_u_dadda_rca16_fa5_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_2(.a(a[15]), .b(b[2]), .out(h_u_dadda_rca16_and_15_2));
  and_gate and_gate_h_u_dadda_rca16_and_14_3(.a(a[14]), .b(b[3]), .out(h_u_dadda_rca16_and_14_3));
  and_gate and_gate_h_u_dadda_rca16_and_13_4(.a(a[13]), .b(b[4]), .out(h_u_dadda_rca16_and_13_4));
  fa fa_h_u_dadda_rca16_fa6_out(.a(h_u_dadda_rca16_and_15_2[0]), .b(h_u_dadda_rca16_and_14_3[0]), .cin(h_u_dadda_rca16_and_13_4[0]), .fa_xor1(h_u_dadda_rca16_fa6_xor1), .fa_or0(h_u_dadda_rca16_fa6_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_3(.a(a[15]), .b(b[3]), .out(h_u_dadda_rca16_and_15_3));
  fa fa_h_u_dadda_rca16_fa7_out(.a(h_u_dadda_rca16_fa6_or0[0]), .b(h_u_dadda_rca16_fa5_or0[0]), .cin(h_u_dadda_rca16_and_15_3[0]), .fa_xor1(h_u_dadda_rca16_fa7_xor1), .fa_or0(h_u_dadda_rca16_fa7_or0));
  and_gate and_gate_h_u_dadda_rca16_and_4_0(.a(a[4]), .b(b[0]), .out(h_u_dadda_rca16_and_4_0));
  and_gate and_gate_h_u_dadda_rca16_and_3_1(.a(a[3]), .b(b[1]), .out(h_u_dadda_rca16_and_3_1));
  ha ha_h_u_dadda_rca16_ha4_out(.a(h_u_dadda_rca16_and_4_0[0]), .b(h_u_dadda_rca16_and_3_1[0]), .ha_xor0(h_u_dadda_rca16_ha4_xor0), .ha_and0(h_u_dadda_rca16_ha4_and0));
  and_gate and_gate_h_u_dadda_rca16_and_5_0(.a(a[5]), .b(b[0]), .out(h_u_dadda_rca16_and_5_0));
  and_gate and_gate_h_u_dadda_rca16_and_4_1(.a(a[4]), .b(b[1]), .out(h_u_dadda_rca16_and_4_1));
  fa fa_h_u_dadda_rca16_fa8_out(.a(h_u_dadda_rca16_ha4_and0[0]), .b(h_u_dadda_rca16_and_5_0[0]), .cin(h_u_dadda_rca16_and_4_1[0]), .fa_xor1(h_u_dadda_rca16_fa8_xor1), .fa_or0(h_u_dadda_rca16_fa8_or0));
  and_gate and_gate_h_u_dadda_rca16_and_3_2(.a(a[3]), .b(b[2]), .out(h_u_dadda_rca16_and_3_2));
  and_gate and_gate_h_u_dadda_rca16_and_2_3(.a(a[2]), .b(b[3]), .out(h_u_dadda_rca16_and_2_3));
  ha ha_h_u_dadda_rca16_ha5_out(.a(h_u_dadda_rca16_and_3_2[0]), .b(h_u_dadda_rca16_and_2_3[0]), .ha_xor0(h_u_dadda_rca16_ha5_xor0), .ha_and0(h_u_dadda_rca16_ha5_and0));
  and_gate and_gate_h_u_dadda_rca16_and_6_0(.a(a[6]), .b(b[0]), .out(h_u_dadda_rca16_and_6_0));
  fa fa_h_u_dadda_rca16_fa9_out(.a(h_u_dadda_rca16_ha5_and0[0]), .b(h_u_dadda_rca16_fa8_or0[0]), .cin(h_u_dadda_rca16_and_6_0[0]), .fa_xor1(h_u_dadda_rca16_fa9_xor1), .fa_or0(h_u_dadda_rca16_fa9_or0));
  and_gate and_gate_h_u_dadda_rca16_and_5_1(.a(a[5]), .b(b[1]), .out(h_u_dadda_rca16_and_5_1));
  and_gate and_gate_h_u_dadda_rca16_and_4_2(.a(a[4]), .b(b[2]), .out(h_u_dadda_rca16_and_4_2));
  and_gate and_gate_h_u_dadda_rca16_and_3_3(.a(a[3]), .b(b[3]), .out(h_u_dadda_rca16_and_3_3));
  fa fa_h_u_dadda_rca16_fa10_out(.a(h_u_dadda_rca16_and_5_1[0]), .b(h_u_dadda_rca16_and_4_2[0]), .cin(h_u_dadda_rca16_and_3_3[0]), .fa_xor1(h_u_dadda_rca16_fa10_xor1), .fa_or0(h_u_dadda_rca16_fa10_or0));
  and_gate and_gate_h_u_dadda_rca16_and_2_4(.a(a[2]), .b(b[4]), .out(h_u_dadda_rca16_and_2_4));
  and_gate and_gate_h_u_dadda_rca16_and_1_5(.a(a[1]), .b(b[5]), .out(h_u_dadda_rca16_and_1_5));
  ha ha_h_u_dadda_rca16_ha6_out(.a(h_u_dadda_rca16_and_2_4[0]), .b(h_u_dadda_rca16_and_1_5[0]), .ha_xor0(h_u_dadda_rca16_ha6_xor0), .ha_and0(h_u_dadda_rca16_ha6_and0));
  fa fa_h_u_dadda_rca16_fa11_out(.a(h_u_dadda_rca16_ha6_and0[0]), .b(h_u_dadda_rca16_fa10_or0[0]), .cin(h_u_dadda_rca16_fa9_or0[0]), .fa_xor1(h_u_dadda_rca16_fa11_xor1), .fa_or0(h_u_dadda_rca16_fa11_or0));
  and_gate and_gate_h_u_dadda_rca16_and_7_0(.a(a[7]), .b(b[0]), .out(h_u_dadda_rca16_and_7_0));
  and_gate and_gate_h_u_dadda_rca16_and_6_1(.a(a[6]), .b(b[1]), .out(h_u_dadda_rca16_and_6_1));
  and_gate and_gate_h_u_dadda_rca16_and_5_2(.a(a[5]), .b(b[2]), .out(h_u_dadda_rca16_and_5_2));
  fa fa_h_u_dadda_rca16_fa12_out(.a(h_u_dadda_rca16_and_7_0[0]), .b(h_u_dadda_rca16_and_6_1[0]), .cin(h_u_dadda_rca16_and_5_2[0]), .fa_xor1(h_u_dadda_rca16_fa12_xor1), .fa_or0(h_u_dadda_rca16_fa12_or0));
  and_gate and_gate_h_u_dadda_rca16_and_4_3(.a(a[4]), .b(b[3]), .out(h_u_dadda_rca16_and_4_3));
  and_gate and_gate_h_u_dadda_rca16_and_3_4(.a(a[3]), .b(b[4]), .out(h_u_dadda_rca16_and_3_4));
  and_gate and_gate_h_u_dadda_rca16_and_2_5(.a(a[2]), .b(b[5]), .out(h_u_dadda_rca16_and_2_5));
  fa fa_h_u_dadda_rca16_fa13_out(.a(h_u_dadda_rca16_and_4_3[0]), .b(h_u_dadda_rca16_and_3_4[0]), .cin(h_u_dadda_rca16_and_2_5[0]), .fa_xor1(h_u_dadda_rca16_fa13_xor1), .fa_or0(h_u_dadda_rca16_fa13_or0));
  and_gate and_gate_h_u_dadda_rca16_and_1_6(.a(a[1]), .b(b[6]), .out(h_u_dadda_rca16_and_1_6));
  and_gate and_gate_h_u_dadda_rca16_and_0_7(.a(a[0]), .b(b[7]), .out(h_u_dadda_rca16_and_0_7));
  ha ha_h_u_dadda_rca16_ha7_out(.a(h_u_dadda_rca16_and_1_6[0]), .b(h_u_dadda_rca16_and_0_7[0]), .ha_xor0(h_u_dadda_rca16_ha7_xor0), .ha_and0(h_u_dadda_rca16_ha7_and0));
  fa fa_h_u_dadda_rca16_fa14_out(.a(h_u_dadda_rca16_ha7_and0[0]), .b(h_u_dadda_rca16_fa13_or0[0]), .cin(h_u_dadda_rca16_fa12_or0[0]), .fa_xor1(h_u_dadda_rca16_fa14_xor1), .fa_or0(h_u_dadda_rca16_fa14_or0));
  and_gate and_gate_h_u_dadda_rca16_and_8_0(.a(a[8]), .b(b[0]), .out(h_u_dadda_rca16_and_8_0));
  and_gate and_gate_h_u_dadda_rca16_and_7_1(.a(a[7]), .b(b[1]), .out(h_u_dadda_rca16_and_7_1));
  fa fa_h_u_dadda_rca16_fa15_out(.a(h_u_dadda_rca16_fa11_or0[0]), .b(h_u_dadda_rca16_and_8_0[0]), .cin(h_u_dadda_rca16_and_7_1[0]), .fa_xor1(h_u_dadda_rca16_fa15_xor1), .fa_or0(h_u_dadda_rca16_fa15_or0));
  and_gate and_gate_h_u_dadda_rca16_and_6_2(.a(a[6]), .b(b[2]), .out(h_u_dadda_rca16_and_6_2));
  and_gate and_gate_h_u_dadda_rca16_and_5_3(.a(a[5]), .b(b[3]), .out(h_u_dadda_rca16_and_5_3));
  and_gate and_gate_h_u_dadda_rca16_and_4_4(.a(a[4]), .b(b[4]), .out(h_u_dadda_rca16_and_4_4));
  fa fa_h_u_dadda_rca16_fa16_out(.a(h_u_dadda_rca16_and_6_2[0]), .b(h_u_dadda_rca16_and_5_3[0]), .cin(h_u_dadda_rca16_and_4_4[0]), .fa_xor1(h_u_dadda_rca16_fa16_xor1), .fa_or0(h_u_dadda_rca16_fa16_or0));
  and_gate and_gate_h_u_dadda_rca16_and_3_5(.a(a[3]), .b(b[5]), .out(h_u_dadda_rca16_and_3_5));
  and_gate and_gate_h_u_dadda_rca16_and_2_6(.a(a[2]), .b(b[6]), .out(h_u_dadda_rca16_and_2_6));
  and_gate and_gate_h_u_dadda_rca16_and_1_7(.a(a[1]), .b(b[7]), .out(h_u_dadda_rca16_and_1_7));
  fa fa_h_u_dadda_rca16_fa17_out(.a(h_u_dadda_rca16_and_3_5[0]), .b(h_u_dadda_rca16_and_2_6[0]), .cin(h_u_dadda_rca16_and_1_7[0]), .fa_xor1(h_u_dadda_rca16_fa17_xor1), .fa_or0(h_u_dadda_rca16_fa17_or0));
  and_gate and_gate_h_u_dadda_rca16_and_0_8(.a(a[0]), .b(b[8]), .out(h_u_dadda_rca16_and_0_8));
  ha ha_h_u_dadda_rca16_ha8_out(.a(h_u_dadda_rca16_and_0_8[0]), .b(h_u_dadda_rca16_fa14_xor1[0]), .ha_xor0(h_u_dadda_rca16_ha8_xor0), .ha_and0(h_u_dadda_rca16_ha8_and0));
  fa fa_h_u_dadda_rca16_fa18_out(.a(h_u_dadda_rca16_ha8_and0[0]), .b(h_u_dadda_rca16_fa17_or0[0]), .cin(h_u_dadda_rca16_fa16_or0[0]), .fa_xor1(h_u_dadda_rca16_fa18_xor1), .fa_or0(h_u_dadda_rca16_fa18_or0));
  and_gate and_gate_h_u_dadda_rca16_and_9_0(.a(a[9]), .b(b[0]), .out(h_u_dadda_rca16_and_9_0));
  fa fa_h_u_dadda_rca16_fa19_out(.a(h_u_dadda_rca16_fa15_or0[0]), .b(h_u_dadda_rca16_fa14_or0[0]), .cin(h_u_dadda_rca16_and_9_0[0]), .fa_xor1(h_u_dadda_rca16_fa19_xor1), .fa_or0(h_u_dadda_rca16_fa19_or0));
  and_gate and_gate_h_u_dadda_rca16_and_8_1(.a(a[8]), .b(b[1]), .out(h_u_dadda_rca16_and_8_1));
  and_gate and_gate_h_u_dadda_rca16_and_7_2(.a(a[7]), .b(b[2]), .out(h_u_dadda_rca16_and_7_2));
  and_gate and_gate_h_u_dadda_rca16_and_6_3(.a(a[6]), .b(b[3]), .out(h_u_dadda_rca16_and_6_3));
  fa fa_h_u_dadda_rca16_fa20_out(.a(h_u_dadda_rca16_and_8_1[0]), .b(h_u_dadda_rca16_and_7_2[0]), .cin(h_u_dadda_rca16_and_6_3[0]), .fa_xor1(h_u_dadda_rca16_fa20_xor1), .fa_or0(h_u_dadda_rca16_fa20_or0));
  and_gate and_gate_h_u_dadda_rca16_and_5_4(.a(a[5]), .b(b[4]), .out(h_u_dadda_rca16_and_5_4));
  and_gate and_gate_h_u_dadda_rca16_and_4_5(.a(a[4]), .b(b[5]), .out(h_u_dadda_rca16_and_4_5));
  and_gate and_gate_h_u_dadda_rca16_and_3_6(.a(a[3]), .b(b[6]), .out(h_u_dadda_rca16_and_3_6));
  fa fa_h_u_dadda_rca16_fa21_out(.a(h_u_dadda_rca16_and_5_4[0]), .b(h_u_dadda_rca16_and_4_5[0]), .cin(h_u_dadda_rca16_and_3_6[0]), .fa_xor1(h_u_dadda_rca16_fa21_xor1), .fa_or0(h_u_dadda_rca16_fa21_or0));
  and_gate and_gate_h_u_dadda_rca16_and_2_7(.a(a[2]), .b(b[7]), .out(h_u_dadda_rca16_and_2_7));
  and_gate and_gate_h_u_dadda_rca16_and_1_8(.a(a[1]), .b(b[8]), .out(h_u_dadda_rca16_and_1_8));
  and_gate and_gate_h_u_dadda_rca16_and_0_9(.a(a[0]), .b(b[9]), .out(h_u_dadda_rca16_and_0_9));
  fa fa_h_u_dadda_rca16_fa22_out(.a(h_u_dadda_rca16_and_2_7[0]), .b(h_u_dadda_rca16_and_1_8[0]), .cin(h_u_dadda_rca16_and_0_9[0]), .fa_xor1(h_u_dadda_rca16_fa22_xor1), .fa_or0(h_u_dadda_rca16_fa22_or0));
  ha ha_h_u_dadda_rca16_ha9_out(.a(h_u_dadda_rca16_fa18_xor1[0]), .b(h_u_dadda_rca16_fa19_xor1[0]), .ha_xor0(h_u_dadda_rca16_ha9_xor0), .ha_and0(h_u_dadda_rca16_ha9_and0));
  fa fa_h_u_dadda_rca16_fa23_out(.a(h_u_dadda_rca16_ha9_and0[0]), .b(h_u_dadda_rca16_fa22_or0[0]), .cin(h_u_dadda_rca16_fa21_or0[0]), .fa_xor1(h_u_dadda_rca16_fa23_xor1), .fa_or0(h_u_dadda_rca16_fa23_or0));
  fa fa_h_u_dadda_rca16_fa24_out(.a(h_u_dadda_rca16_fa20_or0[0]), .b(h_u_dadda_rca16_fa19_or0[0]), .cin(h_u_dadda_rca16_fa18_or0[0]), .fa_xor1(h_u_dadda_rca16_fa24_xor1), .fa_or0(h_u_dadda_rca16_fa24_or0));
  and_gate and_gate_h_u_dadda_rca16_and_10_0(.a(a[10]), .b(b[0]), .out(h_u_dadda_rca16_and_10_0));
  and_gate and_gate_h_u_dadda_rca16_and_9_1(.a(a[9]), .b(b[1]), .out(h_u_dadda_rca16_and_9_1));
  and_gate and_gate_h_u_dadda_rca16_and_8_2(.a(a[8]), .b(b[2]), .out(h_u_dadda_rca16_and_8_2));
  fa fa_h_u_dadda_rca16_fa25_out(.a(h_u_dadda_rca16_and_10_0[0]), .b(h_u_dadda_rca16_and_9_1[0]), .cin(h_u_dadda_rca16_and_8_2[0]), .fa_xor1(h_u_dadda_rca16_fa25_xor1), .fa_or0(h_u_dadda_rca16_fa25_or0));
  and_gate and_gate_h_u_dadda_rca16_and_7_3(.a(a[7]), .b(b[3]), .out(h_u_dadda_rca16_and_7_3));
  and_gate and_gate_h_u_dadda_rca16_and_6_4(.a(a[6]), .b(b[4]), .out(h_u_dadda_rca16_and_6_4));
  and_gate and_gate_h_u_dadda_rca16_and_5_5(.a(a[5]), .b(b[5]), .out(h_u_dadda_rca16_and_5_5));
  fa fa_h_u_dadda_rca16_fa26_out(.a(h_u_dadda_rca16_and_7_3[0]), .b(h_u_dadda_rca16_and_6_4[0]), .cin(h_u_dadda_rca16_and_5_5[0]), .fa_xor1(h_u_dadda_rca16_fa26_xor1), .fa_or0(h_u_dadda_rca16_fa26_or0));
  and_gate and_gate_h_u_dadda_rca16_and_4_6(.a(a[4]), .b(b[6]), .out(h_u_dadda_rca16_and_4_6));
  and_gate and_gate_h_u_dadda_rca16_and_3_7(.a(a[3]), .b(b[7]), .out(h_u_dadda_rca16_and_3_7));
  and_gate and_gate_h_u_dadda_rca16_and_2_8(.a(a[2]), .b(b[8]), .out(h_u_dadda_rca16_and_2_8));
  fa fa_h_u_dadda_rca16_fa27_out(.a(h_u_dadda_rca16_and_4_6[0]), .b(h_u_dadda_rca16_and_3_7[0]), .cin(h_u_dadda_rca16_and_2_8[0]), .fa_xor1(h_u_dadda_rca16_fa27_xor1), .fa_or0(h_u_dadda_rca16_fa27_or0));
  and_gate and_gate_h_u_dadda_rca16_and_1_9(.a(a[1]), .b(b[9]), .out(h_u_dadda_rca16_and_1_9));
  and_gate and_gate_h_u_dadda_rca16_and_0_10(.a(a[0]), .b(b[10]), .out(h_u_dadda_rca16_and_0_10));
  fa fa_h_u_dadda_rca16_fa28_out(.a(h_u_dadda_rca16_and_1_9[0]), .b(h_u_dadda_rca16_and_0_10[0]), .cin(h_u_dadda_rca16_fa23_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa28_xor1), .fa_or0(h_u_dadda_rca16_fa28_or0));
  ha ha_h_u_dadda_rca16_ha10_out(.a(h_u_dadda_rca16_fa24_xor1[0]), .b(h_u_dadda_rca16_fa25_xor1[0]), .ha_xor0(h_u_dadda_rca16_ha10_xor0), .ha_and0(h_u_dadda_rca16_ha10_and0));
  fa fa_h_u_dadda_rca16_fa29_out(.a(h_u_dadda_rca16_ha10_and0[0]), .b(h_u_dadda_rca16_fa28_or0[0]), .cin(h_u_dadda_rca16_fa27_or0[0]), .fa_xor1(h_u_dadda_rca16_fa29_xor1), .fa_or0(h_u_dadda_rca16_fa29_or0));
  fa fa_h_u_dadda_rca16_fa30_out(.a(h_u_dadda_rca16_fa26_or0[0]), .b(h_u_dadda_rca16_fa25_or0[0]), .cin(h_u_dadda_rca16_fa24_or0[0]), .fa_xor1(h_u_dadda_rca16_fa30_xor1), .fa_or0(h_u_dadda_rca16_fa30_or0));
  and_gate and_gate_h_u_dadda_rca16_and_11_0(.a(a[11]), .b(b[0]), .out(h_u_dadda_rca16_and_11_0));
  and_gate and_gate_h_u_dadda_rca16_and_10_1(.a(a[10]), .b(b[1]), .out(h_u_dadda_rca16_and_10_1));
  fa fa_h_u_dadda_rca16_fa31_out(.a(h_u_dadda_rca16_fa23_or0[0]), .b(h_u_dadda_rca16_and_11_0[0]), .cin(h_u_dadda_rca16_and_10_1[0]), .fa_xor1(h_u_dadda_rca16_fa31_xor1), .fa_or0(h_u_dadda_rca16_fa31_or0));
  and_gate and_gate_h_u_dadda_rca16_and_9_2(.a(a[9]), .b(b[2]), .out(h_u_dadda_rca16_and_9_2));
  and_gate and_gate_h_u_dadda_rca16_and_8_3(.a(a[8]), .b(b[3]), .out(h_u_dadda_rca16_and_8_3));
  and_gate and_gate_h_u_dadda_rca16_and_7_4(.a(a[7]), .b(b[4]), .out(h_u_dadda_rca16_and_7_4));
  fa fa_h_u_dadda_rca16_fa32_out(.a(h_u_dadda_rca16_and_9_2[0]), .b(h_u_dadda_rca16_and_8_3[0]), .cin(h_u_dadda_rca16_and_7_4[0]), .fa_xor1(h_u_dadda_rca16_fa32_xor1), .fa_or0(h_u_dadda_rca16_fa32_or0));
  and_gate and_gate_h_u_dadda_rca16_and_6_5(.a(a[6]), .b(b[5]), .out(h_u_dadda_rca16_and_6_5));
  and_gate and_gate_h_u_dadda_rca16_and_5_6(.a(a[5]), .b(b[6]), .out(h_u_dadda_rca16_and_5_6));
  and_gate and_gate_h_u_dadda_rca16_and_4_7(.a(a[4]), .b(b[7]), .out(h_u_dadda_rca16_and_4_7));
  fa fa_h_u_dadda_rca16_fa33_out(.a(h_u_dadda_rca16_and_6_5[0]), .b(h_u_dadda_rca16_and_5_6[0]), .cin(h_u_dadda_rca16_and_4_7[0]), .fa_xor1(h_u_dadda_rca16_fa33_xor1), .fa_or0(h_u_dadda_rca16_fa33_or0));
  and_gate and_gate_h_u_dadda_rca16_and_3_8(.a(a[3]), .b(b[8]), .out(h_u_dadda_rca16_and_3_8));
  and_gate and_gate_h_u_dadda_rca16_and_2_9(.a(a[2]), .b(b[9]), .out(h_u_dadda_rca16_and_2_9));
  and_gate and_gate_h_u_dadda_rca16_and_1_10(.a(a[1]), .b(b[10]), .out(h_u_dadda_rca16_and_1_10));
  fa fa_h_u_dadda_rca16_fa34_out(.a(h_u_dadda_rca16_and_3_8[0]), .b(h_u_dadda_rca16_and_2_9[0]), .cin(h_u_dadda_rca16_and_1_10[0]), .fa_xor1(h_u_dadda_rca16_fa34_xor1), .fa_or0(h_u_dadda_rca16_fa34_or0));
  and_gate and_gate_h_u_dadda_rca16_and_0_11(.a(a[0]), .b(b[11]), .out(h_u_dadda_rca16_and_0_11));
  fa fa_h_u_dadda_rca16_fa35_out(.a(h_u_dadda_rca16_and_0_11[0]), .b(h_u_dadda_rca16_fa29_xor1[0]), .cin(h_u_dadda_rca16_fa30_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa35_xor1), .fa_or0(h_u_dadda_rca16_fa35_or0));
  ha ha_h_u_dadda_rca16_ha11_out(.a(h_u_dadda_rca16_fa31_xor1[0]), .b(h_u_dadda_rca16_fa32_xor1[0]), .ha_xor0(h_u_dadda_rca16_ha11_xor0), .ha_and0(h_u_dadda_rca16_ha11_and0));
  fa fa_h_u_dadda_rca16_fa36_out(.a(h_u_dadda_rca16_ha11_and0[0]), .b(h_u_dadda_rca16_fa35_or0[0]), .cin(h_u_dadda_rca16_fa34_or0[0]), .fa_xor1(h_u_dadda_rca16_fa36_xor1), .fa_or0(h_u_dadda_rca16_fa36_or0));
  fa fa_h_u_dadda_rca16_fa37_out(.a(h_u_dadda_rca16_fa33_or0[0]), .b(h_u_dadda_rca16_fa32_or0[0]), .cin(h_u_dadda_rca16_fa31_or0[0]), .fa_xor1(h_u_dadda_rca16_fa37_xor1), .fa_or0(h_u_dadda_rca16_fa37_or0));
  and_gate and_gate_h_u_dadda_rca16_and_12_0(.a(a[12]), .b(b[0]), .out(h_u_dadda_rca16_and_12_0));
  fa fa_h_u_dadda_rca16_fa38_out(.a(h_u_dadda_rca16_fa30_or0[0]), .b(h_u_dadda_rca16_fa29_or0[0]), .cin(h_u_dadda_rca16_and_12_0[0]), .fa_xor1(h_u_dadda_rca16_fa38_xor1), .fa_or0(h_u_dadda_rca16_fa38_or0));
  and_gate and_gate_h_u_dadda_rca16_and_11_1(.a(a[11]), .b(b[1]), .out(h_u_dadda_rca16_and_11_1));
  and_gate and_gate_h_u_dadda_rca16_and_10_2(.a(a[10]), .b(b[2]), .out(h_u_dadda_rca16_and_10_2));
  and_gate and_gate_h_u_dadda_rca16_and_9_3(.a(a[9]), .b(b[3]), .out(h_u_dadda_rca16_and_9_3));
  fa fa_h_u_dadda_rca16_fa39_out(.a(h_u_dadda_rca16_and_11_1[0]), .b(h_u_dadda_rca16_and_10_2[0]), .cin(h_u_dadda_rca16_and_9_3[0]), .fa_xor1(h_u_dadda_rca16_fa39_xor1), .fa_or0(h_u_dadda_rca16_fa39_or0));
  and_gate and_gate_h_u_dadda_rca16_and_8_4(.a(a[8]), .b(b[4]), .out(h_u_dadda_rca16_and_8_4));
  and_gate and_gate_h_u_dadda_rca16_and_7_5(.a(a[7]), .b(b[5]), .out(h_u_dadda_rca16_and_7_5));
  and_gate and_gate_h_u_dadda_rca16_and_6_6(.a(a[6]), .b(b[6]), .out(h_u_dadda_rca16_and_6_6));
  fa fa_h_u_dadda_rca16_fa40_out(.a(h_u_dadda_rca16_and_8_4[0]), .b(h_u_dadda_rca16_and_7_5[0]), .cin(h_u_dadda_rca16_and_6_6[0]), .fa_xor1(h_u_dadda_rca16_fa40_xor1), .fa_or0(h_u_dadda_rca16_fa40_or0));
  and_gate and_gate_h_u_dadda_rca16_and_5_7(.a(a[5]), .b(b[7]), .out(h_u_dadda_rca16_and_5_7));
  and_gate and_gate_h_u_dadda_rca16_and_4_8(.a(a[4]), .b(b[8]), .out(h_u_dadda_rca16_and_4_8));
  and_gate and_gate_h_u_dadda_rca16_and_3_9(.a(a[3]), .b(b[9]), .out(h_u_dadda_rca16_and_3_9));
  fa fa_h_u_dadda_rca16_fa41_out(.a(h_u_dadda_rca16_and_5_7[0]), .b(h_u_dadda_rca16_and_4_8[0]), .cin(h_u_dadda_rca16_and_3_9[0]), .fa_xor1(h_u_dadda_rca16_fa41_xor1), .fa_or0(h_u_dadda_rca16_fa41_or0));
  and_gate and_gate_h_u_dadda_rca16_and_2_10(.a(a[2]), .b(b[10]), .out(h_u_dadda_rca16_and_2_10));
  and_gate and_gate_h_u_dadda_rca16_and_1_11(.a(a[1]), .b(b[11]), .out(h_u_dadda_rca16_and_1_11));
  and_gate and_gate_h_u_dadda_rca16_and_0_12(.a(a[0]), .b(b[12]), .out(h_u_dadda_rca16_and_0_12));
  fa fa_h_u_dadda_rca16_fa42_out(.a(h_u_dadda_rca16_and_2_10[0]), .b(h_u_dadda_rca16_and_1_11[0]), .cin(h_u_dadda_rca16_and_0_12[0]), .fa_xor1(h_u_dadda_rca16_fa42_xor1), .fa_or0(h_u_dadda_rca16_fa42_or0));
  fa fa_h_u_dadda_rca16_fa43_out(.a(h_u_dadda_rca16_fa36_xor1[0]), .b(h_u_dadda_rca16_fa37_xor1[0]), .cin(h_u_dadda_rca16_fa38_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa43_xor1), .fa_or0(h_u_dadda_rca16_fa43_or0));
  ha ha_h_u_dadda_rca16_ha12_out(.a(h_u_dadda_rca16_fa39_xor1[0]), .b(h_u_dadda_rca16_fa40_xor1[0]), .ha_xor0(h_u_dadda_rca16_ha12_xor0), .ha_and0(h_u_dadda_rca16_ha12_and0));
  fa fa_h_u_dadda_rca16_fa44_out(.a(h_u_dadda_rca16_ha12_and0[0]), .b(h_u_dadda_rca16_fa43_or0[0]), .cin(h_u_dadda_rca16_fa42_or0[0]), .fa_xor1(h_u_dadda_rca16_fa44_xor1), .fa_or0(h_u_dadda_rca16_fa44_or0));
  fa fa_h_u_dadda_rca16_fa45_out(.a(h_u_dadda_rca16_fa41_or0[0]), .b(h_u_dadda_rca16_fa40_or0[0]), .cin(h_u_dadda_rca16_fa39_or0[0]), .fa_xor1(h_u_dadda_rca16_fa45_xor1), .fa_or0(h_u_dadda_rca16_fa45_or0));
  fa fa_h_u_dadda_rca16_fa46_out(.a(h_u_dadda_rca16_fa38_or0[0]), .b(h_u_dadda_rca16_fa37_or0[0]), .cin(h_u_dadda_rca16_fa36_or0[0]), .fa_xor1(h_u_dadda_rca16_fa46_xor1), .fa_or0(h_u_dadda_rca16_fa46_or0));
  and_gate and_gate_h_u_dadda_rca16_and_11_2(.a(a[11]), .b(b[2]), .out(h_u_dadda_rca16_and_11_2));
  and_gate and_gate_h_u_dadda_rca16_and_10_3(.a(a[10]), .b(b[3]), .out(h_u_dadda_rca16_and_10_3));
  and_gate and_gate_h_u_dadda_rca16_and_9_4(.a(a[9]), .b(b[4]), .out(h_u_dadda_rca16_and_9_4));
  fa fa_h_u_dadda_rca16_fa47_out(.a(h_u_dadda_rca16_and_11_2[0]), .b(h_u_dadda_rca16_and_10_3[0]), .cin(h_u_dadda_rca16_and_9_4[0]), .fa_xor1(h_u_dadda_rca16_fa47_xor1), .fa_or0(h_u_dadda_rca16_fa47_or0));
  and_gate and_gate_h_u_dadda_rca16_and_8_5(.a(a[8]), .b(b[5]), .out(h_u_dadda_rca16_and_8_5));
  and_gate and_gate_h_u_dadda_rca16_and_7_6(.a(a[7]), .b(b[6]), .out(h_u_dadda_rca16_and_7_6));
  and_gate and_gate_h_u_dadda_rca16_and_6_7(.a(a[6]), .b(b[7]), .out(h_u_dadda_rca16_and_6_7));
  fa fa_h_u_dadda_rca16_fa48_out(.a(h_u_dadda_rca16_and_8_5[0]), .b(h_u_dadda_rca16_and_7_6[0]), .cin(h_u_dadda_rca16_and_6_7[0]), .fa_xor1(h_u_dadda_rca16_fa48_xor1), .fa_or0(h_u_dadda_rca16_fa48_or0));
  and_gate and_gate_h_u_dadda_rca16_and_5_8(.a(a[5]), .b(b[8]), .out(h_u_dadda_rca16_and_5_8));
  and_gate and_gate_h_u_dadda_rca16_and_4_9(.a(a[4]), .b(b[9]), .out(h_u_dadda_rca16_and_4_9));
  and_gate and_gate_h_u_dadda_rca16_and_3_10(.a(a[3]), .b(b[10]), .out(h_u_dadda_rca16_and_3_10));
  fa fa_h_u_dadda_rca16_fa49_out(.a(h_u_dadda_rca16_and_5_8[0]), .b(h_u_dadda_rca16_and_4_9[0]), .cin(h_u_dadda_rca16_and_3_10[0]), .fa_xor1(h_u_dadda_rca16_fa49_xor1), .fa_or0(h_u_dadda_rca16_fa49_or0));
  and_gate and_gate_h_u_dadda_rca16_and_2_11(.a(a[2]), .b(b[11]), .out(h_u_dadda_rca16_and_2_11));
  and_gate and_gate_h_u_dadda_rca16_and_1_12(.a(a[1]), .b(b[12]), .out(h_u_dadda_rca16_and_1_12));
  and_gate and_gate_h_u_dadda_rca16_and_0_13(.a(a[0]), .b(b[13]), .out(h_u_dadda_rca16_and_0_13));
  fa fa_h_u_dadda_rca16_fa50_out(.a(h_u_dadda_rca16_and_2_11[0]), .b(h_u_dadda_rca16_and_1_12[0]), .cin(h_u_dadda_rca16_and_0_13[0]), .fa_xor1(h_u_dadda_rca16_fa50_xor1), .fa_or0(h_u_dadda_rca16_fa50_or0));
  fa fa_h_u_dadda_rca16_fa51_out(.a(h_u_dadda_rca16_ha0_xor0[0]), .b(h_u_dadda_rca16_fa44_xor1[0]), .cin(h_u_dadda_rca16_fa45_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa51_xor1), .fa_or0(h_u_dadda_rca16_fa51_or0));
  fa fa_h_u_dadda_rca16_fa52_out(.a(h_u_dadda_rca16_fa46_xor1[0]), .b(h_u_dadda_rca16_fa47_xor1[0]), .cin(h_u_dadda_rca16_fa48_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa52_xor1), .fa_or0(h_u_dadda_rca16_fa52_or0));
  fa fa_h_u_dadda_rca16_fa53_out(.a(h_u_dadda_rca16_fa52_or0[0]), .b(h_u_dadda_rca16_fa51_or0[0]), .cin(h_u_dadda_rca16_fa50_or0[0]), .fa_xor1(h_u_dadda_rca16_fa53_xor1), .fa_or0(h_u_dadda_rca16_fa53_or0));
  fa fa_h_u_dadda_rca16_fa54_out(.a(h_u_dadda_rca16_fa49_or0[0]), .b(h_u_dadda_rca16_fa48_or0[0]), .cin(h_u_dadda_rca16_fa47_or0[0]), .fa_xor1(h_u_dadda_rca16_fa54_xor1), .fa_or0(h_u_dadda_rca16_fa54_or0));
  fa fa_h_u_dadda_rca16_fa55_out(.a(h_u_dadda_rca16_fa46_or0[0]), .b(h_u_dadda_rca16_fa45_or0[0]), .cin(h_u_dadda_rca16_fa44_or0[0]), .fa_xor1(h_u_dadda_rca16_fa55_xor1), .fa_or0(h_u_dadda_rca16_fa55_or0));
  and_gate and_gate_h_u_dadda_rca16_and_10_4(.a(a[10]), .b(b[4]), .out(h_u_dadda_rca16_and_10_4));
  and_gate and_gate_h_u_dadda_rca16_and_9_5(.a(a[9]), .b(b[5]), .out(h_u_dadda_rca16_and_9_5));
  and_gate and_gate_h_u_dadda_rca16_and_8_6(.a(a[8]), .b(b[6]), .out(h_u_dadda_rca16_and_8_6));
  fa fa_h_u_dadda_rca16_fa56_out(.a(h_u_dadda_rca16_and_10_4[0]), .b(h_u_dadda_rca16_and_9_5[0]), .cin(h_u_dadda_rca16_and_8_6[0]), .fa_xor1(h_u_dadda_rca16_fa56_xor1), .fa_or0(h_u_dadda_rca16_fa56_or0));
  and_gate and_gate_h_u_dadda_rca16_and_7_7(.a(a[7]), .b(b[7]), .out(h_u_dadda_rca16_and_7_7));
  and_gate and_gate_h_u_dadda_rca16_and_6_8(.a(a[6]), .b(b[8]), .out(h_u_dadda_rca16_and_6_8));
  and_gate and_gate_h_u_dadda_rca16_and_5_9(.a(a[5]), .b(b[9]), .out(h_u_dadda_rca16_and_5_9));
  fa fa_h_u_dadda_rca16_fa57_out(.a(h_u_dadda_rca16_and_7_7[0]), .b(h_u_dadda_rca16_and_6_8[0]), .cin(h_u_dadda_rca16_and_5_9[0]), .fa_xor1(h_u_dadda_rca16_fa57_xor1), .fa_or0(h_u_dadda_rca16_fa57_or0));
  and_gate and_gate_h_u_dadda_rca16_and_4_10(.a(a[4]), .b(b[10]), .out(h_u_dadda_rca16_and_4_10));
  and_gate and_gate_h_u_dadda_rca16_and_3_11(.a(a[3]), .b(b[11]), .out(h_u_dadda_rca16_and_3_11));
  and_gate and_gate_h_u_dadda_rca16_and_2_12(.a(a[2]), .b(b[12]), .out(h_u_dadda_rca16_and_2_12));
  fa fa_h_u_dadda_rca16_fa58_out(.a(h_u_dadda_rca16_and_4_10[0]), .b(h_u_dadda_rca16_and_3_11[0]), .cin(h_u_dadda_rca16_and_2_12[0]), .fa_xor1(h_u_dadda_rca16_fa58_xor1), .fa_or0(h_u_dadda_rca16_fa58_or0));
  and_gate and_gate_h_u_dadda_rca16_and_1_13(.a(a[1]), .b(b[13]), .out(h_u_dadda_rca16_and_1_13));
  and_gate and_gate_h_u_dadda_rca16_and_0_14(.a(a[0]), .b(b[14]), .out(h_u_dadda_rca16_and_0_14));
  fa fa_h_u_dadda_rca16_fa59_out(.a(h_u_dadda_rca16_and_1_13[0]), .b(h_u_dadda_rca16_and_0_14[0]), .cin(h_u_dadda_rca16_fa0_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa59_xor1), .fa_or0(h_u_dadda_rca16_fa59_or0));
  fa fa_h_u_dadda_rca16_fa60_out(.a(h_u_dadda_rca16_ha1_xor0[0]), .b(h_u_dadda_rca16_fa53_xor1[0]), .cin(h_u_dadda_rca16_fa54_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa60_xor1), .fa_or0(h_u_dadda_rca16_fa60_or0));
  fa fa_h_u_dadda_rca16_fa61_out(.a(h_u_dadda_rca16_fa55_xor1[0]), .b(h_u_dadda_rca16_fa56_xor1[0]), .cin(h_u_dadda_rca16_fa57_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa61_xor1), .fa_or0(h_u_dadda_rca16_fa61_or0));
  fa fa_h_u_dadda_rca16_fa62_out(.a(h_u_dadda_rca16_fa61_or0[0]), .b(h_u_dadda_rca16_fa60_or0[0]), .cin(h_u_dadda_rca16_fa59_or0[0]), .fa_xor1(h_u_dadda_rca16_fa62_xor1), .fa_or0(h_u_dadda_rca16_fa62_or0));
  fa fa_h_u_dadda_rca16_fa63_out(.a(h_u_dadda_rca16_fa58_or0[0]), .b(h_u_dadda_rca16_fa57_or0[0]), .cin(h_u_dadda_rca16_fa56_or0[0]), .fa_xor1(h_u_dadda_rca16_fa63_xor1), .fa_or0(h_u_dadda_rca16_fa63_or0));
  fa fa_h_u_dadda_rca16_fa64_out(.a(h_u_dadda_rca16_fa55_or0[0]), .b(h_u_dadda_rca16_fa54_or0[0]), .cin(h_u_dadda_rca16_fa53_or0[0]), .fa_xor1(h_u_dadda_rca16_fa64_xor1), .fa_or0(h_u_dadda_rca16_fa64_or0));
  and_gate and_gate_h_u_dadda_rca16_and_9_6(.a(a[9]), .b(b[6]), .out(h_u_dadda_rca16_and_9_6));
  and_gate and_gate_h_u_dadda_rca16_and_8_7(.a(a[8]), .b(b[7]), .out(h_u_dadda_rca16_and_8_7));
  and_gate and_gate_h_u_dadda_rca16_and_7_8(.a(a[7]), .b(b[8]), .out(h_u_dadda_rca16_and_7_8));
  fa fa_h_u_dadda_rca16_fa65_out(.a(h_u_dadda_rca16_and_9_6[0]), .b(h_u_dadda_rca16_and_8_7[0]), .cin(h_u_dadda_rca16_and_7_8[0]), .fa_xor1(h_u_dadda_rca16_fa65_xor1), .fa_or0(h_u_dadda_rca16_fa65_or0));
  and_gate and_gate_h_u_dadda_rca16_and_6_9(.a(a[6]), .b(b[9]), .out(h_u_dadda_rca16_and_6_9));
  and_gate and_gate_h_u_dadda_rca16_and_5_10(.a(a[5]), .b(b[10]), .out(h_u_dadda_rca16_and_5_10));
  and_gate and_gate_h_u_dadda_rca16_and_4_11(.a(a[4]), .b(b[11]), .out(h_u_dadda_rca16_and_4_11));
  fa fa_h_u_dadda_rca16_fa66_out(.a(h_u_dadda_rca16_and_6_9[0]), .b(h_u_dadda_rca16_and_5_10[0]), .cin(h_u_dadda_rca16_and_4_11[0]), .fa_xor1(h_u_dadda_rca16_fa66_xor1), .fa_or0(h_u_dadda_rca16_fa66_or0));
  and_gate and_gate_h_u_dadda_rca16_and_3_12(.a(a[3]), .b(b[12]), .out(h_u_dadda_rca16_and_3_12));
  and_gate and_gate_h_u_dadda_rca16_and_2_13(.a(a[2]), .b(b[13]), .out(h_u_dadda_rca16_and_2_13));
  and_gate and_gate_h_u_dadda_rca16_and_1_14(.a(a[1]), .b(b[14]), .out(h_u_dadda_rca16_and_1_14));
  fa fa_h_u_dadda_rca16_fa67_out(.a(h_u_dadda_rca16_and_3_12[0]), .b(h_u_dadda_rca16_and_2_13[0]), .cin(h_u_dadda_rca16_and_1_14[0]), .fa_xor1(h_u_dadda_rca16_fa67_xor1), .fa_or0(h_u_dadda_rca16_fa67_or0));
  and_gate and_gate_h_u_dadda_rca16_and_0_15(.a(a[0]), .b(b[15]), .out(h_u_dadda_rca16_and_0_15));
  fa fa_h_u_dadda_rca16_fa68_out(.a(h_u_dadda_rca16_and_0_15[0]), .b(h_u_dadda_rca16_fa1_xor1[0]), .cin(h_u_dadda_rca16_fa2_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa68_xor1), .fa_or0(h_u_dadda_rca16_fa68_or0));
  fa fa_h_u_dadda_rca16_fa69_out(.a(h_u_dadda_rca16_ha2_xor0[0]), .b(h_u_dadda_rca16_fa62_xor1[0]), .cin(h_u_dadda_rca16_fa63_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa69_xor1), .fa_or0(h_u_dadda_rca16_fa69_or0));
  fa fa_h_u_dadda_rca16_fa70_out(.a(h_u_dadda_rca16_fa64_xor1[0]), .b(h_u_dadda_rca16_fa65_xor1[0]), .cin(h_u_dadda_rca16_fa66_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa70_xor1), .fa_or0(h_u_dadda_rca16_fa70_or0));
  fa fa_h_u_dadda_rca16_fa71_out(.a(h_u_dadda_rca16_fa70_or0[0]), .b(h_u_dadda_rca16_fa69_or0[0]), .cin(h_u_dadda_rca16_fa68_or0[0]), .fa_xor1(h_u_dadda_rca16_fa71_xor1), .fa_or0(h_u_dadda_rca16_fa71_or0));
  fa fa_h_u_dadda_rca16_fa72_out(.a(h_u_dadda_rca16_fa67_or0[0]), .b(h_u_dadda_rca16_fa66_or0[0]), .cin(h_u_dadda_rca16_fa65_or0[0]), .fa_xor1(h_u_dadda_rca16_fa72_xor1), .fa_or0(h_u_dadda_rca16_fa72_or0));
  fa fa_h_u_dadda_rca16_fa73_out(.a(h_u_dadda_rca16_fa64_or0[0]), .b(h_u_dadda_rca16_fa63_or0[0]), .cin(h_u_dadda_rca16_fa62_or0[0]), .fa_xor1(h_u_dadda_rca16_fa73_xor1), .fa_or0(h_u_dadda_rca16_fa73_or0));
  and_gate and_gate_h_u_dadda_rca16_and_10_6(.a(a[10]), .b(b[6]), .out(h_u_dadda_rca16_and_10_6));
  and_gate and_gate_h_u_dadda_rca16_and_9_7(.a(a[9]), .b(b[7]), .out(h_u_dadda_rca16_and_9_7));
  and_gate and_gate_h_u_dadda_rca16_and_8_8(.a(a[8]), .b(b[8]), .out(h_u_dadda_rca16_and_8_8));
  fa fa_h_u_dadda_rca16_fa74_out(.a(h_u_dadda_rca16_and_10_6[0]), .b(h_u_dadda_rca16_and_9_7[0]), .cin(h_u_dadda_rca16_and_8_8[0]), .fa_xor1(h_u_dadda_rca16_fa74_xor1), .fa_or0(h_u_dadda_rca16_fa74_or0));
  and_gate and_gate_h_u_dadda_rca16_and_7_9(.a(a[7]), .b(b[9]), .out(h_u_dadda_rca16_and_7_9));
  and_gate and_gate_h_u_dadda_rca16_and_6_10(.a(a[6]), .b(b[10]), .out(h_u_dadda_rca16_and_6_10));
  and_gate and_gate_h_u_dadda_rca16_and_5_11(.a(a[5]), .b(b[11]), .out(h_u_dadda_rca16_and_5_11));
  fa fa_h_u_dadda_rca16_fa75_out(.a(h_u_dadda_rca16_and_7_9[0]), .b(h_u_dadda_rca16_and_6_10[0]), .cin(h_u_dadda_rca16_and_5_11[0]), .fa_xor1(h_u_dadda_rca16_fa75_xor1), .fa_or0(h_u_dadda_rca16_fa75_or0));
  and_gate and_gate_h_u_dadda_rca16_and_4_12(.a(a[4]), .b(b[12]), .out(h_u_dadda_rca16_and_4_12));
  and_gate and_gate_h_u_dadda_rca16_and_3_13(.a(a[3]), .b(b[13]), .out(h_u_dadda_rca16_and_3_13));
  and_gate and_gate_h_u_dadda_rca16_and_2_14(.a(a[2]), .b(b[14]), .out(h_u_dadda_rca16_and_2_14));
  fa fa_h_u_dadda_rca16_fa76_out(.a(h_u_dadda_rca16_and_4_12[0]), .b(h_u_dadda_rca16_and_3_13[0]), .cin(h_u_dadda_rca16_and_2_14[0]), .fa_xor1(h_u_dadda_rca16_fa76_xor1), .fa_or0(h_u_dadda_rca16_fa76_or0));
  and_gate and_gate_h_u_dadda_rca16_and_1_15(.a(a[1]), .b(b[15]), .out(h_u_dadda_rca16_and_1_15));
  fa fa_h_u_dadda_rca16_fa77_out(.a(h_u_dadda_rca16_and_1_15[0]), .b(h_u_dadda_rca16_fa3_xor1[0]), .cin(h_u_dadda_rca16_fa4_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa77_xor1), .fa_or0(h_u_dadda_rca16_fa77_or0));
  fa fa_h_u_dadda_rca16_fa78_out(.a(h_u_dadda_rca16_ha3_xor0[0]), .b(h_u_dadda_rca16_fa71_xor1[0]), .cin(h_u_dadda_rca16_fa72_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa78_xor1), .fa_or0(h_u_dadda_rca16_fa78_or0));
  fa fa_h_u_dadda_rca16_fa79_out(.a(h_u_dadda_rca16_fa73_xor1[0]), .b(h_u_dadda_rca16_fa74_xor1[0]), .cin(h_u_dadda_rca16_fa75_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa79_xor1), .fa_or0(h_u_dadda_rca16_fa79_or0));
  fa fa_h_u_dadda_rca16_fa80_out(.a(h_u_dadda_rca16_fa79_or0[0]), .b(h_u_dadda_rca16_fa78_or0[0]), .cin(h_u_dadda_rca16_fa77_or0[0]), .fa_xor1(h_u_dadda_rca16_fa80_xor1), .fa_or0(h_u_dadda_rca16_fa80_or0));
  fa fa_h_u_dadda_rca16_fa81_out(.a(h_u_dadda_rca16_fa76_or0[0]), .b(h_u_dadda_rca16_fa75_or0[0]), .cin(h_u_dadda_rca16_fa74_or0[0]), .fa_xor1(h_u_dadda_rca16_fa81_xor1), .fa_or0(h_u_dadda_rca16_fa81_or0));
  fa fa_h_u_dadda_rca16_fa82_out(.a(h_u_dadda_rca16_fa73_or0[0]), .b(h_u_dadda_rca16_fa72_or0[0]), .cin(h_u_dadda_rca16_fa71_or0[0]), .fa_xor1(h_u_dadda_rca16_fa82_xor1), .fa_or0(h_u_dadda_rca16_fa82_or0));
  and_gate and_gate_h_u_dadda_rca16_and_12_5(.a(a[12]), .b(b[5]), .out(h_u_dadda_rca16_and_12_5));
  and_gate and_gate_h_u_dadda_rca16_and_11_6(.a(a[11]), .b(b[6]), .out(h_u_dadda_rca16_and_11_6));
  and_gate and_gate_h_u_dadda_rca16_and_10_7(.a(a[10]), .b(b[7]), .out(h_u_dadda_rca16_and_10_7));
  fa fa_h_u_dadda_rca16_fa83_out(.a(h_u_dadda_rca16_and_12_5[0]), .b(h_u_dadda_rca16_and_11_6[0]), .cin(h_u_dadda_rca16_and_10_7[0]), .fa_xor1(h_u_dadda_rca16_fa83_xor1), .fa_or0(h_u_dadda_rca16_fa83_or0));
  and_gate and_gate_h_u_dadda_rca16_and_9_8(.a(a[9]), .b(b[8]), .out(h_u_dadda_rca16_and_9_8));
  and_gate and_gate_h_u_dadda_rca16_and_8_9(.a(a[8]), .b(b[9]), .out(h_u_dadda_rca16_and_8_9));
  and_gate and_gate_h_u_dadda_rca16_and_7_10(.a(a[7]), .b(b[10]), .out(h_u_dadda_rca16_and_7_10));
  fa fa_h_u_dadda_rca16_fa84_out(.a(h_u_dadda_rca16_and_9_8[0]), .b(h_u_dadda_rca16_and_8_9[0]), .cin(h_u_dadda_rca16_and_7_10[0]), .fa_xor1(h_u_dadda_rca16_fa84_xor1), .fa_or0(h_u_dadda_rca16_fa84_or0));
  and_gate and_gate_h_u_dadda_rca16_and_6_11(.a(a[6]), .b(b[11]), .out(h_u_dadda_rca16_and_6_11));
  and_gate and_gate_h_u_dadda_rca16_and_5_12(.a(a[5]), .b(b[12]), .out(h_u_dadda_rca16_and_5_12));
  and_gate and_gate_h_u_dadda_rca16_and_4_13(.a(a[4]), .b(b[13]), .out(h_u_dadda_rca16_and_4_13));
  fa fa_h_u_dadda_rca16_fa85_out(.a(h_u_dadda_rca16_and_6_11[0]), .b(h_u_dadda_rca16_and_5_12[0]), .cin(h_u_dadda_rca16_and_4_13[0]), .fa_xor1(h_u_dadda_rca16_fa85_xor1), .fa_or0(h_u_dadda_rca16_fa85_or0));
  and_gate and_gate_h_u_dadda_rca16_and_3_14(.a(a[3]), .b(b[14]), .out(h_u_dadda_rca16_and_3_14));
  and_gate and_gate_h_u_dadda_rca16_and_2_15(.a(a[2]), .b(b[15]), .out(h_u_dadda_rca16_and_2_15));
  fa fa_h_u_dadda_rca16_fa86_out(.a(h_u_dadda_rca16_and_3_14[0]), .b(h_u_dadda_rca16_and_2_15[0]), .cin(h_u_dadda_rca16_fa5_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa86_xor1), .fa_or0(h_u_dadda_rca16_fa86_or0));
  fa fa_h_u_dadda_rca16_fa87_out(.a(h_u_dadda_rca16_fa6_xor1[0]), .b(h_u_dadda_rca16_fa80_xor1[0]), .cin(h_u_dadda_rca16_fa81_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa87_xor1), .fa_or0(h_u_dadda_rca16_fa87_or0));
  fa fa_h_u_dadda_rca16_fa88_out(.a(h_u_dadda_rca16_fa82_xor1[0]), .b(h_u_dadda_rca16_fa83_xor1[0]), .cin(h_u_dadda_rca16_fa84_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa88_xor1), .fa_or0(h_u_dadda_rca16_fa88_or0));
  fa fa_h_u_dadda_rca16_fa89_out(.a(h_u_dadda_rca16_fa88_or0[0]), .b(h_u_dadda_rca16_fa87_or0[0]), .cin(h_u_dadda_rca16_fa86_or0[0]), .fa_xor1(h_u_dadda_rca16_fa89_xor1), .fa_or0(h_u_dadda_rca16_fa89_or0));
  fa fa_h_u_dadda_rca16_fa90_out(.a(h_u_dadda_rca16_fa85_or0[0]), .b(h_u_dadda_rca16_fa84_or0[0]), .cin(h_u_dadda_rca16_fa83_or0[0]), .fa_xor1(h_u_dadda_rca16_fa90_xor1), .fa_or0(h_u_dadda_rca16_fa90_or0));
  fa fa_h_u_dadda_rca16_fa91_out(.a(h_u_dadda_rca16_fa82_or0[0]), .b(h_u_dadda_rca16_fa81_or0[0]), .cin(h_u_dadda_rca16_fa80_or0[0]), .fa_xor1(h_u_dadda_rca16_fa91_xor1), .fa_or0(h_u_dadda_rca16_fa91_or0));
  and_gate and_gate_h_u_dadda_rca16_and_14_4(.a(a[14]), .b(b[4]), .out(h_u_dadda_rca16_and_14_4));
  and_gate and_gate_h_u_dadda_rca16_and_13_5(.a(a[13]), .b(b[5]), .out(h_u_dadda_rca16_and_13_5));
  and_gate and_gate_h_u_dadda_rca16_and_12_6(.a(a[12]), .b(b[6]), .out(h_u_dadda_rca16_and_12_6));
  fa fa_h_u_dadda_rca16_fa92_out(.a(h_u_dadda_rca16_and_14_4[0]), .b(h_u_dadda_rca16_and_13_5[0]), .cin(h_u_dadda_rca16_and_12_6[0]), .fa_xor1(h_u_dadda_rca16_fa92_xor1), .fa_or0(h_u_dadda_rca16_fa92_or0));
  and_gate and_gate_h_u_dadda_rca16_and_11_7(.a(a[11]), .b(b[7]), .out(h_u_dadda_rca16_and_11_7));
  and_gate and_gate_h_u_dadda_rca16_and_10_8(.a(a[10]), .b(b[8]), .out(h_u_dadda_rca16_and_10_8));
  and_gate and_gate_h_u_dadda_rca16_and_9_9(.a(a[9]), .b(b[9]), .out(h_u_dadda_rca16_and_9_9));
  fa fa_h_u_dadda_rca16_fa93_out(.a(h_u_dadda_rca16_and_11_7[0]), .b(h_u_dadda_rca16_and_10_8[0]), .cin(h_u_dadda_rca16_and_9_9[0]), .fa_xor1(h_u_dadda_rca16_fa93_xor1), .fa_or0(h_u_dadda_rca16_fa93_or0));
  and_gate and_gate_h_u_dadda_rca16_and_8_10(.a(a[8]), .b(b[10]), .out(h_u_dadda_rca16_and_8_10));
  and_gate and_gate_h_u_dadda_rca16_and_7_11(.a(a[7]), .b(b[11]), .out(h_u_dadda_rca16_and_7_11));
  and_gate and_gate_h_u_dadda_rca16_and_6_12(.a(a[6]), .b(b[12]), .out(h_u_dadda_rca16_and_6_12));
  fa fa_h_u_dadda_rca16_fa94_out(.a(h_u_dadda_rca16_and_8_10[0]), .b(h_u_dadda_rca16_and_7_11[0]), .cin(h_u_dadda_rca16_and_6_12[0]), .fa_xor1(h_u_dadda_rca16_fa94_xor1), .fa_or0(h_u_dadda_rca16_fa94_or0));
  and_gate and_gate_h_u_dadda_rca16_and_5_13(.a(a[5]), .b(b[13]), .out(h_u_dadda_rca16_and_5_13));
  and_gate and_gate_h_u_dadda_rca16_and_4_14(.a(a[4]), .b(b[14]), .out(h_u_dadda_rca16_and_4_14));
  and_gate and_gate_h_u_dadda_rca16_and_3_15(.a(a[3]), .b(b[15]), .out(h_u_dadda_rca16_and_3_15));
  fa fa_h_u_dadda_rca16_fa95_out(.a(h_u_dadda_rca16_and_5_13[0]), .b(h_u_dadda_rca16_and_4_14[0]), .cin(h_u_dadda_rca16_and_3_15[0]), .fa_xor1(h_u_dadda_rca16_fa95_xor1), .fa_or0(h_u_dadda_rca16_fa95_or0));
  fa fa_h_u_dadda_rca16_fa96_out(.a(h_u_dadda_rca16_fa7_xor1[0]), .b(h_u_dadda_rca16_fa89_xor1[0]), .cin(h_u_dadda_rca16_fa90_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa96_xor1), .fa_or0(h_u_dadda_rca16_fa96_or0));
  fa fa_h_u_dadda_rca16_fa97_out(.a(h_u_dadda_rca16_fa91_xor1[0]), .b(h_u_dadda_rca16_fa92_xor1[0]), .cin(h_u_dadda_rca16_fa93_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa97_xor1), .fa_or0(h_u_dadda_rca16_fa97_or0));
  fa fa_h_u_dadda_rca16_fa98_out(.a(h_u_dadda_rca16_fa97_or0[0]), .b(h_u_dadda_rca16_fa96_or0[0]), .cin(h_u_dadda_rca16_fa95_or0[0]), .fa_xor1(h_u_dadda_rca16_fa98_xor1), .fa_or0(h_u_dadda_rca16_fa98_or0));
  fa fa_h_u_dadda_rca16_fa99_out(.a(h_u_dadda_rca16_fa94_or0[0]), .b(h_u_dadda_rca16_fa93_or0[0]), .cin(h_u_dadda_rca16_fa92_or0[0]), .fa_xor1(h_u_dadda_rca16_fa99_xor1), .fa_or0(h_u_dadda_rca16_fa99_or0));
  fa fa_h_u_dadda_rca16_fa100_out(.a(h_u_dadda_rca16_fa91_or0[0]), .b(h_u_dadda_rca16_fa90_or0[0]), .cin(h_u_dadda_rca16_fa89_or0[0]), .fa_xor1(h_u_dadda_rca16_fa100_xor1), .fa_or0(h_u_dadda_rca16_fa100_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_4(.a(a[15]), .b(b[4]), .out(h_u_dadda_rca16_and_15_4));
  and_gate and_gate_h_u_dadda_rca16_and_14_5(.a(a[14]), .b(b[5]), .out(h_u_dadda_rca16_and_14_5));
  fa fa_h_u_dadda_rca16_fa101_out(.a(h_u_dadda_rca16_fa7_or0[0]), .b(h_u_dadda_rca16_and_15_4[0]), .cin(h_u_dadda_rca16_and_14_5[0]), .fa_xor1(h_u_dadda_rca16_fa101_xor1), .fa_or0(h_u_dadda_rca16_fa101_or0));
  and_gate and_gate_h_u_dadda_rca16_and_13_6(.a(a[13]), .b(b[6]), .out(h_u_dadda_rca16_and_13_6));
  and_gate and_gate_h_u_dadda_rca16_and_12_7(.a(a[12]), .b(b[7]), .out(h_u_dadda_rca16_and_12_7));
  and_gate and_gate_h_u_dadda_rca16_and_11_8(.a(a[11]), .b(b[8]), .out(h_u_dadda_rca16_and_11_8));
  fa fa_h_u_dadda_rca16_fa102_out(.a(h_u_dadda_rca16_and_13_6[0]), .b(h_u_dadda_rca16_and_12_7[0]), .cin(h_u_dadda_rca16_and_11_8[0]), .fa_xor1(h_u_dadda_rca16_fa102_xor1), .fa_or0(h_u_dadda_rca16_fa102_or0));
  and_gate and_gate_h_u_dadda_rca16_and_10_9(.a(a[10]), .b(b[9]), .out(h_u_dadda_rca16_and_10_9));
  and_gate and_gate_h_u_dadda_rca16_and_9_10(.a(a[9]), .b(b[10]), .out(h_u_dadda_rca16_and_9_10));
  and_gate and_gate_h_u_dadda_rca16_and_8_11(.a(a[8]), .b(b[11]), .out(h_u_dadda_rca16_and_8_11));
  fa fa_h_u_dadda_rca16_fa103_out(.a(h_u_dadda_rca16_and_10_9[0]), .b(h_u_dadda_rca16_and_9_10[0]), .cin(h_u_dadda_rca16_and_8_11[0]), .fa_xor1(h_u_dadda_rca16_fa103_xor1), .fa_or0(h_u_dadda_rca16_fa103_or0));
  and_gate and_gate_h_u_dadda_rca16_and_7_12(.a(a[7]), .b(b[12]), .out(h_u_dadda_rca16_and_7_12));
  and_gate and_gate_h_u_dadda_rca16_and_6_13(.a(a[6]), .b(b[13]), .out(h_u_dadda_rca16_and_6_13));
  and_gate and_gate_h_u_dadda_rca16_and_5_14(.a(a[5]), .b(b[14]), .out(h_u_dadda_rca16_and_5_14));
  fa fa_h_u_dadda_rca16_fa104_out(.a(h_u_dadda_rca16_and_7_12[0]), .b(h_u_dadda_rca16_and_6_13[0]), .cin(h_u_dadda_rca16_and_5_14[0]), .fa_xor1(h_u_dadda_rca16_fa104_xor1), .fa_or0(h_u_dadda_rca16_fa104_or0));
  and_gate and_gate_h_u_dadda_rca16_and_4_15(.a(a[4]), .b(b[15]), .out(h_u_dadda_rca16_and_4_15));
  fa fa_h_u_dadda_rca16_fa105_out(.a(h_u_dadda_rca16_and_4_15[0]), .b(h_u_dadda_rca16_fa98_xor1[0]), .cin(h_u_dadda_rca16_fa99_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa105_xor1), .fa_or0(h_u_dadda_rca16_fa105_or0));
  fa fa_h_u_dadda_rca16_fa106_out(.a(h_u_dadda_rca16_fa100_xor1[0]), .b(h_u_dadda_rca16_fa101_xor1[0]), .cin(h_u_dadda_rca16_fa102_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa106_xor1), .fa_or0(h_u_dadda_rca16_fa106_or0));
  fa fa_h_u_dadda_rca16_fa107_out(.a(h_u_dadda_rca16_fa106_or0[0]), .b(h_u_dadda_rca16_fa105_or0[0]), .cin(h_u_dadda_rca16_fa104_or0[0]), .fa_xor1(h_u_dadda_rca16_fa107_xor1), .fa_or0(h_u_dadda_rca16_fa107_or0));
  fa fa_h_u_dadda_rca16_fa108_out(.a(h_u_dadda_rca16_fa103_or0[0]), .b(h_u_dadda_rca16_fa102_or0[0]), .cin(h_u_dadda_rca16_fa101_or0[0]), .fa_xor1(h_u_dadda_rca16_fa108_xor1), .fa_or0(h_u_dadda_rca16_fa108_or0));
  fa fa_h_u_dadda_rca16_fa109_out(.a(h_u_dadda_rca16_fa100_or0[0]), .b(h_u_dadda_rca16_fa99_or0[0]), .cin(h_u_dadda_rca16_fa98_or0[0]), .fa_xor1(h_u_dadda_rca16_fa109_xor1), .fa_or0(h_u_dadda_rca16_fa109_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_5(.a(a[15]), .b(b[5]), .out(h_u_dadda_rca16_and_15_5));
  and_gate and_gate_h_u_dadda_rca16_and_14_6(.a(a[14]), .b(b[6]), .out(h_u_dadda_rca16_and_14_6));
  and_gate and_gate_h_u_dadda_rca16_and_13_7(.a(a[13]), .b(b[7]), .out(h_u_dadda_rca16_and_13_7));
  fa fa_h_u_dadda_rca16_fa110_out(.a(h_u_dadda_rca16_and_15_5[0]), .b(h_u_dadda_rca16_and_14_6[0]), .cin(h_u_dadda_rca16_and_13_7[0]), .fa_xor1(h_u_dadda_rca16_fa110_xor1), .fa_or0(h_u_dadda_rca16_fa110_or0));
  and_gate and_gate_h_u_dadda_rca16_and_12_8(.a(a[12]), .b(b[8]), .out(h_u_dadda_rca16_and_12_8));
  and_gate and_gate_h_u_dadda_rca16_and_11_9(.a(a[11]), .b(b[9]), .out(h_u_dadda_rca16_and_11_9));
  and_gate and_gate_h_u_dadda_rca16_and_10_10(.a(a[10]), .b(b[10]), .out(h_u_dadda_rca16_and_10_10));
  fa fa_h_u_dadda_rca16_fa111_out(.a(h_u_dadda_rca16_and_12_8[0]), .b(h_u_dadda_rca16_and_11_9[0]), .cin(h_u_dadda_rca16_and_10_10[0]), .fa_xor1(h_u_dadda_rca16_fa111_xor1), .fa_or0(h_u_dadda_rca16_fa111_or0));
  and_gate and_gate_h_u_dadda_rca16_and_9_11(.a(a[9]), .b(b[11]), .out(h_u_dadda_rca16_and_9_11));
  and_gate and_gate_h_u_dadda_rca16_and_8_12(.a(a[8]), .b(b[12]), .out(h_u_dadda_rca16_and_8_12));
  and_gate and_gate_h_u_dadda_rca16_and_7_13(.a(a[7]), .b(b[13]), .out(h_u_dadda_rca16_and_7_13));
  fa fa_h_u_dadda_rca16_fa112_out(.a(h_u_dadda_rca16_and_9_11[0]), .b(h_u_dadda_rca16_and_8_12[0]), .cin(h_u_dadda_rca16_and_7_13[0]), .fa_xor1(h_u_dadda_rca16_fa112_xor1), .fa_or0(h_u_dadda_rca16_fa112_or0));
  and_gate and_gate_h_u_dadda_rca16_and_6_14(.a(a[6]), .b(b[14]), .out(h_u_dadda_rca16_and_6_14));
  and_gate and_gate_h_u_dadda_rca16_and_5_15(.a(a[5]), .b(b[15]), .out(h_u_dadda_rca16_and_5_15));
  fa fa_h_u_dadda_rca16_fa113_out(.a(h_u_dadda_rca16_and_6_14[0]), .b(h_u_dadda_rca16_and_5_15[0]), .cin(h_u_dadda_rca16_fa107_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa113_xor1), .fa_or0(h_u_dadda_rca16_fa113_or0));
  fa fa_h_u_dadda_rca16_fa114_out(.a(h_u_dadda_rca16_fa108_xor1[0]), .b(h_u_dadda_rca16_fa109_xor1[0]), .cin(h_u_dadda_rca16_fa110_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa114_xor1), .fa_or0(h_u_dadda_rca16_fa114_or0));
  fa fa_h_u_dadda_rca16_fa115_out(.a(h_u_dadda_rca16_fa114_or0[0]), .b(h_u_dadda_rca16_fa113_or0[0]), .cin(h_u_dadda_rca16_fa112_or0[0]), .fa_xor1(h_u_dadda_rca16_fa115_xor1), .fa_or0(h_u_dadda_rca16_fa115_or0));
  fa fa_h_u_dadda_rca16_fa116_out(.a(h_u_dadda_rca16_fa111_or0[0]), .b(h_u_dadda_rca16_fa110_or0[0]), .cin(h_u_dadda_rca16_fa109_or0[0]), .fa_xor1(h_u_dadda_rca16_fa116_xor1), .fa_or0(h_u_dadda_rca16_fa116_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_6(.a(a[15]), .b(b[6]), .out(h_u_dadda_rca16_and_15_6));
  fa fa_h_u_dadda_rca16_fa117_out(.a(h_u_dadda_rca16_fa108_or0[0]), .b(h_u_dadda_rca16_fa107_or0[0]), .cin(h_u_dadda_rca16_and_15_6[0]), .fa_xor1(h_u_dadda_rca16_fa117_xor1), .fa_or0(h_u_dadda_rca16_fa117_or0));
  and_gate and_gate_h_u_dadda_rca16_and_14_7(.a(a[14]), .b(b[7]), .out(h_u_dadda_rca16_and_14_7));
  and_gate and_gate_h_u_dadda_rca16_and_13_8(.a(a[13]), .b(b[8]), .out(h_u_dadda_rca16_and_13_8));
  and_gate and_gate_h_u_dadda_rca16_and_12_9(.a(a[12]), .b(b[9]), .out(h_u_dadda_rca16_and_12_9));
  fa fa_h_u_dadda_rca16_fa118_out(.a(h_u_dadda_rca16_and_14_7[0]), .b(h_u_dadda_rca16_and_13_8[0]), .cin(h_u_dadda_rca16_and_12_9[0]), .fa_xor1(h_u_dadda_rca16_fa118_xor1), .fa_or0(h_u_dadda_rca16_fa118_or0));
  and_gate and_gate_h_u_dadda_rca16_and_11_10(.a(a[11]), .b(b[10]), .out(h_u_dadda_rca16_and_11_10));
  and_gate and_gate_h_u_dadda_rca16_and_10_11(.a(a[10]), .b(b[11]), .out(h_u_dadda_rca16_and_10_11));
  and_gate and_gate_h_u_dadda_rca16_and_9_12(.a(a[9]), .b(b[12]), .out(h_u_dadda_rca16_and_9_12));
  fa fa_h_u_dadda_rca16_fa119_out(.a(h_u_dadda_rca16_and_11_10[0]), .b(h_u_dadda_rca16_and_10_11[0]), .cin(h_u_dadda_rca16_and_9_12[0]), .fa_xor1(h_u_dadda_rca16_fa119_xor1), .fa_or0(h_u_dadda_rca16_fa119_or0));
  and_gate and_gate_h_u_dadda_rca16_and_8_13(.a(a[8]), .b(b[13]), .out(h_u_dadda_rca16_and_8_13));
  and_gate and_gate_h_u_dadda_rca16_and_7_14(.a(a[7]), .b(b[14]), .out(h_u_dadda_rca16_and_7_14));
  and_gate and_gate_h_u_dadda_rca16_and_6_15(.a(a[6]), .b(b[15]), .out(h_u_dadda_rca16_and_6_15));
  fa fa_h_u_dadda_rca16_fa120_out(.a(h_u_dadda_rca16_and_8_13[0]), .b(h_u_dadda_rca16_and_7_14[0]), .cin(h_u_dadda_rca16_and_6_15[0]), .fa_xor1(h_u_dadda_rca16_fa120_xor1), .fa_or0(h_u_dadda_rca16_fa120_or0));
  fa fa_h_u_dadda_rca16_fa121_out(.a(h_u_dadda_rca16_fa115_xor1[0]), .b(h_u_dadda_rca16_fa116_xor1[0]), .cin(h_u_dadda_rca16_fa117_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa121_xor1), .fa_or0(h_u_dadda_rca16_fa121_or0));
  fa fa_h_u_dadda_rca16_fa122_out(.a(h_u_dadda_rca16_fa121_or0[0]), .b(h_u_dadda_rca16_fa120_or0[0]), .cin(h_u_dadda_rca16_fa119_or0[0]), .fa_xor1(h_u_dadda_rca16_fa122_xor1), .fa_or0(h_u_dadda_rca16_fa122_or0));
  fa fa_h_u_dadda_rca16_fa123_out(.a(h_u_dadda_rca16_fa118_or0[0]), .b(h_u_dadda_rca16_fa117_or0[0]), .cin(h_u_dadda_rca16_fa116_or0[0]), .fa_xor1(h_u_dadda_rca16_fa123_xor1), .fa_or0(h_u_dadda_rca16_fa123_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_7(.a(a[15]), .b(b[7]), .out(h_u_dadda_rca16_and_15_7));
  and_gate and_gate_h_u_dadda_rca16_and_14_8(.a(a[14]), .b(b[8]), .out(h_u_dadda_rca16_and_14_8));
  fa fa_h_u_dadda_rca16_fa124_out(.a(h_u_dadda_rca16_fa115_or0[0]), .b(h_u_dadda_rca16_and_15_7[0]), .cin(h_u_dadda_rca16_and_14_8[0]), .fa_xor1(h_u_dadda_rca16_fa124_xor1), .fa_or0(h_u_dadda_rca16_fa124_or0));
  and_gate and_gate_h_u_dadda_rca16_and_13_9(.a(a[13]), .b(b[9]), .out(h_u_dadda_rca16_and_13_9));
  and_gate and_gate_h_u_dadda_rca16_and_12_10(.a(a[12]), .b(b[10]), .out(h_u_dadda_rca16_and_12_10));
  and_gate and_gate_h_u_dadda_rca16_and_11_11(.a(a[11]), .b(b[11]), .out(h_u_dadda_rca16_and_11_11));
  fa fa_h_u_dadda_rca16_fa125_out(.a(h_u_dadda_rca16_and_13_9[0]), .b(h_u_dadda_rca16_and_12_10[0]), .cin(h_u_dadda_rca16_and_11_11[0]), .fa_xor1(h_u_dadda_rca16_fa125_xor1), .fa_or0(h_u_dadda_rca16_fa125_or0));
  and_gate and_gate_h_u_dadda_rca16_and_10_12(.a(a[10]), .b(b[12]), .out(h_u_dadda_rca16_and_10_12));
  and_gate and_gate_h_u_dadda_rca16_and_9_13(.a(a[9]), .b(b[13]), .out(h_u_dadda_rca16_and_9_13));
  and_gate and_gate_h_u_dadda_rca16_and_8_14(.a(a[8]), .b(b[14]), .out(h_u_dadda_rca16_and_8_14));
  fa fa_h_u_dadda_rca16_fa126_out(.a(h_u_dadda_rca16_and_10_12[0]), .b(h_u_dadda_rca16_and_9_13[0]), .cin(h_u_dadda_rca16_and_8_14[0]), .fa_xor1(h_u_dadda_rca16_fa126_xor1), .fa_or0(h_u_dadda_rca16_fa126_or0));
  and_gate and_gate_h_u_dadda_rca16_and_7_15(.a(a[7]), .b(b[15]), .out(h_u_dadda_rca16_and_7_15));
  fa fa_h_u_dadda_rca16_fa127_out(.a(h_u_dadda_rca16_and_7_15[0]), .b(h_u_dadda_rca16_fa122_xor1[0]), .cin(h_u_dadda_rca16_fa123_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa127_xor1), .fa_or0(h_u_dadda_rca16_fa127_or0));
  fa fa_h_u_dadda_rca16_fa128_out(.a(h_u_dadda_rca16_fa127_or0[0]), .b(h_u_dadda_rca16_fa126_or0[0]), .cin(h_u_dadda_rca16_fa125_or0[0]), .fa_xor1(h_u_dadda_rca16_fa128_xor1), .fa_or0(h_u_dadda_rca16_fa128_or0));
  fa fa_h_u_dadda_rca16_fa129_out(.a(h_u_dadda_rca16_fa124_or0[0]), .b(h_u_dadda_rca16_fa123_or0[0]), .cin(h_u_dadda_rca16_fa122_or0[0]), .fa_xor1(h_u_dadda_rca16_fa129_xor1), .fa_or0(h_u_dadda_rca16_fa129_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_8(.a(a[15]), .b(b[8]), .out(h_u_dadda_rca16_and_15_8));
  and_gate and_gate_h_u_dadda_rca16_and_14_9(.a(a[14]), .b(b[9]), .out(h_u_dadda_rca16_and_14_9));
  and_gate and_gate_h_u_dadda_rca16_and_13_10(.a(a[13]), .b(b[10]), .out(h_u_dadda_rca16_and_13_10));
  fa fa_h_u_dadda_rca16_fa130_out(.a(h_u_dadda_rca16_and_15_8[0]), .b(h_u_dadda_rca16_and_14_9[0]), .cin(h_u_dadda_rca16_and_13_10[0]), .fa_xor1(h_u_dadda_rca16_fa130_xor1), .fa_or0(h_u_dadda_rca16_fa130_or0));
  and_gate and_gate_h_u_dadda_rca16_and_12_11(.a(a[12]), .b(b[11]), .out(h_u_dadda_rca16_and_12_11));
  and_gate and_gate_h_u_dadda_rca16_and_11_12(.a(a[11]), .b(b[12]), .out(h_u_dadda_rca16_and_11_12));
  and_gate and_gate_h_u_dadda_rca16_and_10_13(.a(a[10]), .b(b[13]), .out(h_u_dadda_rca16_and_10_13));
  fa fa_h_u_dadda_rca16_fa131_out(.a(h_u_dadda_rca16_and_12_11[0]), .b(h_u_dadda_rca16_and_11_12[0]), .cin(h_u_dadda_rca16_and_10_13[0]), .fa_xor1(h_u_dadda_rca16_fa131_xor1), .fa_or0(h_u_dadda_rca16_fa131_or0));
  and_gate and_gate_h_u_dadda_rca16_and_9_14(.a(a[9]), .b(b[14]), .out(h_u_dadda_rca16_and_9_14));
  and_gate and_gate_h_u_dadda_rca16_and_8_15(.a(a[8]), .b(b[15]), .out(h_u_dadda_rca16_and_8_15));
  fa fa_h_u_dadda_rca16_fa132_out(.a(h_u_dadda_rca16_and_9_14[0]), .b(h_u_dadda_rca16_and_8_15[0]), .cin(h_u_dadda_rca16_fa128_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa132_xor1), .fa_or0(h_u_dadda_rca16_fa132_or0));
  fa fa_h_u_dadda_rca16_fa133_out(.a(h_u_dadda_rca16_fa132_or0[0]), .b(h_u_dadda_rca16_fa131_or0[0]), .cin(h_u_dadda_rca16_fa130_or0[0]), .fa_xor1(h_u_dadda_rca16_fa133_xor1), .fa_or0(h_u_dadda_rca16_fa133_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_9(.a(a[15]), .b(b[9]), .out(h_u_dadda_rca16_and_15_9));
  fa fa_h_u_dadda_rca16_fa134_out(.a(h_u_dadda_rca16_fa129_or0[0]), .b(h_u_dadda_rca16_fa128_or0[0]), .cin(h_u_dadda_rca16_and_15_9[0]), .fa_xor1(h_u_dadda_rca16_fa134_xor1), .fa_or0(h_u_dadda_rca16_fa134_or0));
  and_gate and_gate_h_u_dadda_rca16_and_14_10(.a(a[14]), .b(b[10]), .out(h_u_dadda_rca16_and_14_10));
  and_gate and_gate_h_u_dadda_rca16_and_13_11(.a(a[13]), .b(b[11]), .out(h_u_dadda_rca16_and_13_11));
  and_gate and_gate_h_u_dadda_rca16_and_12_12(.a(a[12]), .b(b[12]), .out(h_u_dadda_rca16_and_12_12));
  fa fa_h_u_dadda_rca16_fa135_out(.a(h_u_dadda_rca16_and_14_10[0]), .b(h_u_dadda_rca16_and_13_11[0]), .cin(h_u_dadda_rca16_and_12_12[0]), .fa_xor1(h_u_dadda_rca16_fa135_xor1), .fa_or0(h_u_dadda_rca16_fa135_or0));
  and_gate and_gate_h_u_dadda_rca16_and_11_13(.a(a[11]), .b(b[13]), .out(h_u_dadda_rca16_and_11_13));
  and_gate and_gate_h_u_dadda_rca16_and_10_14(.a(a[10]), .b(b[14]), .out(h_u_dadda_rca16_and_10_14));
  and_gate and_gate_h_u_dadda_rca16_and_9_15(.a(a[9]), .b(b[15]), .out(h_u_dadda_rca16_and_9_15));
  fa fa_h_u_dadda_rca16_fa136_out(.a(h_u_dadda_rca16_and_11_13[0]), .b(h_u_dadda_rca16_and_10_14[0]), .cin(h_u_dadda_rca16_and_9_15[0]), .fa_xor1(h_u_dadda_rca16_fa136_xor1), .fa_or0(h_u_dadda_rca16_fa136_or0));
  fa fa_h_u_dadda_rca16_fa137_out(.a(h_u_dadda_rca16_fa136_or0[0]), .b(h_u_dadda_rca16_fa135_or0[0]), .cin(h_u_dadda_rca16_fa134_or0[0]), .fa_xor1(h_u_dadda_rca16_fa137_xor1), .fa_or0(h_u_dadda_rca16_fa137_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_10(.a(a[15]), .b(b[10]), .out(h_u_dadda_rca16_and_15_10));
  and_gate and_gate_h_u_dadda_rca16_and_14_11(.a(a[14]), .b(b[11]), .out(h_u_dadda_rca16_and_14_11));
  fa fa_h_u_dadda_rca16_fa138_out(.a(h_u_dadda_rca16_fa133_or0[0]), .b(h_u_dadda_rca16_and_15_10[0]), .cin(h_u_dadda_rca16_and_14_11[0]), .fa_xor1(h_u_dadda_rca16_fa138_xor1), .fa_or0(h_u_dadda_rca16_fa138_or0));
  and_gate and_gate_h_u_dadda_rca16_and_13_12(.a(a[13]), .b(b[12]), .out(h_u_dadda_rca16_and_13_12));
  and_gate and_gate_h_u_dadda_rca16_and_12_13(.a(a[12]), .b(b[13]), .out(h_u_dadda_rca16_and_12_13));
  and_gate and_gate_h_u_dadda_rca16_and_11_14(.a(a[11]), .b(b[14]), .out(h_u_dadda_rca16_and_11_14));
  fa fa_h_u_dadda_rca16_fa139_out(.a(h_u_dadda_rca16_and_13_12[0]), .b(h_u_dadda_rca16_and_12_13[0]), .cin(h_u_dadda_rca16_and_11_14[0]), .fa_xor1(h_u_dadda_rca16_fa139_xor1), .fa_or0(h_u_dadda_rca16_fa139_or0));
  fa fa_h_u_dadda_rca16_fa140_out(.a(h_u_dadda_rca16_fa139_or0[0]), .b(h_u_dadda_rca16_fa138_or0[0]), .cin(h_u_dadda_rca16_fa137_or0[0]), .fa_xor1(h_u_dadda_rca16_fa140_xor1), .fa_or0(h_u_dadda_rca16_fa140_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_11(.a(a[15]), .b(b[11]), .out(h_u_dadda_rca16_and_15_11));
  and_gate and_gate_h_u_dadda_rca16_and_14_12(.a(a[14]), .b(b[12]), .out(h_u_dadda_rca16_and_14_12));
  and_gate and_gate_h_u_dadda_rca16_and_13_13(.a(a[13]), .b(b[13]), .out(h_u_dadda_rca16_and_13_13));
  fa fa_h_u_dadda_rca16_fa141_out(.a(h_u_dadda_rca16_and_15_11[0]), .b(h_u_dadda_rca16_and_14_12[0]), .cin(h_u_dadda_rca16_and_13_13[0]), .fa_xor1(h_u_dadda_rca16_fa141_xor1), .fa_or0(h_u_dadda_rca16_fa141_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_12(.a(a[15]), .b(b[12]), .out(h_u_dadda_rca16_and_15_12));
  fa fa_h_u_dadda_rca16_fa142_out(.a(h_u_dadda_rca16_fa141_or0[0]), .b(h_u_dadda_rca16_fa140_or0[0]), .cin(h_u_dadda_rca16_and_15_12[0]), .fa_xor1(h_u_dadda_rca16_fa142_xor1), .fa_or0(h_u_dadda_rca16_fa142_or0));
  and_gate and_gate_h_u_dadda_rca16_and_3_0(.a(a[3]), .b(b[0]), .out(h_u_dadda_rca16_and_3_0));
  and_gate and_gate_h_u_dadda_rca16_and_2_1(.a(a[2]), .b(b[1]), .out(h_u_dadda_rca16_and_2_1));
  ha ha_h_u_dadda_rca16_ha13_out(.a(h_u_dadda_rca16_and_3_0[0]), .b(h_u_dadda_rca16_and_2_1[0]), .ha_xor0(h_u_dadda_rca16_ha13_xor0), .ha_and0(h_u_dadda_rca16_ha13_and0));
  and_gate and_gate_h_u_dadda_rca16_and_2_2(.a(a[2]), .b(b[2]), .out(h_u_dadda_rca16_and_2_2));
  and_gate and_gate_h_u_dadda_rca16_and_1_3(.a(a[1]), .b(b[3]), .out(h_u_dadda_rca16_and_1_3));
  fa fa_h_u_dadda_rca16_fa143_out(.a(h_u_dadda_rca16_ha13_and0[0]), .b(h_u_dadda_rca16_and_2_2[0]), .cin(h_u_dadda_rca16_and_1_3[0]), .fa_xor1(h_u_dadda_rca16_fa143_xor1), .fa_or0(h_u_dadda_rca16_fa143_or0));
  and_gate and_gate_h_u_dadda_rca16_and_1_4(.a(a[1]), .b(b[4]), .out(h_u_dadda_rca16_and_1_4));
  and_gate and_gate_h_u_dadda_rca16_and_0_5(.a(a[0]), .b(b[5]), .out(h_u_dadda_rca16_and_0_5));
  fa fa_h_u_dadda_rca16_fa144_out(.a(h_u_dadda_rca16_fa143_or0[0]), .b(h_u_dadda_rca16_and_1_4[0]), .cin(h_u_dadda_rca16_and_0_5[0]), .fa_xor1(h_u_dadda_rca16_fa144_xor1), .fa_or0(h_u_dadda_rca16_fa144_or0));
  and_gate and_gate_h_u_dadda_rca16_and_0_6(.a(a[0]), .b(b[6]), .out(h_u_dadda_rca16_and_0_6));
  fa fa_h_u_dadda_rca16_fa145_out(.a(h_u_dadda_rca16_fa144_or0[0]), .b(h_u_dadda_rca16_and_0_6[0]), .cin(h_u_dadda_rca16_fa9_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa145_xor1), .fa_or0(h_u_dadda_rca16_fa145_or0));
  fa fa_h_u_dadda_rca16_fa146_out(.a(h_u_dadda_rca16_fa145_or0[0]), .b(h_u_dadda_rca16_fa11_xor1[0]), .cin(h_u_dadda_rca16_fa12_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa146_xor1), .fa_or0(h_u_dadda_rca16_fa146_or0));
  fa fa_h_u_dadda_rca16_fa147_out(.a(h_u_dadda_rca16_fa146_or0[0]), .b(h_u_dadda_rca16_fa15_xor1[0]), .cin(h_u_dadda_rca16_fa16_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa147_xor1), .fa_or0(h_u_dadda_rca16_fa147_or0));
  fa fa_h_u_dadda_rca16_fa148_out(.a(h_u_dadda_rca16_fa147_or0[0]), .b(h_u_dadda_rca16_fa20_xor1[0]), .cin(h_u_dadda_rca16_fa21_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa148_xor1), .fa_or0(h_u_dadda_rca16_fa148_or0));
  fa fa_h_u_dadda_rca16_fa149_out(.a(h_u_dadda_rca16_fa148_or0[0]), .b(h_u_dadda_rca16_fa26_xor1[0]), .cin(h_u_dadda_rca16_fa27_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa149_xor1), .fa_or0(h_u_dadda_rca16_fa149_or0));
  fa fa_h_u_dadda_rca16_fa150_out(.a(h_u_dadda_rca16_fa149_or0[0]), .b(h_u_dadda_rca16_fa33_xor1[0]), .cin(h_u_dadda_rca16_fa34_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa150_xor1), .fa_or0(h_u_dadda_rca16_fa150_or0));
  fa fa_h_u_dadda_rca16_fa151_out(.a(h_u_dadda_rca16_fa150_or0[0]), .b(h_u_dadda_rca16_fa41_xor1[0]), .cin(h_u_dadda_rca16_fa42_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa151_xor1), .fa_or0(h_u_dadda_rca16_fa151_or0));
  fa fa_h_u_dadda_rca16_fa152_out(.a(h_u_dadda_rca16_fa151_or0[0]), .b(h_u_dadda_rca16_fa49_xor1[0]), .cin(h_u_dadda_rca16_fa50_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa152_xor1), .fa_or0(h_u_dadda_rca16_fa152_or0));
  fa fa_h_u_dadda_rca16_fa153_out(.a(h_u_dadda_rca16_fa152_or0[0]), .b(h_u_dadda_rca16_fa58_xor1[0]), .cin(h_u_dadda_rca16_fa59_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa153_xor1), .fa_or0(h_u_dadda_rca16_fa153_or0));
  fa fa_h_u_dadda_rca16_fa154_out(.a(h_u_dadda_rca16_fa153_or0[0]), .b(h_u_dadda_rca16_fa67_xor1[0]), .cin(h_u_dadda_rca16_fa68_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa154_xor1), .fa_or0(h_u_dadda_rca16_fa154_or0));
  fa fa_h_u_dadda_rca16_fa155_out(.a(h_u_dadda_rca16_fa154_or0[0]), .b(h_u_dadda_rca16_fa76_xor1[0]), .cin(h_u_dadda_rca16_fa77_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa155_xor1), .fa_or0(h_u_dadda_rca16_fa155_or0));
  fa fa_h_u_dadda_rca16_fa156_out(.a(h_u_dadda_rca16_fa155_or0[0]), .b(h_u_dadda_rca16_fa85_xor1[0]), .cin(h_u_dadda_rca16_fa86_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa156_xor1), .fa_or0(h_u_dadda_rca16_fa156_or0));
  fa fa_h_u_dadda_rca16_fa157_out(.a(h_u_dadda_rca16_fa156_or0[0]), .b(h_u_dadda_rca16_fa94_xor1[0]), .cin(h_u_dadda_rca16_fa95_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa157_xor1), .fa_or0(h_u_dadda_rca16_fa157_or0));
  fa fa_h_u_dadda_rca16_fa158_out(.a(h_u_dadda_rca16_fa157_or0[0]), .b(h_u_dadda_rca16_fa103_xor1[0]), .cin(h_u_dadda_rca16_fa104_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa158_xor1), .fa_or0(h_u_dadda_rca16_fa158_or0));
  fa fa_h_u_dadda_rca16_fa159_out(.a(h_u_dadda_rca16_fa158_or0[0]), .b(h_u_dadda_rca16_fa111_xor1[0]), .cin(h_u_dadda_rca16_fa112_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa159_xor1), .fa_or0(h_u_dadda_rca16_fa159_or0));
  fa fa_h_u_dadda_rca16_fa160_out(.a(h_u_dadda_rca16_fa159_or0[0]), .b(h_u_dadda_rca16_fa118_xor1[0]), .cin(h_u_dadda_rca16_fa119_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa160_xor1), .fa_or0(h_u_dadda_rca16_fa160_or0));
  fa fa_h_u_dadda_rca16_fa161_out(.a(h_u_dadda_rca16_fa160_or0[0]), .b(h_u_dadda_rca16_fa124_xor1[0]), .cin(h_u_dadda_rca16_fa125_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa161_xor1), .fa_or0(h_u_dadda_rca16_fa161_or0));
  fa fa_h_u_dadda_rca16_fa162_out(.a(h_u_dadda_rca16_fa161_or0[0]), .b(h_u_dadda_rca16_fa129_xor1[0]), .cin(h_u_dadda_rca16_fa130_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa162_xor1), .fa_or0(h_u_dadda_rca16_fa162_or0));
  fa fa_h_u_dadda_rca16_fa163_out(.a(h_u_dadda_rca16_fa162_or0[0]), .b(h_u_dadda_rca16_fa133_xor1[0]), .cin(h_u_dadda_rca16_fa134_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa163_xor1), .fa_or0(h_u_dadda_rca16_fa163_or0));
  and_gate and_gate_h_u_dadda_rca16_and_10_15(.a(a[10]), .b(b[15]), .out(h_u_dadda_rca16_and_10_15));
  fa fa_h_u_dadda_rca16_fa164_out(.a(h_u_dadda_rca16_fa163_or0[0]), .b(h_u_dadda_rca16_and_10_15[0]), .cin(h_u_dadda_rca16_fa137_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa164_xor1), .fa_or0(h_u_dadda_rca16_fa164_or0));
  and_gate and_gate_h_u_dadda_rca16_and_12_14(.a(a[12]), .b(b[14]), .out(h_u_dadda_rca16_and_12_14));
  and_gate and_gate_h_u_dadda_rca16_and_11_15(.a(a[11]), .b(b[15]), .out(h_u_dadda_rca16_and_11_15));
  fa fa_h_u_dadda_rca16_fa165_out(.a(h_u_dadda_rca16_fa164_or0[0]), .b(h_u_dadda_rca16_and_12_14[0]), .cin(h_u_dadda_rca16_and_11_15[0]), .fa_xor1(h_u_dadda_rca16_fa165_xor1), .fa_or0(h_u_dadda_rca16_fa165_or0));
  and_gate and_gate_h_u_dadda_rca16_and_14_13(.a(a[14]), .b(b[13]), .out(h_u_dadda_rca16_and_14_13));
  and_gate and_gate_h_u_dadda_rca16_and_13_14(.a(a[13]), .b(b[14]), .out(h_u_dadda_rca16_and_13_14));
  fa fa_h_u_dadda_rca16_fa166_out(.a(h_u_dadda_rca16_fa165_or0[0]), .b(h_u_dadda_rca16_and_14_13[0]), .cin(h_u_dadda_rca16_and_13_14[0]), .fa_xor1(h_u_dadda_rca16_fa166_xor1), .fa_or0(h_u_dadda_rca16_fa166_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_13(.a(a[15]), .b(b[13]), .out(h_u_dadda_rca16_and_15_13));
  fa fa_h_u_dadda_rca16_fa167_out(.a(h_u_dadda_rca16_fa166_or0[0]), .b(h_u_dadda_rca16_fa142_or0[0]), .cin(h_u_dadda_rca16_and_15_13[0]), .fa_xor1(h_u_dadda_rca16_fa167_xor1), .fa_or0(h_u_dadda_rca16_fa167_or0));
  and_gate and_gate_h_u_dadda_rca16_and_2_0(.a(a[2]), .b(b[0]), .out(h_u_dadda_rca16_and_2_0));
  and_gate and_gate_h_u_dadda_rca16_and_1_1(.a(a[1]), .b(b[1]), .out(h_u_dadda_rca16_and_1_1));
  ha ha_h_u_dadda_rca16_ha14_out(.a(h_u_dadda_rca16_and_2_0[0]), .b(h_u_dadda_rca16_and_1_1[0]), .ha_xor0(h_u_dadda_rca16_ha14_xor0), .ha_and0(h_u_dadda_rca16_ha14_and0));
  and_gate and_gate_h_u_dadda_rca16_and_1_2(.a(a[1]), .b(b[2]), .out(h_u_dadda_rca16_and_1_2));
  and_gate and_gate_h_u_dadda_rca16_and_0_3(.a(a[0]), .b(b[3]), .out(h_u_dadda_rca16_and_0_3));
  fa fa_h_u_dadda_rca16_fa168_out(.a(h_u_dadda_rca16_ha14_and0[0]), .b(h_u_dadda_rca16_and_1_2[0]), .cin(h_u_dadda_rca16_and_0_3[0]), .fa_xor1(h_u_dadda_rca16_fa168_xor1), .fa_or0(h_u_dadda_rca16_fa168_or0));
  and_gate and_gate_h_u_dadda_rca16_and_0_4(.a(a[0]), .b(b[4]), .out(h_u_dadda_rca16_and_0_4));
  fa fa_h_u_dadda_rca16_fa169_out(.a(h_u_dadda_rca16_fa168_or0[0]), .b(h_u_dadda_rca16_and_0_4[0]), .cin(h_u_dadda_rca16_ha4_xor0[0]), .fa_xor1(h_u_dadda_rca16_fa169_xor1), .fa_or0(h_u_dadda_rca16_fa169_or0));
  fa fa_h_u_dadda_rca16_fa170_out(.a(h_u_dadda_rca16_fa169_or0[0]), .b(h_u_dadda_rca16_fa8_xor1[0]), .cin(h_u_dadda_rca16_ha5_xor0[0]), .fa_xor1(h_u_dadda_rca16_fa170_xor1), .fa_or0(h_u_dadda_rca16_fa170_or0));
  fa fa_h_u_dadda_rca16_fa171_out(.a(h_u_dadda_rca16_fa170_or0[0]), .b(h_u_dadda_rca16_fa10_xor1[0]), .cin(h_u_dadda_rca16_ha6_xor0[0]), .fa_xor1(h_u_dadda_rca16_fa171_xor1), .fa_or0(h_u_dadda_rca16_fa171_or0));
  fa fa_h_u_dadda_rca16_fa172_out(.a(h_u_dadda_rca16_fa171_or0[0]), .b(h_u_dadda_rca16_fa13_xor1[0]), .cin(h_u_dadda_rca16_ha7_xor0[0]), .fa_xor1(h_u_dadda_rca16_fa172_xor1), .fa_or0(h_u_dadda_rca16_fa172_or0));
  fa fa_h_u_dadda_rca16_fa173_out(.a(h_u_dadda_rca16_fa172_or0[0]), .b(h_u_dadda_rca16_fa17_xor1[0]), .cin(h_u_dadda_rca16_ha8_xor0[0]), .fa_xor1(h_u_dadda_rca16_fa173_xor1), .fa_or0(h_u_dadda_rca16_fa173_or0));
  fa fa_h_u_dadda_rca16_fa174_out(.a(h_u_dadda_rca16_fa173_or0[0]), .b(h_u_dadda_rca16_fa22_xor1[0]), .cin(h_u_dadda_rca16_ha9_xor0[0]), .fa_xor1(h_u_dadda_rca16_fa174_xor1), .fa_or0(h_u_dadda_rca16_fa174_or0));
  fa fa_h_u_dadda_rca16_fa175_out(.a(h_u_dadda_rca16_fa174_or0[0]), .b(h_u_dadda_rca16_fa28_xor1[0]), .cin(h_u_dadda_rca16_ha10_xor0[0]), .fa_xor1(h_u_dadda_rca16_fa175_xor1), .fa_or0(h_u_dadda_rca16_fa175_or0));
  fa fa_h_u_dadda_rca16_fa176_out(.a(h_u_dadda_rca16_fa175_or0[0]), .b(h_u_dadda_rca16_fa35_xor1[0]), .cin(h_u_dadda_rca16_ha11_xor0[0]), .fa_xor1(h_u_dadda_rca16_fa176_xor1), .fa_or0(h_u_dadda_rca16_fa176_or0));
  fa fa_h_u_dadda_rca16_fa177_out(.a(h_u_dadda_rca16_fa176_or0[0]), .b(h_u_dadda_rca16_fa43_xor1[0]), .cin(h_u_dadda_rca16_ha12_xor0[0]), .fa_xor1(h_u_dadda_rca16_fa177_xor1), .fa_or0(h_u_dadda_rca16_fa177_or0));
  fa fa_h_u_dadda_rca16_fa178_out(.a(h_u_dadda_rca16_fa177_or0[0]), .b(h_u_dadda_rca16_fa51_xor1[0]), .cin(h_u_dadda_rca16_fa52_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa178_xor1), .fa_or0(h_u_dadda_rca16_fa178_or0));
  fa fa_h_u_dadda_rca16_fa179_out(.a(h_u_dadda_rca16_fa178_or0[0]), .b(h_u_dadda_rca16_fa60_xor1[0]), .cin(h_u_dadda_rca16_fa61_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa179_xor1), .fa_or0(h_u_dadda_rca16_fa179_or0));
  fa fa_h_u_dadda_rca16_fa180_out(.a(h_u_dadda_rca16_fa179_or0[0]), .b(h_u_dadda_rca16_fa69_xor1[0]), .cin(h_u_dadda_rca16_fa70_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa180_xor1), .fa_or0(h_u_dadda_rca16_fa180_or0));
  fa fa_h_u_dadda_rca16_fa181_out(.a(h_u_dadda_rca16_fa180_or0[0]), .b(h_u_dadda_rca16_fa78_xor1[0]), .cin(h_u_dadda_rca16_fa79_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa181_xor1), .fa_or0(h_u_dadda_rca16_fa181_or0));
  fa fa_h_u_dadda_rca16_fa182_out(.a(h_u_dadda_rca16_fa181_or0[0]), .b(h_u_dadda_rca16_fa87_xor1[0]), .cin(h_u_dadda_rca16_fa88_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa182_xor1), .fa_or0(h_u_dadda_rca16_fa182_or0));
  fa fa_h_u_dadda_rca16_fa183_out(.a(h_u_dadda_rca16_fa182_or0[0]), .b(h_u_dadda_rca16_fa96_xor1[0]), .cin(h_u_dadda_rca16_fa97_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa183_xor1), .fa_or0(h_u_dadda_rca16_fa183_or0));
  fa fa_h_u_dadda_rca16_fa184_out(.a(h_u_dadda_rca16_fa183_or0[0]), .b(h_u_dadda_rca16_fa105_xor1[0]), .cin(h_u_dadda_rca16_fa106_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa184_xor1), .fa_or0(h_u_dadda_rca16_fa184_or0));
  fa fa_h_u_dadda_rca16_fa185_out(.a(h_u_dadda_rca16_fa184_or0[0]), .b(h_u_dadda_rca16_fa113_xor1[0]), .cin(h_u_dadda_rca16_fa114_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa185_xor1), .fa_or0(h_u_dadda_rca16_fa185_or0));
  fa fa_h_u_dadda_rca16_fa186_out(.a(h_u_dadda_rca16_fa185_or0[0]), .b(h_u_dadda_rca16_fa120_xor1[0]), .cin(h_u_dadda_rca16_fa121_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa186_xor1), .fa_or0(h_u_dadda_rca16_fa186_or0));
  fa fa_h_u_dadda_rca16_fa187_out(.a(h_u_dadda_rca16_fa186_or0[0]), .b(h_u_dadda_rca16_fa126_xor1[0]), .cin(h_u_dadda_rca16_fa127_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa187_xor1), .fa_or0(h_u_dadda_rca16_fa187_or0));
  fa fa_h_u_dadda_rca16_fa188_out(.a(h_u_dadda_rca16_fa187_or0[0]), .b(h_u_dadda_rca16_fa131_xor1[0]), .cin(h_u_dadda_rca16_fa132_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa188_xor1), .fa_or0(h_u_dadda_rca16_fa188_or0));
  fa fa_h_u_dadda_rca16_fa189_out(.a(h_u_dadda_rca16_fa188_or0[0]), .b(h_u_dadda_rca16_fa135_xor1[0]), .cin(h_u_dadda_rca16_fa136_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa189_xor1), .fa_or0(h_u_dadda_rca16_fa189_or0));
  fa fa_h_u_dadda_rca16_fa190_out(.a(h_u_dadda_rca16_fa189_or0[0]), .b(h_u_dadda_rca16_fa138_xor1[0]), .cin(h_u_dadda_rca16_fa139_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa190_xor1), .fa_or0(h_u_dadda_rca16_fa190_or0));
  fa fa_h_u_dadda_rca16_fa191_out(.a(h_u_dadda_rca16_fa190_or0[0]), .b(h_u_dadda_rca16_fa140_xor1[0]), .cin(h_u_dadda_rca16_fa141_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa191_xor1), .fa_or0(h_u_dadda_rca16_fa191_or0));
  and_gate and_gate_h_u_dadda_rca16_and_12_15(.a(a[12]), .b(b[15]), .out(h_u_dadda_rca16_and_12_15));
  fa fa_h_u_dadda_rca16_fa192_out(.a(h_u_dadda_rca16_fa191_or0[0]), .b(h_u_dadda_rca16_and_12_15[0]), .cin(h_u_dadda_rca16_fa142_xor1[0]), .fa_xor1(h_u_dadda_rca16_fa192_xor1), .fa_or0(h_u_dadda_rca16_fa192_or0));
  and_gate and_gate_h_u_dadda_rca16_and_14_14(.a(a[14]), .b(b[14]), .out(h_u_dadda_rca16_and_14_14));
  and_gate and_gate_h_u_dadda_rca16_and_13_15(.a(a[13]), .b(b[15]), .out(h_u_dadda_rca16_and_13_15));
  fa fa_h_u_dadda_rca16_fa193_out(.a(h_u_dadda_rca16_fa192_or0[0]), .b(h_u_dadda_rca16_and_14_14[0]), .cin(h_u_dadda_rca16_and_13_15[0]), .fa_xor1(h_u_dadda_rca16_fa193_xor1), .fa_or0(h_u_dadda_rca16_fa193_or0));
  and_gate and_gate_h_u_dadda_rca16_and_15_14(.a(a[15]), .b(b[14]), .out(h_u_dadda_rca16_and_15_14));
  fa fa_h_u_dadda_rca16_fa194_out(.a(h_u_dadda_rca16_fa193_or0[0]), .b(h_u_dadda_rca16_fa167_or0[0]), .cin(h_u_dadda_rca16_and_15_14[0]), .fa_xor1(h_u_dadda_rca16_fa194_xor1), .fa_or0(h_u_dadda_rca16_fa194_or0));
  and_gate and_gate_h_u_dadda_rca16_and_0_0(.a(a[0]), .b(b[0]), .out(h_u_dadda_rca16_and_0_0));
  and_gate and_gate_h_u_dadda_rca16_and_1_0(.a(a[1]), .b(b[0]), .out(h_u_dadda_rca16_and_1_0));
  and_gate and_gate_h_u_dadda_rca16_and_0_2(.a(a[0]), .b(b[2]), .out(h_u_dadda_rca16_and_0_2));
  and_gate and_gate_h_u_dadda_rca16_and_14_15(.a(a[14]), .b(b[15]), .out(h_u_dadda_rca16_and_14_15));
  and_gate and_gate_h_u_dadda_rca16_and_0_1(.a(a[0]), .b(b[1]), .out(h_u_dadda_rca16_and_0_1));
  and_gate and_gate_h_u_dadda_rca16_and_15_15(.a(a[15]), .b(b[15]), .out(h_u_dadda_rca16_and_15_15));
  assign h_u_dadda_rca16_u_rca30_a[0] = h_u_dadda_rca16_and_1_0[0];
  assign h_u_dadda_rca16_u_rca30_a[1] = h_u_dadda_rca16_and_0_2[0];
  assign h_u_dadda_rca16_u_rca30_a[2] = h_u_dadda_rca16_ha13_xor0[0];
  assign h_u_dadda_rca16_u_rca30_a[3] = h_u_dadda_rca16_fa143_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[4] = h_u_dadda_rca16_fa144_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[5] = h_u_dadda_rca16_fa145_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[6] = h_u_dadda_rca16_fa146_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[7] = h_u_dadda_rca16_fa147_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[8] = h_u_dadda_rca16_fa148_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[9] = h_u_dadda_rca16_fa149_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[10] = h_u_dadda_rca16_fa150_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[11] = h_u_dadda_rca16_fa151_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[12] = h_u_dadda_rca16_fa152_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[13] = h_u_dadda_rca16_fa153_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[14] = h_u_dadda_rca16_fa154_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[15] = h_u_dadda_rca16_fa155_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[16] = h_u_dadda_rca16_fa156_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[17] = h_u_dadda_rca16_fa157_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[18] = h_u_dadda_rca16_fa158_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[19] = h_u_dadda_rca16_fa159_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[20] = h_u_dadda_rca16_fa160_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[21] = h_u_dadda_rca16_fa161_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[22] = h_u_dadda_rca16_fa162_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[23] = h_u_dadda_rca16_fa163_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[24] = h_u_dadda_rca16_fa164_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[25] = h_u_dadda_rca16_fa165_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[26] = h_u_dadda_rca16_fa166_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[27] = h_u_dadda_rca16_fa167_xor1[0];
  assign h_u_dadda_rca16_u_rca30_a[28] = h_u_dadda_rca16_and_14_15[0];
  assign h_u_dadda_rca16_u_rca30_a[29] = h_u_dadda_rca16_fa194_or0[0];
  assign h_u_dadda_rca16_u_rca30_b[0] = h_u_dadda_rca16_and_0_1[0];
  assign h_u_dadda_rca16_u_rca30_b[1] = h_u_dadda_rca16_ha14_xor0[0];
  assign h_u_dadda_rca16_u_rca30_b[2] = h_u_dadda_rca16_fa168_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[3] = h_u_dadda_rca16_fa169_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[4] = h_u_dadda_rca16_fa170_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[5] = h_u_dadda_rca16_fa171_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[6] = h_u_dadda_rca16_fa172_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[7] = h_u_dadda_rca16_fa173_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[8] = h_u_dadda_rca16_fa174_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[9] = h_u_dadda_rca16_fa175_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[10] = h_u_dadda_rca16_fa176_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[11] = h_u_dadda_rca16_fa177_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[12] = h_u_dadda_rca16_fa178_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[13] = h_u_dadda_rca16_fa179_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[14] = h_u_dadda_rca16_fa180_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[15] = h_u_dadda_rca16_fa181_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[16] = h_u_dadda_rca16_fa182_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[17] = h_u_dadda_rca16_fa183_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[18] = h_u_dadda_rca16_fa184_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[19] = h_u_dadda_rca16_fa185_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[20] = h_u_dadda_rca16_fa186_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[21] = h_u_dadda_rca16_fa187_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[22] = h_u_dadda_rca16_fa188_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[23] = h_u_dadda_rca16_fa189_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[24] = h_u_dadda_rca16_fa190_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[25] = h_u_dadda_rca16_fa191_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[26] = h_u_dadda_rca16_fa192_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[27] = h_u_dadda_rca16_fa193_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[28] = h_u_dadda_rca16_fa194_xor1[0];
  assign h_u_dadda_rca16_u_rca30_b[29] = h_u_dadda_rca16_and_15_15[0];
  u_rca30 u_rca30_h_u_dadda_rca16_u_rca30_out(.a(h_u_dadda_rca16_u_rca30_a), .b(h_u_dadda_rca16_u_rca30_b), .u_rca30_out(h_u_dadda_rca16_u_rca30_out));

  assign h_u_dadda_rca16_out[0] = h_u_dadda_rca16_and_0_0[0];
  assign h_u_dadda_rca16_out[1] = h_u_dadda_rca16_u_rca30_out[0];
  assign h_u_dadda_rca16_out[2] = h_u_dadda_rca16_u_rca30_out[1];
  assign h_u_dadda_rca16_out[3] = h_u_dadda_rca16_u_rca30_out[2];
  assign h_u_dadda_rca16_out[4] = h_u_dadda_rca16_u_rca30_out[3];
  assign h_u_dadda_rca16_out[5] = h_u_dadda_rca16_u_rca30_out[4];
  assign h_u_dadda_rca16_out[6] = h_u_dadda_rca16_u_rca30_out[5];
  assign h_u_dadda_rca16_out[7] = h_u_dadda_rca16_u_rca30_out[6];
  assign h_u_dadda_rca16_out[8] = h_u_dadda_rca16_u_rca30_out[7];
  assign h_u_dadda_rca16_out[9] = h_u_dadda_rca16_u_rca30_out[8];
  assign h_u_dadda_rca16_out[10] = h_u_dadda_rca16_u_rca30_out[9];
  assign h_u_dadda_rca16_out[11] = h_u_dadda_rca16_u_rca30_out[10];
  assign h_u_dadda_rca16_out[12] = h_u_dadda_rca16_u_rca30_out[11];
  assign h_u_dadda_rca16_out[13] = h_u_dadda_rca16_u_rca30_out[12];
  assign h_u_dadda_rca16_out[14] = h_u_dadda_rca16_u_rca30_out[13];
  assign h_u_dadda_rca16_out[15] = h_u_dadda_rca16_u_rca30_out[14];
  assign h_u_dadda_rca16_out[16] = h_u_dadda_rca16_u_rca30_out[15];
  assign h_u_dadda_rca16_out[17] = h_u_dadda_rca16_u_rca30_out[16];
  assign h_u_dadda_rca16_out[18] = h_u_dadda_rca16_u_rca30_out[17];
  assign h_u_dadda_rca16_out[19] = h_u_dadda_rca16_u_rca30_out[18];
  assign h_u_dadda_rca16_out[20] = h_u_dadda_rca16_u_rca30_out[19];
  assign h_u_dadda_rca16_out[21] = h_u_dadda_rca16_u_rca30_out[20];
  assign h_u_dadda_rca16_out[22] = h_u_dadda_rca16_u_rca30_out[21];
  assign h_u_dadda_rca16_out[23] = h_u_dadda_rca16_u_rca30_out[22];
  assign h_u_dadda_rca16_out[24] = h_u_dadda_rca16_u_rca30_out[23];
  assign h_u_dadda_rca16_out[25] = h_u_dadda_rca16_u_rca30_out[24];
  assign h_u_dadda_rca16_out[26] = h_u_dadda_rca16_u_rca30_out[25];
  assign h_u_dadda_rca16_out[27] = h_u_dadda_rca16_u_rca30_out[26];
  assign h_u_dadda_rca16_out[28] = h_u_dadda_rca16_u_rca30_out[27];
  assign h_u_dadda_rca16_out[29] = h_u_dadda_rca16_u_rca30_out[28];
  assign h_u_dadda_rca16_out[30] = h_u_dadda_rca16_u_rca30_out[29];
  assign h_u_dadda_rca16_out[31] = h_u_dadda_rca16_u_rca30_out[30];
endmodule