module f_u_cla4(input [3:0] a, input [3:0] b, output [4:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire constant_wire_value_0_a_0;
  wire constant_wire_value_0_b_0;
  wire constant_wire_value_0_y0;
  wire constant_wire_value_0_y1;
  wire constant_wire_0;
  wire f_u_cla4_pg_logic0_a_0;
  wire f_u_cla4_pg_logic0_b_0;
  wire f_u_cla4_pg_logic0_y0;
  wire f_u_cla4_pg_logic0_y1;
  wire f_u_cla4_pg_logic0_y2;
  wire f_u_cla4_xor0_f_u_cla4_pg_logic0_y2;
  wire f_u_cla4_xor0_constant_wire_0;
  wire f_u_cla4_xor0_y0;
  wire f_u_cla4_and0_f_u_cla4_pg_logic0_y0;
  wire f_u_cla4_and0_constant_wire_0;
  wire f_u_cla4_and0_y0;
  wire f_u_cla4_or0_f_u_cla4_pg_logic0_y1;
  wire f_u_cla4_or0_f_u_cla4_and0_y0;
  wire f_u_cla4_or0_y0;
  wire f_u_cla4_pg_logic1_a_1;
  wire f_u_cla4_pg_logic1_b_1;
  wire f_u_cla4_pg_logic1_y0;
  wire f_u_cla4_pg_logic1_y1;
  wire f_u_cla4_pg_logic1_y2;
  wire f_u_cla4_xor1_f_u_cla4_pg_logic1_y2;
  wire f_u_cla4_xor1_f_u_cla4_or0_y0;
  wire f_u_cla4_xor1_y0;
  wire f_u_cla4_and1_f_u_cla4_pg_logic0_y0;
  wire f_u_cla4_and1_constant_wire_0;
  wire f_u_cla4_and1_y0;
  wire f_u_cla4_and2_f_u_cla4_pg_logic1_y0;
  wire f_u_cla4_and2_constant_wire_0;
  wire f_u_cla4_and2_y0;
  wire f_u_cla4_and3_f_u_cla4_and2_y0;
  wire f_u_cla4_and3_f_u_cla4_and1_y0;
  wire f_u_cla4_and3_y0;
  wire f_u_cla4_and4_f_u_cla4_pg_logic1_y0;
  wire f_u_cla4_and4_f_u_cla4_pg_logic0_y1;
  wire f_u_cla4_and4_y0;
  wire f_u_cla4_or1_f_u_cla4_and4_y0;
  wire f_u_cla4_or1_f_u_cla4_and3_y0;
  wire f_u_cla4_or1_y0;
  wire f_u_cla4_or2_f_u_cla4_pg_logic1_y1;
  wire f_u_cla4_or2_f_u_cla4_or1_y0;
  wire f_u_cla4_or2_y0;
  wire f_u_cla4_pg_logic2_a_2;
  wire f_u_cla4_pg_logic2_b_2;
  wire f_u_cla4_pg_logic2_y0;
  wire f_u_cla4_pg_logic2_y1;
  wire f_u_cla4_pg_logic2_y2;
  wire f_u_cla4_xor2_f_u_cla4_pg_logic2_y2;
  wire f_u_cla4_xor2_f_u_cla4_or2_y0;
  wire f_u_cla4_xor2_y0;
  wire f_u_cla4_and5_f_u_cla4_pg_logic0_y0;
  wire f_u_cla4_and5_constant_wire_0;
  wire f_u_cla4_and5_y0;
  wire f_u_cla4_and6_f_u_cla4_pg_logic1_y0;
  wire f_u_cla4_and6_constant_wire_0;
  wire f_u_cla4_and6_y0;
  wire f_u_cla4_and7_f_u_cla4_and6_y0;
  wire f_u_cla4_and7_f_u_cla4_and5_y0;
  wire f_u_cla4_and7_y0;
  wire f_u_cla4_and8_f_u_cla4_pg_logic2_y0;
  wire f_u_cla4_and8_constant_wire_0;
  wire f_u_cla4_and8_y0;
  wire f_u_cla4_and9_f_u_cla4_and8_y0;
  wire f_u_cla4_and9_f_u_cla4_and7_y0;
  wire f_u_cla4_and9_y0;
  wire f_u_cla4_and10_f_u_cla4_pg_logic1_y0;
  wire f_u_cla4_and10_f_u_cla4_pg_logic0_y1;
  wire f_u_cla4_and10_y0;
  wire f_u_cla4_and11_f_u_cla4_pg_logic2_y0;
  wire f_u_cla4_and11_f_u_cla4_pg_logic0_y1;
  wire f_u_cla4_and11_y0;
  wire f_u_cla4_and12_f_u_cla4_and11_y0;
  wire f_u_cla4_and12_f_u_cla4_and10_y0;
  wire f_u_cla4_and12_y0;
  wire f_u_cla4_and13_f_u_cla4_pg_logic2_y0;
  wire f_u_cla4_and13_f_u_cla4_pg_logic1_y1;
  wire f_u_cla4_and13_y0;
  wire f_u_cla4_or3_f_u_cla4_and13_y0;
  wire f_u_cla4_or3_f_u_cla4_and9_y0;
  wire f_u_cla4_or3_y0;
  wire f_u_cla4_or4_f_u_cla4_or3_y0;
  wire f_u_cla4_or4_f_u_cla4_and12_y0;
  wire f_u_cla4_or4_y0;
  wire f_u_cla4_or5_f_u_cla4_pg_logic2_y1;
  wire f_u_cla4_or5_f_u_cla4_or4_y0;
  wire f_u_cla4_or5_y0;
  wire f_u_cla4_pg_logic3_a_3;
  wire f_u_cla4_pg_logic3_b_3;
  wire f_u_cla4_pg_logic3_y0;
  wire f_u_cla4_pg_logic3_y1;
  wire f_u_cla4_pg_logic3_y2;
  wire f_u_cla4_xor3_f_u_cla4_pg_logic3_y2;
  wire f_u_cla4_xor3_f_u_cla4_or5_y0;
  wire f_u_cla4_xor3_y0;
  wire f_u_cla4_and14_f_u_cla4_pg_logic0_y0;
  wire f_u_cla4_and14_constant_wire_0;
  wire f_u_cla4_and14_y0;
  wire f_u_cla4_and15_f_u_cla4_pg_logic1_y0;
  wire f_u_cla4_and15_constant_wire_0;
  wire f_u_cla4_and15_y0;
  wire f_u_cla4_and16_f_u_cla4_and15_y0;
  wire f_u_cla4_and16_f_u_cla4_and14_y0;
  wire f_u_cla4_and16_y0;
  wire f_u_cla4_and17_f_u_cla4_pg_logic2_y0;
  wire f_u_cla4_and17_constant_wire_0;
  wire f_u_cla4_and17_y0;
  wire f_u_cla4_and18_f_u_cla4_and17_y0;
  wire f_u_cla4_and18_f_u_cla4_and16_y0;
  wire f_u_cla4_and18_y0;
  wire f_u_cla4_and19_f_u_cla4_pg_logic3_y0;
  wire f_u_cla4_and19_constant_wire_0;
  wire f_u_cla4_and19_y0;
  wire f_u_cla4_and20_f_u_cla4_and19_y0;
  wire f_u_cla4_and20_f_u_cla4_and18_y0;
  wire f_u_cla4_and20_y0;
  wire f_u_cla4_and21_f_u_cla4_pg_logic1_y0;
  wire f_u_cla4_and21_f_u_cla4_pg_logic0_y1;
  wire f_u_cla4_and21_y0;
  wire f_u_cla4_and22_f_u_cla4_pg_logic2_y0;
  wire f_u_cla4_and22_f_u_cla4_pg_logic0_y1;
  wire f_u_cla4_and22_y0;
  wire f_u_cla4_and23_f_u_cla4_and22_y0;
  wire f_u_cla4_and23_f_u_cla4_and21_y0;
  wire f_u_cla4_and23_y0;
  wire f_u_cla4_and24_f_u_cla4_pg_logic3_y0;
  wire f_u_cla4_and24_f_u_cla4_pg_logic0_y1;
  wire f_u_cla4_and24_y0;
  wire f_u_cla4_and25_f_u_cla4_and24_y0;
  wire f_u_cla4_and25_f_u_cla4_and23_y0;
  wire f_u_cla4_and25_y0;
  wire f_u_cla4_and26_f_u_cla4_pg_logic2_y0;
  wire f_u_cla4_and26_f_u_cla4_pg_logic1_y1;
  wire f_u_cla4_and26_y0;
  wire f_u_cla4_and27_f_u_cla4_pg_logic3_y0;
  wire f_u_cla4_and27_f_u_cla4_pg_logic1_y1;
  wire f_u_cla4_and27_y0;
  wire f_u_cla4_and28_f_u_cla4_and27_y0;
  wire f_u_cla4_and28_f_u_cla4_and26_y0;
  wire f_u_cla4_and28_y0;
  wire f_u_cla4_and29_f_u_cla4_pg_logic3_y0;
  wire f_u_cla4_and29_f_u_cla4_pg_logic2_y1;
  wire f_u_cla4_and29_y0;
  wire f_u_cla4_or6_f_u_cla4_and29_y0;
  wire f_u_cla4_or6_f_u_cla4_and20_y0;
  wire f_u_cla4_or6_y0;
  wire f_u_cla4_or7_f_u_cla4_or6_y0;
  wire f_u_cla4_or7_f_u_cla4_and25_y0;
  wire f_u_cla4_or7_y0;
  wire f_u_cla4_or8_f_u_cla4_or7_y0;
  wire f_u_cla4_or8_f_u_cla4_and28_y0;
  wire f_u_cla4_or8_y0;
  wire f_u_cla4_or9_f_u_cla4_pg_logic3_y1;
  wire f_u_cla4_or9_f_u_cla4_or8_y0;
  wire f_u_cla4_or9_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign constant_wire_value_0_a_0 = a_0;
  assign constant_wire_value_0_b_0 = b_0;
  assign constant_wire_value_0_y0 = constant_wire_value_0_a_0 ^ constant_wire_value_0_b_0;
  assign constant_wire_value_0_y1 = ~(constant_wire_value_0_a_0 ^ constant_wire_value_0_b_0);
  assign constant_wire_0 = ~(constant_wire_value_0_y0 | constant_wire_value_0_y1);
  assign f_u_cla4_pg_logic0_a_0 = a_0;
  assign f_u_cla4_pg_logic0_b_0 = b_0;
  assign f_u_cla4_pg_logic0_y0 = f_u_cla4_pg_logic0_a_0 | f_u_cla4_pg_logic0_b_0;
  assign f_u_cla4_pg_logic0_y1 = f_u_cla4_pg_logic0_a_0 & f_u_cla4_pg_logic0_b_0;
  assign f_u_cla4_pg_logic0_y2 = f_u_cla4_pg_logic0_a_0 ^ f_u_cla4_pg_logic0_b_0;
  assign f_u_cla4_xor0_f_u_cla4_pg_logic0_y2 = f_u_cla4_pg_logic0_y2;
  assign f_u_cla4_xor0_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_xor0_y0 = f_u_cla4_xor0_f_u_cla4_pg_logic0_y2 ^ f_u_cla4_xor0_constant_wire_0;
  assign f_u_cla4_and0_f_u_cla4_pg_logic0_y0 = f_u_cla4_pg_logic0_y0;
  assign f_u_cla4_and0_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and0_y0 = f_u_cla4_and0_f_u_cla4_pg_logic0_y0 & f_u_cla4_and0_constant_wire_0;
  assign f_u_cla4_or0_f_u_cla4_pg_logic0_y1 = f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_or0_f_u_cla4_and0_y0 = f_u_cla4_and0_y0;
  assign f_u_cla4_or0_y0 = f_u_cla4_or0_f_u_cla4_pg_logic0_y1 | f_u_cla4_or0_f_u_cla4_and0_y0;
  assign f_u_cla4_pg_logic1_a_1 = a_1;
  assign f_u_cla4_pg_logic1_b_1 = b_1;
  assign f_u_cla4_pg_logic1_y0 = f_u_cla4_pg_logic1_a_1 | f_u_cla4_pg_logic1_b_1;
  assign f_u_cla4_pg_logic1_y1 = f_u_cla4_pg_logic1_a_1 & f_u_cla4_pg_logic1_b_1;
  assign f_u_cla4_pg_logic1_y2 = f_u_cla4_pg_logic1_a_1 ^ f_u_cla4_pg_logic1_b_1;
  assign f_u_cla4_xor1_f_u_cla4_pg_logic1_y2 = f_u_cla4_pg_logic1_y2;
  assign f_u_cla4_xor1_f_u_cla4_or0_y0 = f_u_cla4_or0_y0;
  assign f_u_cla4_xor1_y0 = f_u_cla4_xor1_f_u_cla4_pg_logic1_y2 ^ f_u_cla4_xor1_f_u_cla4_or0_y0;
  assign f_u_cla4_and1_f_u_cla4_pg_logic0_y0 = f_u_cla4_pg_logic0_y0;
  assign f_u_cla4_and1_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and1_y0 = f_u_cla4_and1_f_u_cla4_pg_logic0_y0 & f_u_cla4_and1_constant_wire_0;
  assign f_u_cla4_and2_f_u_cla4_pg_logic1_y0 = f_u_cla4_pg_logic1_y0;
  assign f_u_cla4_and2_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and2_y0 = f_u_cla4_and2_f_u_cla4_pg_logic1_y0 & f_u_cla4_and2_constant_wire_0;
  assign f_u_cla4_and3_f_u_cla4_and2_y0 = f_u_cla4_and2_y0;
  assign f_u_cla4_and3_f_u_cla4_and1_y0 = f_u_cla4_and1_y0;
  assign f_u_cla4_and3_y0 = f_u_cla4_and3_f_u_cla4_and2_y0 & f_u_cla4_and3_f_u_cla4_and1_y0;
  assign f_u_cla4_and4_f_u_cla4_pg_logic1_y0 = f_u_cla4_pg_logic1_y0;
  assign f_u_cla4_and4_f_u_cla4_pg_logic0_y1 = f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and4_y0 = f_u_cla4_and4_f_u_cla4_pg_logic1_y0 & f_u_cla4_and4_f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_or1_f_u_cla4_and4_y0 = f_u_cla4_and4_y0;
  assign f_u_cla4_or1_f_u_cla4_and3_y0 = f_u_cla4_and3_y0;
  assign f_u_cla4_or1_y0 = f_u_cla4_or1_f_u_cla4_and4_y0 | f_u_cla4_or1_f_u_cla4_and3_y0;
  assign f_u_cla4_or2_f_u_cla4_pg_logic1_y1 = f_u_cla4_pg_logic1_y1;
  assign f_u_cla4_or2_f_u_cla4_or1_y0 = f_u_cla4_or1_y0;
  assign f_u_cla4_or2_y0 = f_u_cla4_or2_f_u_cla4_pg_logic1_y1 | f_u_cla4_or2_f_u_cla4_or1_y0;
  assign f_u_cla4_pg_logic2_a_2 = a_2;
  assign f_u_cla4_pg_logic2_b_2 = b_2;
  assign f_u_cla4_pg_logic2_y0 = f_u_cla4_pg_logic2_a_2 | f_u_cla4_pg_logic2_b_2;
  assign f_u_cla4_pg_logic2_y1 = f_u_cla4_pg_logic2_a_2 & f_u_cla4_pg_logic2_b_2;
  assign f_u_cla4_pg_logic2_y2 = f_u_cla4_pg_logic2_a_2 ^ f_u_cla4_pg_logic2_b_2;
  assign f_u_cla4_xor2_f_u_cla4_pg_logic2_y2 = f_u_cla4_pg_logic2_y2;
  assign f_u_cla4_xor2_f_u_cla4_or2_y0 = f_u_cla4_or2_y0;
  assign f_u_cla4_xor2_y0 = f_u_cla4_xor2_f_u_cla4_pg_logic2_y2 ^ f_u_cla4_xor2_f_u_cla4_or2_y0;
  assign f_u_cla4_and5_f_u_cla4_pg_logic0_y0 = f_u_cla4_pg_logic0_y0;
  assign f_u_cla4_and5_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and5_y0 = f_u_cla4_and5_f_u_cla4_pg_logic0_y0 & f_u_cla4_and5_constant_wire_0;
  assign f_u_cla4_and6_f_u_cla4_pg_logic1_y0 = f_u_cla4_pg_logic1_y0;
  assign f_u_cla4_and6_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and6_y0 = f_u_cla4_and6_f_u_cla4_pg_logic1_y0 & f_u_cla4_and6_constant_wire_0;
  assign f_u_cla4_and7_f_u_cla4_and6_y0 = f_u_cla4_and6_y0;
  assign f_u_cla4_and7_f_u_cla4_and5_y0 = f_u_cla4_and5_y0;
  assign f_u_cla4_and7_y0 = f_u_cla4_and7_f_u_cla4_and6_y0 & f_u_cla4_and7_f_u_cla4_and5_y0;
  assign f_u_cla4_and8_f_u_cla4_pg_logic2_y0 = f_u_cla4_pg_logic2_y0;
  assign f_u_cla4_and8_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and8_y0 = f_u_cla4_and8_f_u_cla4_pg_logic2_y0 & f_u_cla4_and8_constant_wire_0;
  assign f_u_cla4_and9_f_u_cla4_and8_y0 = f_u_cla4_and8_y0;
  assign f_u_cla4_and9_f_u_cla4_and7_y0 = f_u_cla4_and7_y0;
  assign f_u_cla4_and9_y0 = f_u_cla4_and9_f_u_cla4_and8_y0 & f_u_cla4_and9_f_u_cla4_and7_y0;
  assign f_u_cla4_and10_f_u_cla4_pg_logic1_y0 = f_u_cla4_pg_logic1_y0;
  assign f_u_cla4_and10_f_u_cla4_pg_logic0_y1 = f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and10_y0 = f_u_cla4_and10_f_u_cla4_pg_logic1_y0 & f_u_cla4_and10_f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and11_f_u_cla4_pg_logic2_y0 = f_u_cla4_pg_logic2_y0;
  assign f_u_cla4_and11_f_u_cla4_pg_logic0_y1 = f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and11_y0 = f_u_cla4_and11_f_u_cla4_pg_logic2_y0 & f_u_cla4_and11_f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and12_f_u_cla4_and11_y0 = f_u_cla4_and11_y0;
  assign f_u_cla4_and12_f_u_cla4_and10_y0 = f_u_cla4_and10_y0;
  assign f_u_cla4_and12_y0 = f_u_cla4_and12_f_u_cla4_and11_y0 & f_u_cla4_and12_f_u_cla4_and10_y0;
  assign f_u_cla4_and13_f_u_cla4_pg_logic2_y0 = f_u_cla4_pg_logic2_y0;
  assign f_u_cla4_and13_f_u_cla4_pg_logic1_y1 = f_u_cla4_pg_logic1_y1;
  assign f_u_cla4_and13_y0 = f_u_cla4_and13_f_u_cla4_pg_logic2_y0 & f_u_cla4_and13_f_u_cla4_pg_logic1_y1;
  assign f_u_cla4_or3_f_u_cla4_and13_y0 = f_u_cla4_and13_y0;
  assign f_u_cla4_or3_f_u_cla4_and9_y0 = f_u_cla4_and9_y0;
  assign f_u_cla4_or3_y0 = f_u_cla4_or3_f_u_cla4_and13_y0 | f_u_cla4_or3_f_u_cla4_and9_y0;
  assign f_u_cla4_or4_f_u_cla4_or3_y0 = f_u_cla4_or3_y0;
  assign f_u_cla4_or4_f_u_cla4_and12_y0 = f_u_cla4_and12_y0;
  assign f_u_cla4_or4_y0 = f_u_cla4_or4_f_u_cla4_or3_y0 | f_u_cla4_or4_f_u_cla4_and12_y0;
  assign f_u_cla4_or5_f_u_cla4_pg_logic2_y1 = f_u_cla4_pg_logic2_y1;
  assign f_u_cla4_or5_f_u_cla4_or4_y0 = f_u_cla4_or4_y0;
  assign f_u_cla4_or5_y0 = f_u_cla4_or5_f_u_cla4_pg_logic2_y1 | f_u_cla4_or5_f_u_cla4_or4_y0;
  assign f_u_cla4_pg_logic3_a_3 = a_3;
  assign f_u_cla4_pg_logic3_b_3 = b_3;
  assign f_u_cla4_pg_logic3_y0 = f_u_cla4_pg_logic3_a_3 | f_u_cla4_pg_logic3_b_3;
  assign f_u_cla4_pg_logic3_y1 = f_u_cla4_pg_logic3_a_3 & f_u_cla4_pg_logic3_b_3;
  assign f_u_cla4_pg_logic3_y2 = f_u_cla4_pg_logic3_a_3 ^ f_u_cla4_pg_logic3_b_3;
  assign f_u_cla4_xor3_f_u_cla4_pg_logic3_y2 = f_u_cla4_pg_logic3_y2;
  assign f_u_cla4_xor3_f_u_cla4_or5_y0 = f_u_cla4_or5_y0;
  assign f_u_cla4_xor3_y0 = f_u_cla4_xor3_f_u_cla4_pg_logic3_y2 ^ f_u_cla4_xor3_f_u_cla4_or5_y0;
  assign f_u_cla4_and14_f_u_cla4_pg_logic0_y0 = f_u_cla4_pg_logic0_y0;
  assign f_u_cla4_and14_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and14_y0 = f_u_cla4_and14_f_u_cla4_pg_logic0_y0 & f_u_cla4_and14_constant_wire_0;
  assign f_u_cla4_and15_f_u_cla4_pg_logic1_y0 = f_u_cla4_pg_logic1_y0;
  assign f_u_cla4_and15_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and15_y0 = f_u_cla4_and15_f_u_cla4_pg_logic1_y0 & f_u_cla4_and15_constant_wire_0;
  assign f_u_cla4_and16_f_u_cla4_and15_y0 = f_u_cla4_and15_y0;
  assign f_u_cla4_and16_f_u_cla4_and14_y0 = f_u_cla4_and14_y0;
  assign f_u_cla4_and16_y0 = f_u_cla4_and16_f_u_cla4_and15_y0 & f_u_cla4_and16_f_u_cla4_and14_y0;
  assign f_u_cla4_and17_f_u_cla4_pg_logic2_y0 = f_u_cla4_pg_logic2_y0;
  assign f_u_cla4_and17_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and17_y0 = f_u_cla4_and17_f_u_cla4_pg_logic2_y0 & f_u_cla4_and17_constant_wire_0;
  assign f_u_cla4_and18_f_u_cla4_and17_y0 = f_u_cla4_and17_y0;
  assign f_u_cla4_and18_f_u_cla4_and16_y0 = f_u_cla4_and16_y0;
  assign f_u_cla4_and18_y0 = f_u_cla4_and18_f_u_cla4_and17_y0 & f_u_cla4_and18_f_u_cla4_and16_y0;
  assign f_u_cla4_and19_f_u_cla4_pg_logic3_y0 = f_u_cla4_pg_logic3_y0;
  assign f_u_cla4_and19_constant_wire_0 = constant_wire_0;
  assign f_u_cla4_and19_y0 = f_u_cla4_and19_f_u_cla4_pg_logic3_y0 & f_u_cla4_and19_constant_wire_0;
  assign f_u_cla4_and20_f_u_cla4_and19_y0 = f_u_cla4_and19_y0;
  assign f_u_cla4_and20_f_u_cla4_and18_y0 = f_u_cla4_and18_y0;
  assign f_u_cla4_and20_y0 = f_u_cla4_and20_f_u_cla4_and19_y0 & f_u_cla4_and20_f_u_cla4_and18_y0;
  assign f_u_cla4_and21_f_u_cla4_pg_logic1_y0 = f_u_cla4_pg_logic1_y0;
  assign f_u_cla4_and21_f_u_cla4_pg_logic0_y1 = f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and21_y0 = f_u_cla4_and21_f_u_cla4_pg_logic1_y0 & f_u_cla4_and21_f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and22_f_u_cla4_pg_logic2_y0 = f_u_cla4_pg_logic2_y0;
  assign f_u_cla4_and22_f_u_cla4_pg_logic0_y1 = f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and22_y0 = f_u_cla4_and22_f_u_cla4_pg_logic2_y0 & f_u_cla4_and22_f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and23_f_u_cla4_and22_y0 = f_u_cla4_and22_y0;
  assign f_u_cla4_and23_f_u_cla4_and21_y0 = f_u_cla4_and21_y0;
  assign f_u_cla4_and23_y0 = f_u_cla4_and23_f_u_cla4_and22_y0 & f_u_cla4_and23_f_u_cla4_and21_y0;
  assign f_u_cla4_and24_f_u_cla4_pg_logic3_y0 = f_u_cla4_pg_logic3_y0;
  assign f_u_cla4_and24_f_u_cla4_pg_logic0_y1 = f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and24_y0 = f_u_cla4_and24_f_u_cla4_pg_logic3_y0 & f_u_cla4_and24_f_u_cla4_pg_logic0_y1;
  assign f_u_cla4_and25_f_u_cla4_and24_y0 = f_u_cla4_and24_y0;
  assign f_u_cla4_and25_f_u_cla4_and23_y0 = f_u_cla4_and23_y0;
  assign f_u_cla4_and25_y0 = f_u_cla4_and25_f_u_cla4_and24_y0 & f_u_cla4_and25_f_u_cla4_and23_y0;
  assign f_u_cla4_and26_f_u_cla4_pg_logic2_y0 = f_u_cla4_pg_logic2_y0;
  assign f_u_cla4_and26_f_u_cla4_pg_logic1_y1 = f_u_cla4_pg_logic1_y1;
  assign f_u_cla4_and26_y0 = f_u_cla4_and26_f_u_cla4_pg_logic2_y0 & f_u_cla4_and26_f_u_cla4_pg_logic1_y1;
  assign f_u_cla4_and27_f_u_cla4_pg_logic3_y0 = f_u_cla4_pg_logic3_y0;
  assign f_u_cla4_and27_f_u_cla4_pg_logic1_y1 = f_u_cla4_pg_logic1_y1;
  assign f_u_cla4_and27_y0 = f_u_cla4_and27_f_u_cla4_pg_logic3_y0 & f_u_cla4_and27_f_u_cla4_pg_logic1_y1;
  assign f_u_cla4_and28_f_u_cla4_and27_y0 = f_u_cla4_and27_y0;
  assign f_u_cla4_and28_f_u_cla4_and26_y0 = f_u_cla4_and26_y0;
  assign f_u_cla4_and28_y0 = f_u_cla4_and28_f_u_cla4_and27_y0 & f_u_cla4_and28_f_u_cla4_and26_y0;
  assign f_u_cla4_and29_f_u_cla4_pg_logic3_y0 = f_u_cla4_pg_logic3_y0;
  assign f_u_cla4_and29_f_u_cla4_pg_logic2_y1 = f_u_cla4_pg_logic2_y1;
  assign f_u_cla4_and29_y0 = f_u_cla4_and29_f_u_cla4_pg_logic3_y0 & f_u_cla4_and29_f_u_cla4_pg_logic2_y1;
  assign f_u_cla4_or6_f_u_cla4_and29_y0 = f_u_cla4_and29_y0;
  assign f_u_cla4_or6_f_u_cla4_and20_y0 = f_u_cla4_and20_y0;
  assign f_u_cla4_or6_y0 = f_u_cla4_or6_f_u_cla4_and29_y0 | f_u_cla4_or6_f_u_cla4_and20_y0;
  assign f_u_cla4_or7_f_u_cla4_or6_y0 = f_u_cla4_or6_y0;
  assign f_u_cla4_or7_f_u_cla4_and25_y0 = f_u_cla4_and25_y0;
  assign f_u_cla4_or7_y0 = f_u_cla4_or7_f_u_cla4_or6_y0 | f_u_cla4_or7_f_u_cla4_and25_y0;
  assign f_u_cla4_or8_f_u_cla4_or7_y0 = f_u_cla4_or7_y0;
  assign f_u_cla4_or8_f_u_cla4_and28_y0 = f_u_cla4_and28_y0;
  assign f_u_cla4_or8_y0 = f_u_cla4_or8_f_u_cla4_or7_y0 | f_u_cla4_or8_f_u_cla4_and28_y0;
  assign f_u_cla4_or9_f_u_cla4_pg_logic3_y1 = f_u_cla4_pg_logic3_y1;
  assign f_u_cla4_or9_f_u_cla4_or8_y0 = f_u_cla4_or8_y0;
  assign f_u_cla4_or9_y0 = f_u_cla4_or9_f_u_cla4_pg_logic3_y1 | f_u_cla4_or9_f_u_cla4_or8_y0;

  assign out[0] = f_u_cla4_xor0_y0;
  assign out[1] = f_u_cla4_xor1_y0;
  assign out[2] = f_u_cla4_xor2_y0;
  assign out[3] = f_u_cla4_xor3_y0;
  assign out[4] = f_u_cla4_or9_y0;
endmodule