module s_CSAwallace_rca16(input [15:0] a, input [15:0] b, output [31:0] s_CSAwallace_rca16_out);
  wire s_CSAwallace_rca16_and_0_0;
  wire s_CSAwallace_rca16_and_1_0;
  wire s_CSAwallace_rca16_and_2_0;
  wire s_CSAwallace_rca16_and_3_0;
  wire s_CSAwallace_rca16_and_4_0;
  wire s_CSAwallace_rca16_and_5_0;
  wire s_CSAwallace_rca16_and_6_0;
  wire s_CSAwallace_rca16_and_7_0;
  wire s_CSAwallace_rca16_and_8_0;
  wire s_CSAwallace_rca16_and_9_0;
  wire s_CSAwallace_rca16_and_10_0;
  wire s_CSAwallace_rca16_and_11_0;
  wire s_CSAwallace_rca16_and_12_0;
  wire s_CSAwallace_rca16_and_13_0;
  wire s_CSAwallace_rca16_and_14_0;
  wire s_CSAwallace_rca16_nand_15_0;
  wire s_CSAwallace_rca16_and_0_1;
  wire s_CSAwallace_rca16_and_1_1;
  wire s_CSAwallace_rca16_and_2_1;
  wire s_CSAwallace_rca16_and_3_1;
  wire s_CSAwallace_rca16_and_4_1;
  wire s_CSAwallace_rca16_and_5_1;
  wire s_CSAwallace_rca16_and_6_1;
  wire s_CSAwallace_rca16_and_7_1;
  wire s_CSAwallace_rca16_and_8_1;
  wire s_CSAwallace_rca16_and_9_1;
  wire s_CSAwallace_rca16_and_10_1;
  wire s_CSAwallace_rca16_and_11_1;
  wire s_CSAwallace_rca16_and_12_1;
  wire s_CSAwallace_rca16_and_13_1;
  wire s_CSAwallace_rca16_and_14_1;
  wire s_CSAwallace_rca16_nand_15_1;
  wire s_CSAwallace_rca16_and_0_2;
  wire s_CSAwallace_rca16_and_1_2;
  wire s_CSAwallace_rca16_and_2_2;
  wire s_CSAwallace_rca16_and_3_2;
  wire s_CSAwallace_rca16_and_4_2;
  wire s_CSAwallace_rca16_and_5_2;
  wire s_CSAwallace_rca16_and_6_2;
  wire s_CSAwallace_rca16_and_7_2;
  wire s_CSAwallace_rca16_and_8_2;
  wire s_CSAwallace_rca16_and_9_2;
  wire s_CSAwallace_rca16_and_10_2;
  wire s_CSAwallace_rca16_and_11_2;
  wire s_CSAwallace_rca16_and_12_2;
  wire s_CSAwallace_rca16_and_13_2;
  wire s_CSAwallace_rca16_and_14_2;
  wire s_CSAwallace_rca16_nand_15_2;
  wire s_CSAwallace_rca16_and_0_3;
  wire s_CSAwallace_rca16_and_1_3;
  wire s_CSAwallace_rca16_and_2_3;
  wire s_CSAwallace_rca16_and_3_3;
  wire s_CSAwallace_rca16_and_4_3;
  wire s_CSAwallace_rca16_and_5_3;
  wire s_CSAwallace_rca16_and_6_3;
  wire s_CSAwallace_rca16_and_7_3;
  wire s_CSAwallace_rca16_and_8_3;
  wire s_CSAwallace_rca16_and_9_3;
  wire s_CSAwallace_rca16_and_10_3;
  wire s_CSAwallace_rca16_and_11_3;
  wire s_CSAwallace_rca16_and_12_3;
  wire s_CSAwallace_rca16_and_13_3;
  wire s_CSAwallace_rca16_and_14_3;
  wire s_CSAwallace_rca16_nand_15_3;
  wire s_CSAwallace_rca16_and_0_4;
  wire s_CSAwallace_rca16_and_1_4;
  wire s_CSAwallace_rca16_and_2_4;
  wire s_CSAwallace_rca16_and_3_4;
  wire s_CSAwallace_rca16_and_4_4;
  wire s_CSAwallace_rca16_and_5_4;
  wire s_CSAwallace_rca16_and_6_4;
  wire s_CSAwallace_rca16_and_7_4;
  wire s_CSAwallace_rca16_and_8_4;
  wire s_CSAwallace_rca16_and_9_4;
  wire s_CSAwallace_rca16_and_10_4;
  wire s_CSAwallace_rca16_and_11_4;
  wire s_CSAwallace_rca16_and_12_4;
  wire s_CSAwallace_rca16_and_13_4;
  wire s_CSAwallace_rca16_and_14_4;
  wire s_CSAwallace_rca16_nand_15_4;
  wire s_CSAwallace_rca16_and_0_5;
  wire s_CSAwallace_rca16_and_1_5;
  wire s_CSAwallace_rca16_and_2_5;
  wire s_CSAwallace_rca16_and_3_5;
  wire s_CSAwallace_rca16_and_4_5;
  wire s_CSAwallace_rca16_and_5_5;
  wire s_CSAwallace_rca16_and_6_5;
  wire s_CSAwallace_rca16_and_7_5;
  wire s_CSAwallace_rca16_and_8_5;
  wire s_CSAwallace_rca16_and_9_5;
  wire s_CSAwallace_rca16_and_10_5;
  wire s_CSAwallace_rca16_and_11_5;
  wire s_CSAwallace_rca16_and_12_5;
  wire s_CSAwallace_rca16_and_13_5;
  wire s_CSAwallace_rca16_and_14_5;
  wire s_CSAwallace_rca16_nand_15_5;
  wire s_CSAwallace_rca16_and_0_6;
  wire s_CSAwallace_rca16_and_1_6;
  wire s_CSAwallace_rca16_and_2_6;
  wire s_CSAwallace_rca16_and_3_6;
  wire s_CSAwallace_rca16_and_4_6;
  wire s_CSAwallace_rca16_and_5_6;
  wire s_CSAwallace_rca16_and_6_6;
  wire s_CSAwallace_rca16_and_7_6;
  wire s_CSAwallace_rca16_and_8_6;
  wire s_CSAwallace_rca16_and_9_6;
  wire s_CSAwallace_rca16_and_10_6;
  wire s_CSAwallace_rca16_and_11_6;
  wire s_CSAwallace_rca16_and_12_6;
  wire s_CSAwallace_rca16_and_13_6;
  wire s_CSAwallace_rca16_and_14_6;
  wire s_CSAwallace_rca16_nand_15_6;
  wire s_CSAwallace_rca16_and_0_7;
  wire s_CSAwallace_rca16_and_1_7;
  wire s_CSAwallace_rca16_and_2_7;
  wire s_CSAwallace_rca16_and_3_7;
  wire s_CSAwallace_rca16_and_4_7;
  wire s_CSAwallace_rca16_and_5_7;
  wire s_CSAwallace_rca16_and_6_7;
  wire s_CSAwallace_rca16_and_7_7;
  wire s_CSAwallace_rca16_and_8_7;
  wire s_CSAwallace_rca16_and_9_7;
  wire s_CSAwallace_rca16_and_10_7;
  wire s_CSAwallace_rca16_and_11_7;
  wire s_CSAwallace_rca16_and_12_7;
  wire s_CSAwallace_rca16_and_13_7;
  wire s_CSAwallace_rca16_and_14_7;
  wire s_CSAwallace_rca16_nand_15_7;
  wire s_CSAwallace_rca16_and_0_8;
  wire s_CSAwallace_rca16_and_1_8;
  wire s_CSAwallace_rca16_and_2_8;
  wire s_CSAwallace_rca16_and_3_8;
  wire s_CSAwallace_rca16_and_4_8;
  wire s_CSAwallace_rca16_and_5_8;
  wire s_CSAwallace_rca16_and_6_8;
  wire s_CSAwallace_rca16_and_7_8;
  wire s_CSAwallace_rca16_and_8_8;
  wire s_CSAwallace_rca16_and_9_8;
  wire s_CSAwallace_rca16_and_10_8;
  wire s_CSAwallace_rca16_and_11_8;
  wire s_CSAwallace_rca16_and_12_8;
  wire s_CSAwallace_rca16_and_13_8;
  wire s_CSAwallace_rca16_and_14_8;
  wire s_CSAwallace_rca16_nand_15_8;
  wire s_CSAwallace_rca16_and_0_9;
  wire s_CSAwallace_rca16_and_1_9;
  wire s_CSAwallace_rca16_and_2_9;
  wire s_CSAwallace_rca16_and_3_9;
  wire s_CSAwallace_rca16_and_4_9;
  wire s_CSAwallace_rca16_and_5_9;
  wire s_CSAwallace_rca16_and_6_9;
  wire s_CSAwallace_rca16_and_7_9;
  wire s_CSAwallace_rca16_and_8_9;
  wire s_CSAwallace_rca16_and_9_9;
  wire s_CSAwallace_rca16_and_10_9;
  wire s_CSAwallace_rca16_and_11_9;
  wire s_CSAwallace_rca16_and_12_9;
  wire s_CSAwallace_rca16_and_13_9;
  wire s_CSAwallace_rca16_and_14_9;
  wire s_CSAwallace_rca16_nand_15_9;
  wire s_CSAwallace_rca16_and_0_10;
  wire s_CSAwallace_rca16_and_1_10;
  wire s_CSAwallace_rca16_and_2_10;
  wire s_CSAwallace_rca16_and_3_10;
  wire s_CSAwallace_rca16_and_4_10;
  wire s_CSAwallace_rca16_and_5_10;
  wire s_CSAwallace_rca16_and_6_10;
  wire s_CSAwallace_rca16_and_7_10;
  wire s_CSAwallace_rca16_and_8_10;
  wire s_CSAwallace_rca16_and_9_10;
  wire s_CSAwallace_rca16_and_10_10;
  wire s_CSAwallace_rca16_and_11_10;
  wire s_CSAwallace_rca16_and_12_10;
  wire s_CSAwallace_rca16_and_13_10;
  wire s_CSAwallace_rca16_and_14_10;
  wire s_CSAwallace_rca16_nand_15_10;
  wire s_CSAwallace_rca16_and_0_11;
  wire s_CSAwallace_rca16_and_1_11;
  wire s_CSAwallace_rca16_and_2_11;
  wire s_CSAwallace_rca16_and_3_11;
  wire s_CSAwallace_rca16_and_4_11;
  wire s_CSAwallace_rca16_and_5_11;
  wire s_CSAwallace_rca16_and_6_11;
  wire s_CSAwallace_rca16_and_7_11;
  wire s_CSAwallace_rca16_and_8_11;
  wire s_CSAwallace_rca16_and_9_11;
  wire s_CSAwallace_rca16_and_10_11;
  wire s_CSAwallace_rca16_and_11_11;
  wire s_CSAwallace_rca16_and_12_11;
  wire s_CSAwallace_rca16_and_13_11;
  wire s_CSAwallace_rca16_and_14_11;
  wire s_CSAwallace_rca16_nand_15_11;
  wire s_CSAwallace_rca16_and_0_12;
  wire s_CSAwallace_rca16_and_1_12;
  wire s_CSAwallace_rca16_and_2_12;
  wire s_CSAwallace_rca16_and_3_12;
  wire s_CSAwallace_rca16_and_4_12;
  wire s_CSAwallace_rca16_and_5_12;
  wire s_CSAwallace_rca16_and_6_12;
  wire s_CSAwallace_rca16_and_7_12;
  wire s_CSAwallace_rca16_and_8_12;
  wire s_CSAwallace_rca16_and_9_12;
  wire s_CSAwallace_rca16_and_10_12;
  wire s_CSAwallace_rca16_and_11_12;
  wire s_CSAwallace_rca16_and_12_12;
  wire s_CSAwallace_rca16_and_13_12;
  wire s_CSAwallace_rca16_and_14_12;
  wire s_CSAwallace_rca16_nand_15_12;
  wire s_CSAwallace_rca16_and_0_13;
  wire s_CSAwallace_rca16_and_1_13;
  wire s_CSAwallace_rca16_and_2_13;
  wire s_CSAwallace_rca16_and_3_13;
  wire s_CSAwallace_rca16_and_4_13;
  wire s_CSAwallace_rca16_and_5_13;
  wire s_CSAwallace_rca16_and_6_13;
  wire s_CSAwallace_rca16_and_7_13;
  wire s_CSAwallace_rca16_and_8_13;
  wire s_CSAwallace_rca16_and_9_13;
  wire s_CSAwallace_rca16_and_10_13;
  wire s_CSAwallace_rca16_and_11_13;
  wire s_CSAwallace_rca16_and_12_13;
  wire s_CSAwallace_rca16_and_13_13;
  wire s_CSAwallace_rca16_and_14_13;
  wire s_CSAwallace_rca16_nand_15_13;
  wire s_CSAwallace_rca16_and_0_14;
  wire s_CSAwallace_rca16_and_1_14;
  wire s_CSAwallace_rca16_and_2_14;
  wire s_CSAwallace_rca16_and_3_14;
  wire s_CSAwallace_rca16_and_4_14;
  wire s_CSAwallace_rca16_and_5_14;
  wire s_CSAwallace_rca16_and_6_14;
  wire s_CSAwallace_rca16_and_7_14;
  wire s_CSAwallace_rca16_and_8_14;
  wire s_CSAwallace_rca16_and_9_14;
  wire s_CSAwallace_rca16_and_10_14;
  wire s_CSAwallace_rca16_and_11_14;
  wire s_CSAwallace_rca16_and_12_14;
  wire s_CSAwallace_rca16_and_13_14;
  wire s_CSAwallace_rca16_and_14_14;
  wire s_CSAwallace_rca16_nand_15_14;
  wire s_CSAwallace_rca16_nand_0_15;
  wire s_CSAwallace_rca16_nand_1_15;
  wire s_CSAwallace_rca16_nand_2_15;
  wire s_CSAwallace_rca16_nand_3_15;
  wire s_CSAwallace_rca16_nand_4_15;
  wire s_CSAwallace_rca16_nand_5_15;
  wire s_CSAwallace_rca16_nand_6_15;
  wire s_CSAwallace_rca16_nand_7_15;
  wire s_CSAwallace_rca16_nand_8_15;
  wire s_CSAwallace_rca16_nand_9_15;
  wire s_CSAwallace_rca16_nand_10_15;
  wire s_CSAwallace_rca16_nand_11_15;
  wire s_CSAwallace_rca16_nand_12_15;
  wire s_CSAwallace_rca16_nand_13_15;
  wire s_CSAwallace_rca16_nand_14_15;
  wire s_CSAwallace_rca16_and_15_15;
  wire s_CSAwallace_rca16_csa0_csa_component_fa1_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa1_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa2_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa2_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa2_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa2_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa2_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa3_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa3_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa3_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa3_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa3_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa4_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa4_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa4_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa4_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa4_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa5_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa5_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa5_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa5_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa5_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa6_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa6_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa6_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa6_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa6_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa7_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa7_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa7_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa7_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa7_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa8_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa8_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa8_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa8_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa8_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa9_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa9_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa9_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa10_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa10_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa10_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa11_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa11_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa11_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa0_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa0_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa4_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa4_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa5_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa5_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa5_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa5_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa5_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa6_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa6_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa6_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa6_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa6_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa7_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa7_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa7_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa7_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa7_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa8_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa8_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa8_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa8_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa8_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa9_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa9_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa9_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa10_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa10_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa10_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa11_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa11_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa11_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa1_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa1_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa7_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa7_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa8_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa8_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa8_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa8_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa8_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa9_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa9_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa9_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa10_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa10_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa10_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa11_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa11_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa11_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa21_and0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa2_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa2_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa11_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa11_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa11_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa21_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa22_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa23_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa23_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa23_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa23_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa23_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa24_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa24_and0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa24_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa24_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa24_or0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa25_xor0;
  wire s_CSAwallace_rca16_csa3_csa_component_fa25_xor1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa25_and1;
  wire s_CSAwallace_rca16_csa3_csa_component_fa25_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa21_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa22_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa23_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa23_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa23_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa23_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa23_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa24_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa24_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa24_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa24_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa24_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa25_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa25_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa25_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa25_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa25_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa26_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa26_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa26_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa26_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa26_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa27_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa27_and0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa27_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa27_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa27_or0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa28_xor0;
  wire s_CSAwallace_rca16_csa4_csa_component_fa28_xor1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa28_and1;
  wire s_CSAwallace_rca16_csa4_csa_component_fa28_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa2_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa2_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa3_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa3_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa3_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa3_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa3_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa4_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa4_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa4_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa4_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa4_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa5_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa5_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa5_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa5_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa5_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa6_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa6_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa6_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa6_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa6_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa7_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa7_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa7_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa7_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa7_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa8_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa8_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa8_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa8_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa8_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa9_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa9_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa9_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa10_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa10_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa10_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa11_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa11_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa11_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa5_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa5_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa6_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa6_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa7_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa7_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa8_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa8_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa8_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa8_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa8_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa9_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa9_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa9_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa10_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa10_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa10_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa11_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa11_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa11_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa23_xor0;
  wire s_CSAwallace_rca16_csa6_csa_component_fa23_xor1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa23_and1;
  wire s_CSAwallace_rca16_csa6_csa_component_fa23_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa21_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa22_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa23_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa23_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa23_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa23_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa23_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa24_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa24_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa24_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa24_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa24_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa25_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa25_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa25_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa25_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa25_or0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa26_xor0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa26_and0;
  wire s_CSAwallace_rca16_csa7_csa_component_fa26_xor1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa26_and1;
  wire s_CSAwallace_rca16_csa7_csa_component_fa26_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa3_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa3_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa4_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa4_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa5_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa5_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa5_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa5_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa5_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa6_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa6_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa6_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa6_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa6_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa7_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa7_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa7_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa7_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa7_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa8_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa8_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa8_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa8_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa8_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa9_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa9_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa9_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa10_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa10_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa10_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa11_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa11_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa11_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa8_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa8_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa21_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa22_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa23_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa23_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa23_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa23_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa23_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa24_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa24_and0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa24_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa24_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa24_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa25_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa25_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa25_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa25_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa26_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa26_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa26_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa26_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa27_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa27_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa27_and1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa27_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa28_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa28_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa28_or0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa29_xor0;
  wire s_CSAwallace_rca16_csa9_csa_component_fa29_xor1;
  wire s_CSAwallace_rca16_csa9_csa_component_fa29_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa4_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa4_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa5_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa5_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa6_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa6_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa7_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa7_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa7_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa7_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa7_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa8_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa8_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa8_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa8_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa8_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa9_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa9_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa9_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa10_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa10_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa10_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa11_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa11_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa11_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa21_and0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa23_xor0;
  wire s_CSAwallace_rca16_csa10_csa_component_fa23_xor1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa23_and1;
  wire s_CSAwallace_rca16_csa10_csa_component_fa23_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa21_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa22_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa23_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa23_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa23_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa23_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa23_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa24_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa24_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa24_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa24_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa24_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa25_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa25_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa25_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa25_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa25_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa26_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa26_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa26_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa26_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa26_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa27_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa27_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa27_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa27_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa27_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa28_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa28_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa28_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa28_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa28_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa29_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa29_and0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa29_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa29_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa29_or0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa30_xor0;
  wire s_CSAwallace_rca16_csa11_csa_component_fa30_xor1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa30_and1;
  wire s_CSAwallace_rca16_csa11_csa_component_fa30_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa5_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa5_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa6_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa6_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa7_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa7_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa8_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa8_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa10_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa10_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa10_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa11_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa11_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa11_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa12_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa12_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa12_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa13_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa13_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa13_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa14_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa14_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa14_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa21_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa22_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa23_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa23_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa23_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa23_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa23_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa24_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa24_and0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa24_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa24_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa24_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa25_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa25_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa25_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa25_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa26_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa26_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa26_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa26_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa27_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa27_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa27_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa27_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa28_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa28_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa28_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa28_or0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa29_xor0;
  wire s_CSAwallace_rca16_csa12_csa_component_fa29_xor1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa29_and1;
  wire s_CSAwallace_rca16_csa12_csa_component_fa29_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa6_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa6_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa7_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa7_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa8_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa8_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa9_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa9_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa10_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa10_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa11_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa11_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa12_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa12_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa13_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa13_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa14_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa14_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa15_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa15_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa15_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa15_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa15_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa16_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa16_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa16_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa16_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa16_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa17_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa17_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa17_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa17_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa17_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa18_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa18_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa18_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa18_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa18_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa19_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa19_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa19_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa19_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa19_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa20_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa20_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa20_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa20_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa20_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa21_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa21_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa21_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa21_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa21_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa22_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa22_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa22_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa22_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa22_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa23_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa23_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa23_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa23_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa23_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa24_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa24_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa24_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa24_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa24_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa25_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa25_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa25_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa25_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa25_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa26_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa26_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa26_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa26_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa26_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa27_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa27_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa27_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa27_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa27_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa28_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa28_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa28_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa28_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa28_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa29_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa29_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa29_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa29_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa29_or0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa30_xor0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa30_and0;
  wire s_CSAwallace_rca16_csa13_csa_component_fa30_xor1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa30_and1;
  wire s_CSAwallace_rca16_csa13_csa_component_fa30_or0;
  wire s_CSAwallace_rca16_u_rca32_fa7_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa7_and0;
  wire s_CSAwallace_rca16_u_rca32_fa8_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa8_and0;
  wire s_CSAwallace_rca16_u_rca32_fa8_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa8_and1;
  wire s_CSAwallace_rca16_u_rca32_fa8_or0;
  wire s_CSAwallace_rca16_u_rca32_fa9_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa9_and0;
  wire s_CSAwallace_rca16_u_rca32_fa9_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa9_and1;
  wire s_CSAwallace_rca16_u_rca32_fa9_or0;
  wire s_CSAwallace_rca16_u_rca32_fa10_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa10_and0;
  wire s_CSAwallace_rca16_u_rca32_fa10_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa10_and1;
  wire s_CSAwallace_rca16_u_rca32_fa10_or0;
  wire s_CSAwallace_rca16_u_rca32_fa11_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa11_and0;
  wire s_CSAwallace_rca16_u_rca32_fa11_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa11_and1;
  wire s_CSAwallace_rca16_u_rca32_fa11_or0;
  wire s_CSAwallace_rca16_u_rca32_fa12_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa12_and0;
  wire s_CSAwallace_rca16_u_rca32_fa12_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa12_and1;
  wire s_CSAwallace_rca16_u_rca32_fa12_or0;
  wire s_CSAwallace_rca16_u_rca32_fa13_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa13_and0;
  wire s_CSAwallace_rca16_u_rca32_fa13_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa13_and1;
  wire s_CSAwallace_rca16_u_rca32_fa13_or0;
  wire s_CSAwallace_rca16_u_rca32_fa14_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa14_and0;
  wire s_CSAwallace_rca16_u_rca32_fa14_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa14_and1;
  wire s_CSAwallace_rca16_u_rca32_fa14_or0;
  wire s_CSAwallace_rca16_u_rca32_fa15_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa15_and0;
  wire s_CSAwallace_rca16_u_rca32_fa15_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa15_and1;
  wire s_CSAwallace_rca16_u_rca32_fa15_or0;
  wire s_CSAwallace_rca16_u_rca32_fa16_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa16_and0;
  wire s_CSAwallace_rca16_u_rca32_fa16_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa16_and1;
  wire s_CSAwallace_rca16_u_rca32_fa16_or0;
  wire s_CSAwallace_rca16_u_rca32_fa17_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa17_and0;
  wire s_CSAwallace_rca16_u_rca32_fa17_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa17_and1;
  wire s_CSAwallace_rca16_u_rca32_fa17_or0;
  wire s_CSAwallace_rca16_u_rca32_fa18_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa18_and0;
  wire s_CSAwallace_rca16_u_rca32_fa18_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa18_and1;
  wire s_CSAwallace_rca16_u_rca32_fa18_or0;
  wire s_CSAwallace_rca16_u_rca32_fa19_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa19_and0;
  wire s_CSAwallace_rca16_u_rca32_fa19_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa19_and1;
  wire s_CSAwallace_rca16_u_rca32_fa19_or0;
  wire s_CSAwallace_rca16_u_rca32_fa20_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa20_and0;
  wire s_CSAwallace_rca16_u_rca32_fa20_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa20_and1;
  wire s_CSAwallace_rca16_u_rca32_fa20_or0;
  wire s_CSAwallace_rca16_u_rca32_fa21_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa21_and0;
  wire s_CSAwallace_rca16_u_rca32_fa21_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa21_and1;
  wire s_CSAwallace_rca16_u_rca32_fa21_or0;
  wire s_CSAwallace_rca16_u_rca32_fa22_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa22_and0;
  wire s_CSAwallace_rca16_u_rca32_fa22_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa22_and1;
  wire s_CSAwallace_rca16_u_rca32_fa22_or0;
  wire s_CSAwallace_rca16_u_rca32_fa23_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa23_and0;
  wire s_CSAwallace_rca16_u_rca32_fa23_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa23_and1;
  wire s_CSAwallace_rca16_u_rca32_fa23_or0;
  wire s_CSAwallace_rca16_u_rca32_fa24_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa24_and0;
  wire s_CSAwallace_rca16_u_rca32_fa24_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa24_and1;
  wire s_CSAwallace_rca16_u_rca32_fa24_or0;
  wire s_CSAwallace_rca16_u_rca32_fa25_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa25_and0;
  wire s_CSAwallace_rca16_u_rca32_fa25_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa25_and1;
  wire s_CSAwallace_rca16_u_rca32_fa25_or0;
  wire s_CSAwallace_rca16_u_rca32_fa26_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa26_and0;
  wire s_CSAwallace_rca16_u_rca32_fa26_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa26_and1;
  wire s_CSAwallace_rca16_u_rca32_fa26_or0;
  wire s_CSAwallace_rca16_u_rca32_fa27_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa27_and0;
  wire s_CSAwallace_rca16_u_rca32_fa27_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa27_and1;
  wire s_CSAwallace_rca16_u_rca32_fa27_or0;
  wire s_CSAwallace_rca16_u_rca32_fa28_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa28_and0;
  wire s_CSAwallace_rca16_u_rca32_fa28_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa28_and1;
  wire s_CSAwallace_rca16_u_rca32_fa28_or0;
  wire s_CSAwallace_rca16_u_rca32_fa29_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa29_and0;
  wire s_CSAwallace_rca16_u_rca32_fa29_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa29_and1;
  wire s_CSAwallace_rca16_u_rca32_fa29_or0;
  wire s_CSAwallace_rca16_u_rca32_fa30_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa30_and0;
  wire s_CSAwallace_rca16_u_rca32_fa30_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa30_and1;
  wire s_CSAwallace_rca16_u_rca32_fa30_or0;
  wire s_CSAwallace_rca16_u_rca32_fa31_xor0;
  wire s_CSAwallace_rca16_u_rca32_fa31_and0;
  wire s_CSAwallace_rca16_u_rca32_fa31_xor1;
  wire s_CSAwallace_rca16_u_rca32_fa31_and1;
  wire s_CSAwallace_rca16_u_rca32_fa31_or0;
  wire s_CSAwallace_rca16_xor0;

  assign s_CSAwallace_rca16_and_0_0 = a[0] & b[0];
  assign s_CSAwallace_rca16_and_1_0 = a[1] & b[0];
  assign s_CSAwallace_rca16_and_2_0 = a[2] & b[0];
  assign s_CSAwallace_rca16_and_3_0 = a[3] & b[0];
  assign s_CSAwallace_rca16_and_4_0 = a[4] & b[0];
  assign s_CSAwallace_rca16_and_5_0 = a[5] & b[0];
  assign s_CSAwallace_rca16_and_6_0 = a[6] & b[0];
  assign s_CSAwallace_rca16_and_7_0 = a[7] & b[0];
  assign s_CSAwallace_rca16_and_8_0 = a[8] & b[0];
  assign s_CSAwallace_rca16_and_9_0 = a[9] & b[0];
  assign s_CSAwallace_rca16_and_10_0 = a[10] & b[0];
  assign s_CSAwallace_rca16_and_11_0 = a[11] & b[0];
  assign s_CSAwallace_rca16_and_12_0 = a[12] & b[0];
  assign s_CSAwallace_rca16_and_13_0 = a[13] & b[0];
  assign s_CSAwallace_rca16_and_14_0 = a[14] & b[0];
  assign s_CSAwallace_rca16_nand_15_0 = ~(a[15] & b[0]);
  assign s_CSAwallace_rca16_and_0_1 = a[0] & b[1];
  assign s_CSAwallace_rca16_and_1_1 = a[1] & b[1];
  assign s_CSAwallace_rca16_and_2_1 = a[2] & b[1];
  assign s_CSAwallace_rca16_and_3_1 = a[3] & b[1];
  assign s_CSAwallace_rca16_and_4_1 = a[4] & b[1];
  assign s_CSAwallace_rca16_and_5_1 = a[5] & b[1];
  assign s_CSAwallace_rca16_and_6_1 = a[6] & b[1];
  assign s_CSAwallace_rca16_and_7_1 = a[7] & b[1];
  assign s_CSAwallace_rca16_and_8_1 = a[8] & b[1];
  assign s_CSAwallace_rca16_and_9_1 = a[9] & b[1];
  assign s_CSAwallace_rca16_and_10_1 = a[10] & b[1];
  assign s_CSAwallace_rca16_and_11_1 = a[11] & b[1];
  assign s_CSAwallace_rca16_and_12_1 = a[12] & b[1];
  assign s_CSAwallace_rca16_and_13_1 = a[13] & b[1];
  assign s_CSAwallace_rca16_and_14_1 = a[14] & b[1];
  assign s_CSAwallace_rca16_nand_15_1 = ~(a[15] & b[1]);
  assign s_CSAwallace_rca16_and_0_2 = a[0] & b[2];
  assign s_CSAwallace_rca16_and_1_2 = a[1] & b[2];
  assign s_CSAwallace_rca16_and_2_2 = a[2] & b[2];
  assign s_CSAwallace_rca16_and_3_2 = a[3] & b[2];
  assign s_CSAwallace_rca16_and_4_2 = a[4] & b[2];
  assign s_CSAwallace_rca16_and_5_2 = a[5] & b[2];
  assign s_CSAwallace_rca16_and_6_2 = a[6] & b[2];
  assign s_CSAwallace_rca16_and_7_2 = a[7] & b[2];
  assign s_CSAwallace_rca16_and_8_2 = a[8] & b[2];
  assign s_CSAwallace_rca16_and_9_2 = a[9] & b[2];
  assign s_CSAwallace_rca16_and_10_2 = a[10] & b[2];
  assign s_CSAwallace_rca16_and_11_2 = a[11] & b[2];
  assign s_CSAwallace_rca16_and_12_2 = a[12] & b[2];
  assign s_CSAwallace_rca16_and_13_2 = a[13] & b[2];
  assign s_CSAwallace_rca16_and_14_2 = a[14] & b[2];
  assign s_CSAwallace_rca16_nand_15_2 = ~(a[15] & b[2]);
  assign s_CSAwallace_rca16_and_0_3 = a[0] & b[3];
  assign s_CSAwallace_rca16_and_1_3 = a[1] & b[3];
  assign s_CSAwallace_rca16_and_2_3 = a[2] & b[3];
  assign s_CSAwallace_rca16_and_3_3 = a[3] & b[3];
  assign s_CSAwallace_rca16_and_4_3 = a[4] & b[3];
  assign s_CSAwallace_rca16_and_5_3 = a[5] & b[3];
  assign s_CSAwallace_rca16_and_6_3 = a[6] & b[3];
  assign s_CSAwallace_rca16_and_7_3 = a[7] & b[3];
  assign s_CSAwallace_rca16_and_8_3 = a[8] & b[3];
  assign s_CSAwallace_rca16_and_9_3 = a[9] & b[3];
  assign s_CSAwallace_rca16_and_10_3 = a[10] & b[3];
  assign s_CSAwallace_rca16_and_11_3 = a[11] & b[3];
  assign s_CSAwallace_rca16_and_12_3 = a[12] & b[3];
  assign s_CSAwallace_rca16_and_13_3 = a[13] & b[3];
  assign s_CSAwallace_rca16_and_14_3 = a[14] & b[3];
  assign s_CSAwallace_rca16_nand_15_3 = ~(a[15] & b[3]);
  assign s_CSAwallace_rca16_and_0_4 = a[0] & b[4];
  assign s_CSAwallace_rca16_and_1_4 = a[1] & b[4];
  assign s_CSAwallace_rca16_and_2_4 = a[2] & b[4];
  assign s_CSAwallace_rca16_and_3_4 = a[3] & b[4];
  assign s_CSAwallace_rca16_and_4_4 = a[4] & b[4];
  assign s_CSAwallace_rca16_and_5_4 = a[5] & b[4];
  assign s_CSAwallace_rca16_and_6_4 = a[6] & b[4];
  assign s_CSAwallace_rca16_and_7_4 = a[7] & b[4];
  assign s_CSAwallace_rca16_and_8_4 = a[8] & b[4];
  assign s_CSAwallace_rca16_and_9_4 = a[9] & b[4];
  assign s_CSAwallace_rca16_and_10_4 = a[10] & b[4];
  assign s_CSAwallace_rca16_and_11_4 = a[11] & b[4];
  assign s_CSAwallace_rca16_and_12_4 = a[12] & b[4];
  assign s_CSAwallace_rca16_and_13_4 = a[13] & b[4];
  assign s_CSAwallace_rca16_and_14_4 = a[14] & b[4];
  assign s_CSAwallace_rca16_nand_15_4 = ~(a[15] & b[4]);
  assign s_CSAwallace_rca16_and_0_5 = a[0] & b[5];
  assign s_CSAwallace_rca16_and_1_5 = a[1] & b[5];
  assign s_CSAwallace_rca16_and_2_5 = a[2] & b[5];
  assign s_CSAwallace_rca16_and_3_5 = a[3] & b[5];
  assign s_CSAwallace_rca16_and_4_5 = a[4] & b[5];
  assign s_CSAwallace_rca16_and_5_5 = a[5] & b[5];
  assign s_CSAwallace_rca16_and_6_5 = a[6] & b[5];
  assign s_CSAwallace_rca16_and_7_5 = a[7] & b[5];
  assign s_CSAwallace_rca16_and_8_5 = a[8] & b[5];
  assign s_CSAwallace_rca16_and_9_5 = a[9] & b[5];
  assign s_CSAwallace_rca16_and_10_5 = a[10] & b[5];
  assign s_CSAwallace_rca16_and_11_5 = a[11] & b[5];
  assign s_CSAwallace_rca16_and_12_5 = a[12] & b[5];
  assign s_CSAwallace_rca16_and_13_5 = a[13] & b[5];
  assign s_CSAwallace_rca16_and_14_5 = a[14] & b[5];
  assign s_CSAwallace_rca16_nand_15_5 = ~(a[15] & b[5]);
  assign s_CSAwallace_rca16_and_0_6 = a[0] & b[6];
  assign s_CSAwallace_rca16_and_1_6 = a[1] & b[6];
  assign s_CSAwallace_rca16_and_2_6 = a[2] & b[6];
  assign s_CSAwallace_rca16_and_3_6 = a[3] & b[6];
  assign s_CSAwallace_rca16_and_4_6 = a[4] & b[6];
  assign s_CSAwallace_rca16_and_5_6 = a[5] & b[6];
  assign s_CSAwallace_rca16_and_6_6 = a[6] & b[6];
  assign s_CSAwallace_rca16_and_7_6 = a[7] & b[6];
  assign s_CSAwallace_rca16_and_8_6 = a[8] & b[6];
  assign s_CSAwallace_rca16_and_9_6 = a[9] & b[6];
  assign s_CSAwallace_rca16_and_10_6 = a[10] & b[6];
  assign s_CSAwallace_rca16_and_11_6 = a[11] & b[6];
  assign s_CSAwallace_rca16_and_12_6 = a[12] & b[6];
  assign s_CSAwallace_rca16_and_13_6 = a[13] & b[6];
  assign s_CSAwallace_rca16_and_14_6 = a[14] & b[6];
  assign s_CSAwallace_rca16_nand_15_6 = ~(a[15] & b[6]);
  assign s_CSAwallace_rca16_and_0_7 = a[0] & b[7];
  assign s_CSAwallace_rca16_and_1_7 = a[1] & b[7];
  assign s_CSAwallace_rca16_and_2_7 = a[2] & b[7];
  assign s_CSAwallace_rca16_and_3_7 = a[3] & b[7];
  assign s_CSAwallace_rca16_and_4_7 = a[4] & b[7];
  assign s_CSAwallace_rca16_and_5_7 = a[5] & b[7];
  assign s_CSAwallace_rca16_and_6_7 = a[6] & b[7];
  assign s_CSAwallace_rca16_and_7_7 = a[7] & b[7];
  assign s_CSAwallace_rca16_and_8_7 = a[8] & b[7];
  assign s_CSAwallace_rca16_and_9_7 = a[9] & b[7];
  assign s_CSAwallace_rca16_and_10_7 = a[10] & b[7];
  assign s_CSAwallace_rca16_and_11_7 = a[11] & b[7];
  assign s_CSAwallace_rca16_and_12_7 = a[12] & b[7];
  assign s_CSAwallace_rca16_and_13_7 = a[13] & b[7];
  assign s_CSAwallace_rca16_and_14_7 = a[14] & b[7];
  assign s_CSAwallace_rca16_nand_15_7 = ~(a[15] & b[7]);
  assign s_CSAwallace_rca16_and_0_8 = a[0] & b[8];
  assign s_CSAwallace_rca16_and_1_8 = a[1] & b[8];
  assign s_CSAwallace_rca16_and_2_8 = a[2] & b[8];
  assign s_CSAwallace_rca16_and_3_8 = a[3] & b[8];
  assign s_CSAwallace_rca16_and_4_8 = a[4] & b[8];
  assign s_CSAwallace_rca16_and_5_8 = a[5] & b[8];
  assign s_CSAwallace_rca16_and_6_8 = a[6] & b[8];
  assign s_CSAwallace_rca16_and_7_8 = a[7] & b[8];
  assign s_CSAwallace_rca16_and_8_8 = a[8] & b[8];
  assign s_CSAwallace_rca16_and_9_8 = a[9] & b[8];
  assign s_CSAwallace_rca16_and_10_8 = a[10] & b[8];
  assign s_CSAwallace_rca16_and_11_8 = a[11] & b[8];
  assign s_CSAwallace_rca16_and_12_8 = a[12] & b[8];
  assign s_CSAwallace_rca16_and_13_8 = a[13] & b[8];
  assign s_CSAwallace_rca16_and_14_8 = a[14] & b[8];
  assign s_CSAwallace_rca16_nand_15_8 = ~(a[15] & b[8]);
  assign s_CSAwallace_rca16_and_0_9 = a[0] & b[9];
  assign s_CSAwallace_rca16_and_1_9 = a[1] & b[9];
  assign s_CSAwallace_rca16_and_2_9 = a[2] & b[9];
  assign s_CSAwallace_rca16_and_3_9 = a[3] & b[9];
  assign s_CSAwallace_rca16_and_4_9 = a[4] & b[9];
  assign s_CSAwallace_rca16_and_5_9 = a[5] & b[9];
  assign s_CSAwallace_rca16_and_6_9 = a[6] & b[9];
  assign s_CSAwallace_rca16_and_7_9 = a[7] & b[9];
  assign s_CSAwallace_rca16_and_8_9 = a[8] & b[9];
  assign s_CSAwallace_rca16_and_9_9 = a[9] & b[9];
  assign s_CSAwallace_rca16_and_10_9 = a[10] & b[9];
  assign s_CSAwallace_rca16_and_11_9 = a[11] & b[9];
  assign s_CSAwallace_rca16_and_12_9 = a[12] & b[9];
  assign s_CSAwallace_rca16_and_13_9 = a[13] & b[9];
  assign s_CSAwallace_rca16_and_14_9 = a[14] & b[9];
  assign s_CSAwallace_rca16_nand_15_9 = ~(a[15] & b[9]);
  assign s_CSAwallace_rca16_and_0_10 = a[0] & b[10];
  assign s_CSAwallace_rca16_and_1_10 = a[1] & b[10];
  assign s_CSAwallace_rca16_and_2_10 = a[2] & b[10];
  assign s_CSAwallace_rca16_and_3_10 = a[3] & b[10];
  assign s_CSAwallace_rca16_and_4_10 = a[4] & b[10];
  assign s_CSAwallace_rca16_and_5_10 = a[5] & b[10];
  assign s_CSAwallace_rca16_and_6_10 = a[6] & b[10];
  assign s_CSAwallace_rca16_and_7_10 = a[7] & b[10];
  assign s_CSAwallace_rca16_and_8_10 = a[8] & b[10];
  assign s_CSAwallace_rca16_and_9_10 = a[9] & b[10];
  assign s_CSAwallace_rca16_and_10_10 = a[10] & b[10];
  assign s_CSAwallace_rca16_and_11_10 = a[11] & b[10];
  assign s_CSAwallace_rca16_and_12_10 = a[12] & b[10];
  assign s_CSAwallace_rca16_and_13_10 = a[13] & b[10];
  assign s_CSAwallace_rca16_and_14_10 = a[14] & b[10];
  assign s_CSAwallace_rca16_nand_15_10 = ~(a[15] & b[10]);
  assign s_CSAwallace_rca16_and_0_11 = a[0] & b[11];
  assign s_CSAwallace_rca16_and_1_11 = a[1] & b[11];
  assign s_CSAwallace_rca16_and_2_11 = a[2] & b[11];
  assign s_CSAwallace_rca16_and_3_11 = a[3] & b[11];
  assign s_CSAwallace_rca16_and_4_11 = a[4] & b[11];
  assign s_CSAwallace_rca16_and_5_11 = a[5] & b[11];
  assign s_CSAwallace_rca16_and_6_11 = a[6] & b[11];
  assign s_CSAwallace_rca16_and_7_11 = a[7] & b[11];
  assign s_CSAwallace_rca16_and_8_11 = a[8] & b[11];
  assign s_CSAwallace_rca16_and_9_11 = a[9] & b[11];
  assign s_CSAwallace_rca16_and_10_11 = a[10] & b[11];
  assign s_CSAwallace_rca16_and_11_11 = a[11] & b[11];
  assign s_CSAwallace_rca16_and_12_11 = a[12] & b[11];
  assign s_CSAwallace_rca16_and_13_11 = a[13] & b[11];
  assign s_CSAwallace_rca16_and_14_11 = a[14] & b[11];
  assign s_CSAwallace_rca16_nand_15_11 = ~(a[15] & b[11]);
  assign s_CSAwallace_rca16_and_0_12 = a[0] & b[12];
  assign s_CSAwallace_rca16_and_1_12 = a[1] & b[12];
  assign s_CSAwallace_rca16_and_2_12 = a[2] & b[12];
  assign s_CSAwallace_rca16_and_3_12 = a[3] & b[12];
  assign s_CSAwallace_rca16_and_4_12 = a[4] & b[12];
  assign s_CSAwallace_rca16_and_5_12 = a[5] & b[12];
  assign s_CSAwallace_rca16_and_6_12 = a[6] & b[12];
  assign s_CSAwallace_rca16_and_7_12 = a[7] & b[12];
  assign s_CSAwallace_rca16_and_8_12 = a[8] & b[12];
  assign s_CSAwallace_rca16_and_9_12 = a[9] & b[12];
  assign s_CSAwallace_rca16_and_10_12 = a[10] & b[12];
  assign s_CSAwallace_rca16_and_11_12 = a[11] & b[12];
  assign s_CSAwallace_rca16_and_12_12 = a[12] & b[12];
  assign s_CSAwallace_rca16_and_13_12 = a[13] & b[12];
  assign s_CSAwallace_rca16_and_14_12 = a[14] & b[12];
  assign s_CSAwallace_rca16_nand_15_12 = ~(a[15] & b[12]);
  assign s_CSAwallace_rca16_and_0_13 = a[0] & b[13];
  assign s_CSAwallace_rca16_and_1_13 = a[1] & b[13];
  assign s_CSAwallace_rca16_and_2_13 = a[2] & b[13];
  assign s_CSAwallace_rca16_and_3_13 = a[3] & b[13];
  assign s_CSAwallace_rca16_and_4_13 = a[4] & b[13];
  assign s_CSAwallace_rca16_and_5_13 = a[5] & b[13];
  assign s_CSAwallace_rca16_and_6_13 = a[6] & b[13];
  assign s_CSAwallace_rca16_and_7_13 = a[7] & b[13];
  assign s_CSAwallace_rca16_and_8_13 = a[8] & b[13];
  assign s_CSAwallace_rca16_and_9_13 = a[9] & b[13];
  assign s_CSAwallace_rca16_and_10_13 = a[10] & b[13];
  assign s_CSAwallace_rca16_and_11_13 = a[11] & b[13];
  assign s_CSAwallace_rca16_and_12_13 = a[12] & b[13];
  assign s_CSAwallace_rca16_and_13_13 = a[13] & b[13];
  assign s_CSAwallace_rca16_and_14_13 = a[14] & b[13];
  assign s_CSAwallace_rca16_nand_15_13 = ~(a[15] & b[13]);
  assign s_CSAwallace_rca16_and_0_14 = a[0] & b[14];
  assign s_CSAwallace_rca16_and_1_14 = a[1] & b[14];
  assign s_CSAwallace_rca16_and_2_14 = a[2] & b[14];
  assign s_CSAwallace_rca16_and_3_14 = a[3] & b[14];
  assign s_CSAwallace_rca16_and_4_14 = a[4] & b[14];
  assign s_CSAwallace_rca16_and_5_14 = a[5] & b[14];
  assign s_CSAwallace_rca16_and_6_14 = a[6] & b[14];
  assign s_CSAwallace_rca16_and_7_14 = a[7] & b[14];
  assign s_CSAwallace_rca16_and_8_14 = a[8] & b[14];
  assign s_CSAwallace_rca16_and_9_14 = a[9] & b[14];
  assign s_CSAwallace_rca16_and_10_14 = a[10] & b[14];
  assign s_CSAwallace_rca16_and_11_14 = a[11] & b[14];
  assign s_CSAwallace_rca16_and_12_14 = a[12] & b[14];
  assign s_CSAwallace_rca16_and_13_14 = a[13] & b[14];
  assign s_CSAwallace_rca16_and_14_14 = a[14] & b[14];
  assign s_CSAwallace_rca16_nand_15_14 = ~(a[15] & b[14]);
  assign s_CSAwallace_rca16_nand_0_15 = ~(a[0] & b[15]);
  assign s_CSAwallace_rca16_nand_1_15 = ~(a[1] & b[15]);
  assign s_CSAwallace_rca16_nand_2_15 = ~(a[2] & b[15]);
  assign s_CSAwallace_rca16_nand_3_15 = ~(a[3] & b[15]);
  assign s_CSAwallace_rca16_nand_4_15 = ~(a[4] & b[15]);
  assign s_CSAwallace_rca16_nand_5_15 = ~(a[5] & b[15]);
  assign s_CSAwallace_rca16_nand_6_15 = ~(a[6] & b[15]);
  assign s_CSAwallace_rca16_nand_7_15 = ~(a[7] & b[15]);
  assign s_CSAwallace_rca16_nand_8_15 = ~(a[8] & b[15]);
  assign s_CSAwallace_rca16_nand_9_15 = ~(a[9] & b[15]);
  assign s_CSAwallace_rca16_nand_10_15 = ~(a[10] & b[15]);
  assign s_CSAwallace_rca16_nand_11_15 = ~(a[11] & b[15]);
  assign s_CSAwallace_rca16_nand_12_15 = ~(a[12] & b[15]);
  assign s_CSAwallace_rca16_nand_13_15 = ~(a[13] & b[15]);
  assign s_CSAwallace_rca16_nand_14_15 = ~(a[14] & b[15]);
  assign s_CSAwallace_rca16_and_15_15 = a[15] & b[15];
  assign s_CSAwallace_rca16_csa0_csa_component_fa1_xor0 = s_CSAwallace_rca16_and_1_0 ^ s_CSAwallace_rca16_and_0_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa1_and0 = s_CSAwallace_rca16_and_1_0 & s_CSAwallace_rca16_and_0_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa2_xor0 = s_CSAwallace_rca16_and_2_0 ^ s_CSAwallace_rca16_and_1_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa2_and0 = s_CSAwallace_rca16_and_2_0 & s_CSAwallace_rca16_and_1_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa2_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa2_xor0 ^ s_CSAwallace_rca16_and_0_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa2_and1 = s_CSAwallace_rca16_csa0_csa_component_fa2_xor0 & s_CSAwallace_rca16_and_0_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa2_or0 = s_CSAwallace_rca16_csa0_csa_component_fa2_and0 | s_CSAwallace_rca16_csa0_csa_component_fa2_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa3_xor0 = s_CSAwallace_rca16_and_3_0 ^ s_CSAwallace_rca16_and_2_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa3_and0 = s_CSAwallace_rca16_and_3_0 & s_CSAwallace_rca16_and_2_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa3_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa3_xor0 ^ s_CSAwallace_rca16_and_1_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa3_and1 = s_CSAwallace_rca16_csa0_csa_component_fa3_xor0 & s_CSAwallace_rca16_and_1_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa3_or0 = s_CSAwallace_rca16_csa0_csa_component_fa3_and0 | s_CSAwallace_rca16_csa0_csa_component_fa3_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa4_xor0 = s_CSAwallace_rca16_and_4_0 ^ s_CSAwallace_rca16_and_3_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa4_and0 = s_CSAwallace_rca16_and_4_0 & s_CSAwallace_rca16_and_3_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa4_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa4_xor0 ^ s_CSAwallace_rca16_and_2_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa4_and1 = s_CSAwallace_rca16_csa0_csa_component_fa4_xor0 & s_CSAwallace_rca16_and_2_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa4_or0 = s_CSAwallace_rca16_csa0_csa_component_fa4_and0 | s_CSAwallace_rca16_csa0_csa_component_fa4_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa5_xor0 = s_CSAwallace_rca16_and_5_0 ^ s_CSAwallace_rca16_and_4_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa5_and0 = s_CSAwallace_rca16_and_5_0 & s_CSAwallace_rca16_and_4_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa5_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa5_xor0 ^ s_CSAwallace_rca16_and_3_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa5_and1 = s_CSAwallace_rca16_csa0_csa_component_fa5_xor0 & s_CSAwallace_rca16_and_3_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa5_or0 = s_CSAwallace_rca16_csa0_csa_component_fa5_and0 | s_CSAwallace_rca16_csa0_csa_component_fa5_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa6_xor0 = s_CSAwallace_rca16_and_6_0 ^ s_CSAwallace_rca16_and_5_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa6_and0 = s_CSAwallace_rca16_and_6_0 & s_CSAwallace_rca16_and_5_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa6_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa6_xor0 ^ s_CSAwallace_rca16_and_4_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa6_and1 = s_CSAwallace_rca16_csa0_csa_component_fa6_xor0 & s_CSAwallace_rca16_and_4_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa6_or0 = s_CSAwallace_rca16_csa0_csa_component_fa6_and0 | s_CSAwallace_rca16_csa0_csa_component_fa6_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa7_xor0 = s_CSAwallace_rca16_and_7_0 ^ s_CSAwallace_rca16_and_6_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa7_and0 = s_CSAwallace_rca16_and_7_0 & s_CSAwallace_rca16_and_6_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa7_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa7_xor0 ^ s_CSAwallace_rca16_and_5_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa7_and1 = s_CSAwallace_rca16_csa0_csa_component_fa7_xor0 & s_CSAwallace_rca16_and_5_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa7_or0 = s_CSAwallace_rca16_csa0_csa_component_fa7_and0 | s_CSAwallace_rca16_csa0_csa_component_fa7_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa8_xor0 = s_CSAwallace_rca16_and_8_0 ^ s_CSAwallace_rca16_and_7_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa8_and0 = s_CSAwallace_rca16_and_8_0 & s_CSAwallace_rca16_and_7_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa8_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa8_xor0 ^ s_CSAwallace_rca16_and_6_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa8_and1 = s_CSAwallace_rca16_csa0_csa_component_fa8_xor0 & s_CSAwallace_rca16_and_6_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa8_or0 = s_CSAwallace_rca16_csa0_csa_component_fa8_and0 | s_CSAwallace_rca16_csa0_csa_component_fa8_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa9_xor0 = s_CSAwallace_rca16_and_9_0 ^ s_CSAwallace_rca16_and_8_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa9_and0 = s_CSAwallace_rca16_and_9_0 & s_CSAwallace_rca16_and_8_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa9_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa9_xor0 ^ s_CSAwallace_rca16_and_7_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa9_and1 = s_CSAwallace_rca16_csa0_csa_component_fa9_xor0 & s_CSAwallace_rca16_and_7_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa9_or0 = s_CSAwallace_rca16_csa0_csa_component_fa9_and0 | s_CSAwallace_rca16_csa0_csa_component_fa9_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa10_xor0 = s_CSAwallace_rca16_and_10_0 ^ s_CSAwallace_rca16_and_9_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa10_and0 = s_CSAwallace_rca16_and_10_0 & s_CSAwallace_rca16_and_9_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa10_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa10_xor0 ^ s_CSAwallace_rca16_and_8_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa10_and1 = s_CSAwallace_rca16_csa0_csa_component_fa10_xor0 & s_CSAwallace_rca16_and_8_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa10_or0 = s_CSAwallace_rca16_csa0_csa_component_fa10_and0 | s_CSAwallace_rca16_csa0_csa_component_fa10_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa11_xor0 = s_CSAwallace_rca16_and_11_0 ^ s_CSAwallace_rca16_and_10_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa11_and0 = s_CSAwallace_rca16_and_11_0 & s_CSAwallace_rca16_and_10_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa11_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_and_9_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa11_and1 = s_CSAwallace_rca16_csa0_csa_component_fa11_xor0 & s_CSAwallace_rca16_and_9_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa11_or0 = s_CSAwallace_rca16_csa0_csa_component_fa11_and0 | s_CSAwallace_rca16_csa0_csa_component_fa11_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa12_xor0 = s_CSAwallace_rca16_and_12_0 ^ s_CSAwallace_rca16_and_11_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa12_and0 = s_CSAwallace_rca16_and_12_0 & s_CSAwallace_rca16_and_11_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_and_10_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa12_and1 = s_CSAwallace_rca16_csa0_csa_component_fa12_xor0 & s_CSAwallace_rca16_and_10_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa12_or0 = s_CSAwallace_rca16_csa0_csa_component_fa12_and0 | s_CSAwallace_rca16_csa0_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa13_xor0 = s_CSAwallace_rca16_and_13_0 ^ s_CSAwallace_rca16_and_12_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa13_and0 = s_CSAwallace_rca16_and_13_0 & s_CSAwallace_rca16_and_12_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_and_11_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa13_and1 = s_CSAwallace_rca16_csa0_csa_component_fa13_xor0 & s_CSAwallace_rca16_and_11_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa13_or0 = s_CSAwallace_rca16_csa0_csa_component_fa13_and0 | s_CSAwallace_rca16_csa0_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa14_xor0 = s_CSAwallace_rca16_and_14_0 ^ s_CSAwallace_rca16_and_13_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa14_and0 = s_CSAwallace_rca16_and_14_0 & s_CSAwallace_rca16_and_13_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_and_12_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa14_and1 = s_CSAwallace_rca16_csa0_csa_component_fa14_xor0 & s_CSAwallace_rca16_and_12_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa14_or0 = s_CSAwallace_rca16_csa0_csa_component_fa14_and0 | s_CSAwallace_rca16_csa0_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa15_xor0 = s_CSAwallace_rca16_nand_15_0 ^ s_CSAwallace_rca16_and_14_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa15_and0 = s_CSAwallace_rca16_nand_15_0 & s_CSAwallace_rca16_and_14_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_and_13_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa15_and1 = s_CSAwallace_rca16_csa0_csa_component_fa15_xor0 & s_CSAwallace_rca16_and_13_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa15_or0 = s_CSAwallace_rca16_csa0_csa_component_fa15_and0 | s_CSAwallace_rca16_csa0_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa16_xor0 = ~s_CSAwallace_rca16_nand_15_1;
  assign s_CSAwallace_rca16_csa0_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa0_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_and_14_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa16_and1 = s_CSAwallace_rca16_csa0_csa_component_fa16_xor0 & s_CSAwallace_rca16_and_14_2;
  assign s_CSAwallace_rca16_csa0_csa_component_fa16_or0 = s_CSAwallace_rca16_nand_15_1 | s_CSAwallace_rca16_csa0_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa4_xor0 = s_CSAwallace_rca16_and_1_3 ^ s_CSAwallace_rca16_and_0_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa4_and0 = s_CSAwallace_rca16_and_1_3 & s_CSAwallace_rca16_and_0_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa5_xor0 = s_CSAwallace_rca16_and_2_3 ^ s_CSAwallace_rca16_and_1_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa5_and0 = s_CSAwallace_rca16_and_2_3 & s_CSAwallace_rca16_and_1_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa5_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa5_xor0 ^ s_CSAwallace_rca16_and_0_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa5_and1 = s_CSAwallace_rca16_csa1_csa_component_fa5_xor0 & s_CSAwallace_rca16_and_0_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa5_or0 = s_CSAwallace_rca16_csa1_csa_component_fa5_and0 | s_CSAwallace_rca16_csa1_csa_component_fa5_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa6_xor0 = s_CSAwallace_rca16_and_3_3 ^ s_CSAwallace_rca16_and_2_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa6_and0 = s_CSAwallace_rca16_and_3_3 & s_CSAwallace_rca16_and_2_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa6_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa6_xor0 ^ s_CSAwallace_rca16_and_1_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa6_and1 = s_CSAwallace_rca16_csa1_csa_component_fa6_xor0 & s_CSAwallace_rca16_and_1_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa6_or0 = s_CSAwallace_rca16_csa1_csa_component_fa6_and0 | s_CSAwallace_rca16_csa1_csa_component_fa6_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa7_xor0 = s_CSAwallace_rca16_and_4_3 ^ s_CSAwallace_rca16_and_3_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa7_and0 = s_CSAwallace_rca16_and_4_3 & s_CSAwallace_rca16_and_3_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa7_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa7_xor0 ^ s_CSAwallace_rca16_and_2_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa7_and1 = s_CSAwallace_rca16_csa1_csa_component_fa7_xor0 & s_CSAwallace_rca16_and_2_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa7_or0 = s_CSAwallace_rca16_csa1_csa_component_fa7_and0 | s_CSAwallace_rca16_csa1_csa_component_fa7_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa8_xor0 = s_CSAwallace_rca16_and_5_3 ^ s_CSAwallace_rca16_and_4_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa8_and0 = s_CSAwallace_rca16_and_5_3 & s_CSAwallace_rca16_and_4_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa8_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa8_xor0 ^ s_CSAwallace_rca16_and_3_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa8_and1 = s_CSAwallace_rca16_csa1_csa_component_fa8_xor0 & s_CSAwallace_rca16_and_3_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa8_or0 = s_CSAwallace_rca16_csa1_csa_component_fa8_and0 | s_CSAwallace_rca16_csa1_csa_component_fa8_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa9_xor0 = s_CSAwallace_rca16_and_6_3 ^ s_CSAwallace_rca16_and_5_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa9_and0 = s_CSAwallace_rca16_and_6_3 & s_CSAwallace_rca16_and_5_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa9_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa9_xor0 ^ s_CSAwallace_rca16_and_4_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa9_and1 = s_CSAwallace_rca16_csa1_csa_component_fa9_xor0 & s_CSAwallace_rca16_and_4_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa9_or0 = s_CSAwallace_rca16_csa1_csa_component_fa9_and0 | s_CSAwallace_rca16_csa1_csa_component_fa9_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa10_xor0 = s_CSAwallace_rca16_and_7_3 ^ s_CSAwallace_rca16_and_6_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa10_and0 = s_CSAwallace_rca16_and_7_3 & s_CSAwallace_rca16_and_6_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa10_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa10_xor0 ^ s_CSAwallace_rca16_and_5_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa10_and1 = s_CSAwallace_rca16_csa1_csa_component_fa10_xor0 & s_CSAwallace_rca16_and_5_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa10_or0 = s_CSAwallace_rca16_csa1_csa_component_fa10_and0 | s_CSAwallace_rca16_csa1_csa_component_fa10_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa11_xor0 = s_CSAwallace_rca16_and_8_3 ^ s_CSAwallace_rca16_and_7_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa11_and0 = s_CSAwallace_rca16_and_8_3 & s_CSAwallace_rca16_and_7_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa11_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_and_6_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa11_and1 = s_CSAwallace_rca16_csa1_csa_component_fa11_xor0 & s_CSAwallace_rca16_and_6_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa11_or0 = s_CSAwallace_rca16_csa1_csa_component_fa11_and0 | s_CSAwallace_rca16_csa1_csa_component_fa11_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa12_xor0 = s_CSAwallace_rca16_and_9_3 ^ s_CSAwallace_rca16_and_8_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa12_and0 = s_CSAwallace_rca16_and_9_3 & s_CSAwallace_rca16_and_8_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_and_7_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa12_and1 = s_CSAwallace_rca16_csa1_csa_component_fa12_xor0 & s_CSAwallace_rca16_and_7_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa12_or0 = s_CSAwallace_rca16_csa1_csa_component_fa12_and0 | s_CSAwallace_rca16_csa1_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa13_xor0 = s_CSAwallace_rca16_and_10_3 ^ s_CSAwallace_rca16_and_9_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa13_and0 = s_CSAwallace_rca16_and_10_3 & s_CSAwallace_rca16_and_9_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_and_8_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa13_and1 = s_CSAwallace_rca16_csa1_csa_component_fa13_xor0 & s_CSAwallace_rca16_and_8_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa13_or0 = s_CSAwallace_rca16_csa1_csa_component_fa13_and0 | s_CSAwallace_rca16_csa1_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa14_xor0 = s_CSAwallace_rca16_and_11_3 ^ s_CSAwallace_rca16_and_10_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa14_and0 = s_CSAwallace_rca16_and_11_3 & s_CSAwallace_rca16_and_10_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_and_9_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa14_and1 = s_CSAwallace_rca16_csa1_csa_component_fa14_xor0 & s_CSAwallace_rca16_and_9_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa14_or0 = s_CSAwallace_rca16_csa1_csa_component_fa14_and0 | s_CSAwallace_rca16_csa1_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa15_xor0 = s_CSAwallace_rca16_and_12_3 ^ s_CSAwallace_rca16_and_11_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa15_and0 = s_CSAwallace_rca16_and_12_3 & s_CSAwallace_rca16_and_11_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_and_10_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa15_and1 = s_CSAwallace_rca16_csa1_csa_component_fa15_xor0 & s_CSAwallace_rca16_and_10_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa15_or0 = s_CSAwallace_rca16_csa1_csa_component_fa15_and0 | s_CSAwallace_rca16_csa1_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa16_xor0 = s_CSAwallace_rca16_and_13_3 ^ s_CSAwallace_rca16_and_12_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa16_and0 = s_CSAwallace_rca16_and_13_3 & s_CSAwallace_rca16_and_12_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_and_11_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa16_and1 = s_CSAwallace_rca16_csa1_csa_component_fa16_xor0 & s_CSAwallace_rca16_and_11_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa16_or0 = s_CSAwallace_rca16_csa1_csa_component_fa16_and0 | s_CSAwallace_rca16_csa1_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa17_xor0 = s_CSAwallace_rca16_and_14_3 ^ s_CSAwallace_rca16_and_13_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa17_and0 = s_CSAwallace_rca16_and_14_3 & s_CSAwallace_rca16_and_13_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_and_12_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa17_and1 = s_CSAwallace_rca16_csa1_csa_component_fa17_xor0 & s_CSAwallace_rca16_and_12_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa17_or0 = s_CSAwallace_rca16_csa1_csa_component_fa17_and0 | s_CSAwallace_rca16_csa1_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa18_xor0 = s_CSAwallace_rca16_nand_15_3 ^ s_CSAwallace_rca16_and_14_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa18_and0 = s_CSAwallace_rca16_nand_15_3 & s_CSAwallace_rca16_and_14_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_and_13_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa18_and1 = s_CSAwallace_rca16_csa1_csa_component_fa18_xor0 & s_CSAwallace_rca16_and_13_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa18_or0 = s_CSAwallace_rca16_csa1_csa_component_fa18_and0 | s_CSAwallace_rca16_csa1_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa1_csa_component_fa19_xor0 = ~s_CSAwallace_rca16_nand_15_4;
  assign s_CSAwallace_rca16_csa1_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa1_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_and_14_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa19_and1 = s_CSAwallace_rca16_csa1_csa_component_fa19_xor0 & s_CSAwallace_rca16_and_14_5;
  assign s_CSAwallace_rca16_csa1_csa_component_fa19_or0 = s_CSAwallace_rca16_nand_15_4 | s_CSAwallace_rca16_csa1_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa7_xor0 = s_CSAwallace_rca16_and_1_6 ^ s_CSAwallace_rca16_and_0_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa7_and0 = s_CSAwallace_rca16_and_1_6 & s_CSAwallace_rca16_and_0_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa8_xor0 = s_CSAwallace_rca16_and_2_6 ^ s_CSAwallace_rca16_and_1_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa8_and0 = s_CSAwallace_rca16_and_2_6 & s_CSAwallace_rca16_and_1_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa8_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa8_xor0 ^ s_CSAwallace_rca16_and_0_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa8_and1 = s_CSAwallace_rca16_csa2_csa_component_fa8_xor0 & s_CSAwallace_rca16_and_0_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa8_or0 = s_CSAwallace_rca16_csa2_csa_component_fa8_and0 | s_CSAwallace_rca16_csa2_csa_component_fa8_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa9_xor0 = s_CSAwallace_rca16_and_3_6 ^ s_CSAwallace_rca16_and_2_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa9_and0 = s_CSAwallace_rca16_and_3_6 & s_CSAwallace_rca16_and_2_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa9_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa9_xor0 ^ s_CSAwallace_rca16_and_1_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa9_and1 = s_CSAwallace_rca16_csa2_csa_component_fa9_xor0 & s_CSAwallace_rca16_and_1_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa9_or0 = s_CSAwallace_rca16_csa2_csa_component_fa9_and0 | s_CSAwallace_rca16_csa2_csa_component_fa9_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa10_xor0 = s_CSAwallace_rca16_and_4_6 ^ s_CSAwallace_rca16_and_3_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa10_and0 = s_CSAwallace_rca16_and_4_6 & s_CSAwallace_rca16_and_3_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa10_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa10_xor0 ^ s_CSAwallace_rca16_and_2_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa10_and1 = s_CSAwallace_rca16_csa2_csa_component_fa10_xor0 & s_CSAwallace_rca16_and_2_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa10_or0 = s_CSAwallace_rca16_csa2_csa_component_fa10_and0 | s_CSAwallace_rca16_csa2_csa_component_fa10_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa11_xor0 = s_CSAwallace_rca16_and_5_6 ^ s_CSAwallace_rca16_and_4_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa11_and0 = s_CSAwallace_rca16_and_5_6 & s_CSAwallace_rca16_and_4_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa11_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_and_3_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa11_and1 = s_CSAwallace_rca16_csa2_csa_component_fa11_xor0 & s_CSAwallace_rca16_and_3_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa11_or0 = s_CSAwallace_rca16_csa2_csa_component_fa11_and0 | s_CSAwallace_rca16_csa2_csa_component_fa11_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa12_xor0 = s_CSAwallace_rca16_and_6_6 ^ s_CSAwallace_rca16_and_5_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa12_and0 = s_CSAwallace_rca16_and_6_6 & s_CSAwallace_rca16_and_5_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_and_4_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa12_and1 = s_CSAwallace_rca16_csa2_csa_component_fa12_xor0 & s_CSAwallace_rca16_and_4_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa12_or0 = s_CSAwallace_rca16_csa2_csa_component_fa12_and0 | s_CSAwallace_rca16_csa2_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa13_xor0 = s_CSAwallace_rca16_and_7_6 ^ s_CSAwallace_rca16_and_6_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa13_and0 = s_CSAwallace_rca16_and_7_6 & s_CSAwallace_rca16_and_6_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_and_5_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa13_and1 = s_CSAwallace_rca16_csa2_csa_component_fa13_xor0 & s_CSAwallace_rca16_and_5_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa13_or0 = s_CSAwallace_rca16_csa2_csa_component_fa13_and0 | s_CSAwallace_rca16_csa2_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa14_xor0 = s_CSAwallace_rca16_and_8_6 ^ s_CSAwallace_rca16_and_7_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa14_and0 = s_CSAwallace_rca16_and_8_6 & s_CSAwallace_rca16_and_7_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_and_6_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa14_and1 = s_CSAwallace_rca16_csa2_csa_component_fa14_xor0 & s_CSAwallace_rca16_and_6_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa14_or0 = s_CSAwallace_rca16_csa2_csa_component_fa14_and0 | s_CSAwallace_rca16_csa2_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa15_xor0 = s_CSAwallace_rca16_and_9_6 ^ s_CSAwallace_rca16_and_8_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa15_and0 = s_CSAwallace_rca16_and_9_6 & s_CSAwallace_rca16_and_8_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_and_7_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa15_and1 = s_CSAwallace_rca16_csa2_csa_component_fa15_xor0 & s_CSAwallace_rca16_and_7_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa15_or0 = s_CSAwallace_rca16_csa2_csa_component_fa15_and0 | s_CSAwallace_rca16_csa2_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa16_xor0 = s_CSAwallace_rca16_and_10_6 ^ s_CSAwallace_rca16_and_9_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa16_and0 = s_CSAwallace_rca16_and_10_6 & s_CSAwallace_rca16_and_9_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_and_8_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa16_and1 = s_CSAwallace_rca16_csa2_csa_component_fa16_xor0 & s_CSAwallace_rca16_and_8_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa16_or0 = s_CSAwallace_rca16_csa2_csa_component_fa16_and0 | s_CSAwallace_rca16_csa2_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa17_xor0 = s_CSAwallace_rca16_and_11_6 ^ s_CSAwallace_rca16_and_10_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa17_and0 = s_CSAwallace_rca16_and_11_6 & s_CSAwallace_rca16_and_10_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_and_9_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa17_and1 = s_CSAwallace_rca16_csa2_csa_component_fa17_xor0 & s_CSAwallace_rca16_and_9_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa17_or0 = s_CSAwallace_rca16_csa2_csa_component_fa17_and0 | s_CSAwallace_rca16_csa2_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa18_xor0 = s_CSAwallace_rca16_and_12_6 ^ s_CSAwallace_rca16_and_11_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa18_and0 = s_CSAwallace_rca16_and_12_6 & s_CSAwallace_rca16_and_11_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_and_10_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa18_and1 = s_CSAwallace_rca16_csa2_csa_component_fa18_xor0 & s_CSAwallace_rca16_and_10_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa18_or0 = s_CSAwallace_rca16_csa2_csa_component_fa18_and0 | s_CSAwallace_rca16_csa2_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa19_xor0 = s_CSAwallace_rca16_and_13_6 ^ s_CSAwallace_rca16_and_12_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa19_and0 = s_CSAwallace_rca16_and_13_6 & s_CSAwallace_rca16_and_12_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_and_11_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa19_and1 = s_CSAwallace_rca16_csa2_csa_component_fa19_xor0 & s_CSAwallace_rca16_and_11_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa19_or0 = s_CSAwallace_rca16_csa2_csa_component_fa19_and0 | s_CSAwallace_rca16_csa2_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa20_xor0 = s_CSAwallace_rca16_and_14_6 ^ s_CSAwallace_rca16_and_13_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa20_and0 = s_CSAwallace_rca16_and_14_6 & s_CSAwallace_rca16_and_13_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_and_12_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa20_and1 = s_CSAwallace_rca16_csa2_csa_component_fa20_xor0 & s_CSAwallace_rca16_and_12_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa20_or0 = s_CSAwallace_rca16_csa2_csa_component_fa20_and0 | s_CSAwallace_rca16_csa2_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa21_xor0 = s_CSAwallace_rca16_nand_15_6 ^ s_CSAwallace_rca16_and_14_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa21_and0 = s_CSAwallace_rca16_nand_15_6 & s_CSAwallace_rca16_and_14_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_and_13_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa21_and1 = s_CSAwallace_rca16_csa2_csa_component_fa21_xor0 & s_CSAwallace_rca16_and_13_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa21_or0 = s_CSAwallace_rca16_csa2_csa_component_fa21_and0 | s_CSAwallace_rca16_csa2_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa2_csa_component_fa22_xor0 = ~s_CSAwallace_rca16_nand_15_7;
  assign s_CSAwallace_rca16_csa2_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa2_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_and_14_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa22_and1 = s_CSAwallace_rca16_csa2_csa_component_fa22_xor0 & s_CSAwallace_rca16_and_14_8;
  assign s_CSAwallace_rca16_csa2_csa_component_fa22_or0 = s_CSAwallace_rca16_nand_15_7 | s_CSAwallace_rca16_csa2_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa10_xor0 = s_CSAwallace_rca16_and_1_9 ^ s_CSAwallace_rca16_and_0_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa10_and0 = s_CSAwallace_rca16_and_1_9 & s_CSAwallace_rca16_and_0_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa11_xor0 = s_CSAwallace_rca16_and_2_9 ^ s_CSAwallace_rca16_and_1_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa11_and0 = s_CSAwallace_rca16_and_2_9 & s_CSAwallace_rca16_and_1_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa11_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_and_0_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa11_and1 = s_CSAwallace_rca16_csa3_csa_component_fa11_xor0 & s_CSAwallace_rca16_and_0_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa11_or0 = s_CSAwallace_rca16_csa3_csa_component_fa11_and0 | s_CSAwallace_rca16_csa3_csa_component_fa11_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa12_xor0 = s_CSAwallace_rca16_and_3_9 ^ s_CSAwallace_rca16_and_2_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa12_and0 = s_CSAwallace_rca16_and_3_9 & s_CSAwallace_rca16_and_2_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_and_1_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa12_and1 = s_CSAwallace_rca16_csa3_csa_component_fa12_xor0 & s_CSAwallace_rca16_and_1_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa12_or0 = s_CSAwallace_rca16_csa3_csa_component_fa12_and0 | s_CSAwallace_rca16_csa3_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa13_xor0 = s_CSAwallace_rca16_and_4_9 ^ s_CSAwallace_rca16_and_3_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa13_and0 = s_CSAwallace_rca16_and_4_9 & s_CSAwallace_rca16_and_3_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_and_2_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa13_and1 = s_CSAwallace_rca16_csa3_csa_component_fa13_xor0 & s_CSAwallace_rca16_and_2_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa13_or0 = s_CSAwallace_rca16_csa3_csa_component_fa13_and0 | s_CSAwallace_rca16_csa3_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa14_xor0 = s_CSAwallace_rca16_and_5_9 ^ s_CSAwallace_rca16_and_4_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa14_and0 = s_CSAwallace_rca16_and_5_9 & s_CSAwallace_rca16_and_4_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_and_3_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa14_and1 = s_CSAwallace_rca16_csa3_csa_component_fa14_xor0 & s_CSAwallace_rca16_and_3_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa14_or0 = s_CSAwallace_rca16_csa3_csa_component_fa14_and0 | s_CSAwallace_rca16_csa3_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa15_xor0 = s_CSAwallace_rca16_and_6_9 ^ s_CSAwallace_rca16_and_5_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa15_and0 = s_CSAwallace_rca16_and_6_9 & s_CSAwallace_rca16_and_5_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_and_4_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa15_and1 = s_CSAwallace_rca16_csa3_csa_component_fa15_xor0 & s_CSAwallace_rca16_and_4_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa15_or0 = s_CSAwallace_rca16_csa3_csa_component_fa15_and0 | s_CSAwallace_rca16_csa3_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa16_xor0 = s_CSAwallace_rca16_and_7_9 ^ s_CSAwallace_rca16_and_6_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa16_and0 = s_CSAwallace_rca16_and_7_9 & s_CSAwallace_rca16_and_6_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_and_5_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa16_and1 = s_CSAwallace_rca16_csa3_csa_component_fa16_xor0 & s_CSAwallace_rca16_and_5_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa16_or0 = s_CSAwallace_rca16_csa3_csa_component_fa16_and0 | s_CSAwallace_rca16_csa3_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa17_xor0 = s_CSAwallace_rca16_and_8_9 ^ s_CSAwallace_rca16_and_7_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa17_and0 = s_CSAwallace_rca16_and_8_9 & s_CSAwallace_rca16_and_7_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_and_6_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa17_and1 = s_CSAwallace_rca16_csa3_csa_component_fa17_xor0 & s_CSAwallace_rca16_and_6_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa17_or0 = s_CSAwallace_rca16_csa3_csa_component_fa17_and0 | s_CSAwallace_rca16_csa3_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa18_xor0 = s_CSAwallace_rca16_and_9_9 ^ s_CSAwallace_rca16_and_8_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa18_and0 = s_CSAwallace_rca16_and_9_9 & s_CSAwallace_rca16_and_8_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_and_7_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa18_and1 = s_CSAwallace_rca16_csa3_csa_component_fa18_xor0 & s_CSAwallace_rca16_and_7_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa18_or0 = s_CSAwallace_rca16_csa3_csa_component_fa18_and0 | s_CSAwallace_rca16_csa3_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa19_xor0 = s_CSAwallace_rca16_and_10_9 ^ s_CSAwallace_rca16_and_9_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa19_and0 = s_CSAwallace_rca16_and_10_9 & s_CSAwallace_rca16_and_9_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_and_8_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa19_and1 = s_CSAwallace_rca16_csa3_csa_component_fa19_xor0 & s_CSAwallace_rca16_and_8_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa19_or0 = s_CSAwallace_rca16_csa3_csa_component_fa19_and0 | s_CSAwallace_rca16_csa3_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa20_xor0 = s_CSAwallace_rca16_and_11_9 ^ s_CSAwallace_rca16_and_10_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa20_and0 = s_CSAwallace_rca16_and_11_9 & s_CSAwallace_rca16_and_10_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_and_9_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa20_and1 = s_CSAwallace_rca16_csa3_csa_component_fa20_xor0 & s_CSAwallace_rca16_and_9_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa20_or0 = s_CSAwallace_rca16_csa3_csa_component_fa20_and0 | s_CSAwallace_rca16_csa3_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa21_xor0 = s_CSAwallace_rca16_and_12_9 ^ s_CSAwallace_rca16_and_11_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa21_and0 = s_CSAwallace_rca16_and_12_9 & s_CSAwallace_rca16_and_11_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_and_10_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa21_and1 = s_CSAwallace_rca16_csa3_csa_component_fa21_xor0 & s_CSAwallace_rca16_and_10_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa21_or0 = s_CSAwallace_rca16_csa3_csa_component_fa21_and0 | s_CSAwallace_rca16_csa3_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa22_xor0 = s_CSAwallace_rca16_and_13_9 ^ s_CSAwallace_rca16_and_12_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa22_and0 = s_CSAwallace_rca16_and_13_9 & s_CSAwallace_rca16_and_12_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_and_11_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa22_and1 = s_CSAwallace_rca16_csa3_csa_component_fa22_xor0 & s_CSAwallace_rca16_and_11_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa22_or0 = s_CSAwallace_rca16_csa3_csa_component_fa22_and0 | s_CSAwallace_rca16_csa3_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa23_xor0 = s_CSAwallace_rca16_and_14_9 ^ s_CSAwallace_rca16_and_13_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa23_and0 = s_CSAwallace_rca16_and_14_9 & s_CSAwallace_rca16_and_13_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa23_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa23_xor0 ^ s_CSAwallace_rca16_and_12_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa23_and1 = s_CSAwallace_rca16_csa3_csa_component_fa23_xor0 & s_CSAwallace_rca16_and_12_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa23_or0 = s_CSAwallace_rca16_csa3_csa_component_fa23_and0 | s_CSAwallace_rca16_csa3_csa_component_fa23_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa24_xor0 = s_CSAwallace_rca16_nand_15_9 ^ s_CSAwallace_rca16_and_14_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa24_and0 = s_CSAwallace_rca16_nand_15_9 & s_CSAwallace_rca16_and_14_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa24_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa24_xor0 ^ s_CSAwallace_rca16_and_13_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa24_and1 = s_CSAwallace_rca16_csa3_csa_component_fa24_xor0 & s_CSAwallace_rca16_and_13_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa24_or0 = s_CSAwallace_rca16_csa3_csa_component_fa24_and0 | s_CSAwallace_rca16_csa3_csa_component_fa24_and1;
  assign s_CSAwallace_rca16_csa3_csa_component_fa25_xor0 = ~s_CSAwallace_rca16_nand_15_10;
  assign s_CSAwallace_rca16_csa3_csa_component_fa25_xor1 = s_CSAwallace_rca16_csa3_csa_component_fa25_xor0 ^ s_CSAwallace_rca16_and_14_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa25_and1 = s_CSAwallace_rca16_csa3_csa_component_fa25_xor0 & s_CSAwallace_rca16_and_14_11;
  assign s_CSAwallace_rca16_csa3_csa_component_fa25_or0 = s_CSAwallace_rca16_nand_15_10 | s_CSAwallace_rca16_csa3_csa_component_fa25_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa13_xor0 = s_CSAwallace_rca16_and_1_12 ^ s_CSAwallace_rca16_and_0_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa13_and0 = s_CSAwallace_rca16_and_1_12 & s_CSAwallace_rca16_and_0_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa14_xor0 = s_CSAwallace_rca16_and_2_12 ^ s_CSAwallace_rca16_and_1_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa14_and0 = s_CSAwallace_rca16_and_2_12 & s_CSAwallace_rca16_and_1_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_and_0_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa14_and1 = s_CSAwallace_rca16_csa4_csa_component_fa14_xor0 & s_CSAwallace_rca16_and_0_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa14_or0 = s_CSAwallace_rca16_csa4_csa_component_fa14_and0 | s_CSAwallace_rca16_csa4_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa15_xor0 = s_CSAwallace_rca16_and_3_12 ^ s_CSAwallace_rca16_and_2_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa15_and0 = s_CSAwallace_rca16_and_3_12 & s_CSAwallace_rca16_and_2_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_and_1_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa15_and1 = s_CSAwallace_rca16_csa4_csa_component_fa15_xor0 & s_CSAwallace_rca16_and_1_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa15_or0 = s_CSAwallace_rca16_csa4_csa_component_fa15_and0 | s_CSAwallace_rca16_csa4_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa16_xor0 = s_CSAwallace_rca16_and_4_12 ^ s_CSAwallace_rca16_and_3_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa16_and0 = s_CSAwallace_rca16_and_4_12 & s_CSAwallace_rca16_and_3_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_and_2_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa16_and1 = s_CSAwallace_rca16_csa4_csa_component_fa16_xor0 & s_CSAwallace_rca16_and_2_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa16_or0 = s_CSAwallace_rca16_csa4_csa_component_fa16_and0 | s_CSAwallace_rca16_csa4_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa17_xor0 = s_CSAwallace_rca16_and_5_12 ^ s_CSAwallace_rca16_and_4_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa17_and0 = s_CSAwallace_rca16_and_5_12 & s_CSAwallace_rca16_and_4_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_and_3_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa17_and1 = s_CSAwallace_rca16_csa4_csa_component_fa17_xor0 & s_CSAwallace_rca16_and_3_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa17_or0 = s_CSAwallace_rca16_csa4_csa_component_fa17_and0 | s_CSAwallace_rca16_csa4_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa18_xor0 = s_CSAwallace_rca16_and_6_12 ^ s_CSAwallace_rca16_and_5_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa18_and0 = s_CSAwallace_rca16_and_6_12 & s_CSAwallace_rca16_and_5_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_and_4_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa18_and1 = s_CSAwallace_rca16_csa4_csa_component_fa18_xor0 & s_CSAwallace_rca16_and_4_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa18_or0 = s_CSAwallace_rca16_csa4_csa_component_fa18_and0 | s_CSAwallace_rca16_csa4_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa19_xor0 = s_CSAwallace_rca16_and_7_12 ^ s_CSAwallace_rca16_and_6_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa19_and0 = s_CSAwallace_rca16_and_7_12 & s_CSAwallace_rca16_and_6_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_and_5_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa19_and1 = s_CSAwallace_rca16_csa4_csa_component_fa19_xor0 & s_CSAwallace_rca16_and_5_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa19_or0 = s_CSAwallace_rca16_csa4_csa_component_fa19_and0 | s_CSAwallace_rca16_csa4_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa20_xor0 = s_CSAwallace_rca16_and_8_12 ^ s_CSAwallace_rca16_and_7_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa20_and0 = s_CSAwallace_rca16_and_8_12 & s_CSAwallace_rca16_and_7_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_and_6_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa20_and1 = s_CSAwallace_rca16_csa4_csa_component_fa20_xor0 & s_CSAwallace_rca16_and_6_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa20_or0 = s_CSAwallace_rca16_csa4_csa_component_fa20_and0 | s_CSAwallace_rca16_csa4_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa21_xor0 = s_CSAwallace_rca16_and_9_12 ^ s_CSAwallace_rca16_and_8_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa21_and0 = s_CSAwallace_rca16_and_9_12 & s_CSAwallace_rca16_and_8_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_and_7_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa21_and1 = s_CSAwallace_rca16_csa4_csa_component_fa21_xor0 & s_CSAwallace_rca16_and_7_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa21_or0 = s_CSAwallace_rca16_csa4_csa_component_fa21_and0 | s_CSAwallace_rca16_csa4_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa22_xor0 = s_CSAwallace_rca16_and_10_12 ^ s_CSAwallace_rca16_and_9_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa22_and0 = s_CSAwallace_rca16_and_10_12 & s_CSAwallace_rca16_and_9_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_and_8_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa22_and1 = s_CSAwallace_rca16_csa4_csa_component_fa22_xor0 & s_CSAwallace_rca16_and_8_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa22_or0 = s_CSAwallace_rca16_csa4_csa_component_fa22_and0 | s_CSAwallace_rca16_csa4_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa23_xor0 = s_CSAwallace_rca16_and_11_12 ^ s_CSAwallace_rca16_and_10_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa23_and0 = s_CSAwallace_rca16_and_11_12 & s_CSAwallace_rca16_and_10_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa23_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa23_xor0 ^ s_CSAwallace_rca16_and_9_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa23_and1 = s_CSAwallace_rca16_csa4_csa_component_fa23_xor0 & s_CSAwallace_rca16_and_9_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa23_or0 = s_CSAwallace_rca16_csa4_csa_component_fa23_and0 | s_CSAwallace_rca16_csa4_csa_component_fa23_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa24_xor0 = s_CSAwallace_rca16_and_12_12 ^ s_CSAwallace_rca16_and_11_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa24_and0 = s_CSAwallace_rca16_and_12_12 & s_CSAwallace_rca16_and_11_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa24_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa24_xor0 ^ s_CSAwallace_rca16_and_10_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa24_and1 = s_CSAwallace_rca16_csa4_csa_component_fa24_xor0 & s_CSAwallace_rca16_and_10_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa24_or0 = s_CSAwallace_rca16_csa4_csa_component_fa24_and0 | s_CSAwallace_rca16_csa4_csa_component_fa24_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa25_xor0 = s_CSAwallace_rca16_and_13_12 ^ s_CSAwallace_rca16_and_12_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa25_and0 = s_CSAwallace_rca16_and_13_12 & s_CSAwallace_rca16_and_12_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa25_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa25_xor0 ^ s_CSAwallace_rca16_and_11_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa25_and1 = s_CSAwallace_rca16_csa4_csa_component_fa25_xor0 & s_CSAwallace_rca16_and_11_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa25_or0 = s_CSAwallace_rca16_csa4_csa_component_fa25_and0 | s_CSAwallace_rca16_csa4_csa_component_fa25_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa26_xor0 = s_CSAwallace_rca16_and_14_12 ^ s_CSAwallace_rca16_and_13_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa26_and0 = s_CSAwallace_rca16_and_14_12 & s_CSAwallace_rca16_and_13_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa26_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa26_xor0 ^ s_CSAwallace_rca16_and_12_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa26_and1 = s_CSAwallace_rca16_csa4_csa_component_fa26_xor0 & s_CSAwallace_rca16_and_12_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa26_or0 = s_CSAwallace_rca16_csa4_csa_component_fa26_and0 | s_CSAwallace_rca16_csa4_csa_component_fa26_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa27_xor0 = s_CSAwallace_rca16_nand_15_12 ^ s_CSAwallace_rca16_and_14_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa27_and0 = s_CSAwallace_rca16_nand_15_12 & s_CSAwallace_rca16_and_14_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa27_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa27_xor0 ^ s_CSAwallace_rca16_and_13_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa27_and1 = s_CSAwallace_rca16_csa4_csa_component_fa27_xor0 & s_CSAwallace_rca16_and_13_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa27_or0 = s_CSAwallace_rca16_csa4_csa_component_fa27_and0 | s_CSAwallace_rca16_csa4_csa_component_fa27_and1;
  assign s_CSAwallace_rca16_csa4_csa_component_fa28_xor0 = ~s_CSAwallace_rca16_nand_15_13;
  assign s_CSAwallace_rca16_csa4_csa_component_fa28_xor1 = s_CSAwallace_rca16_csa4_csa_component_fa28_xor0 ^ s_CSAwallace_rca16_and_14_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa28_and1 = s_CSAwallace_rca16_csa4_csa_component_fa28_xor0 & s_CSAwallace_rca16_and_14_14;
  assign s_CSAwallace_rca16_csa4_csa_component_fa28_or0 = s_CSAwallace_rca16_nand_15_13 | s_CSAwallace_rca16_csa4_csa_component_fa28_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa2_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa2_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa1_and0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa2_and0 = s_CSAwallace_rca16_csa0_csa_component_fa2_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa1_and0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa3_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa3_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa2_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa3_and0 = s_CSAwallace_rca16_csa0_csa_component_fa3_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa2_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa3_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa3_xor0 ^ s_CSAwallace_rca16_and_0_3;
  assign s_CSAwallace_rca16_csa5_csa_component_fa3_and1 = s_CSAwallace_rca16_csa5_csa_component_fa3_xor0 & s_CSAwallace_rca16_and_0_3;
  assign s_CSAwallace_rca16_csa5_csa_component_fa3_or0 = s_CSAwallace_rca16_csa5_csa_component_fa3_and0 | s_CSAwallace_rca16_csa5_csa_component_fa3_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa4_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa4_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa3_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa4_and0 = s_CSAwallace_rca16_csa0_csa_component_fa4_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa3_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa4_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa4_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa4_xor0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa4_and1 = s_CSAwallace_rca16_csa5_csa_component_fa4_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa4_xor0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa4_or0 = s_CSAwallace_rca16_csa5_csa_component_fa4_and0 | s_CSAwallace_rca16_csa5_csa_component_fa4_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa5_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa5_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa4_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa5_and0 = s_CSAwallace_rca16_csa0_csa_component_fa5_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa4_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa5_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa5_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa5_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa5_and1 = s_CSAwallace_rca16_csa5_csa_component_fa5_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa5_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa5_or0 = s_CSAwallace_rca16_csa5_csa_component_fa5_and0 | s_CSAwallace_rca16_csa5_csa_component_fa5_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa6_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa6_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa5_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa6_and0 = s_CSAwallace_rca16_csa0_csa_component_fa6_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa5_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa6_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa6_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa6_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa6_and1 = s_CSAwallace_rca16_csa5_csa_component_fa6_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa6_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa6_or0 = s_CSAwallace_rca16_csa5_csa_component_fa6_and0 | s_CSAwallace_rca16_csa5_csa_component_fa6_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa7_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa7_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa6_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa7_and0 = s_CSAwallace_rca16_csa0_csa_component_fa7_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa6_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa7_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa7_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa7_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa7_and1 = s_CSAwallace_rca16_csa5_csa_component_fa7_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa7_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa7_or0 = s_CSAwallace_rca16_csa5_csa_component_fa7_and0 | s_CSAwallace_rca16_csa5_csa_component_fa7_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa8_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa8_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa7_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa8_and0 = s_CSAwallace_rca16_csa0_csa_component_fa8_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa7_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa8_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa8_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa8_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa8_and1 = s_CSAwallace_rca16_csa5_csa_component_fa8_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa8_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa8_or0 = s_CSAwallace_rca16_csa5_csa_component_fa8_and0 | s_CSAwallace_rca16_csa5_csa_component_fa8_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa9_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa9_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa9_and0 = s_CSAwallace_rca16_csa0_csa_component_fa9_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa9_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa9_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa9_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa9_and1 = s_CSAwallace_rca16_csa5_csa_component_fa9_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa9_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa9_or0 = s_CSAwallace_rca16_csa5_csa_component_fa9_and0 | s_CSAwallace_rca16_csa5_csa_component_fa9_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa10_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa10_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa10_and0 = s_CSAwallace_rca16_csa0_csa_component_fa10_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa10_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa10_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa10_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa10_and1 = s_CSAwallace_rca16_csa5_csa_component_fa10_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa10_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa10_or0 = s_CSAwallace_rca16_csa5_csa_component_fa10_and0 | s_CSAwallace_rca16_csa5_csa_component_fa10_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa11_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa11_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa11_and0 = s_CSAwallace_rca16_csa0_csa_component_fa11_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa11_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa11_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa11_and1 = s_CSAwallace_rca16_csa5_csa_component_fa11_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa11_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa11_or0 = s_CSAwallace_rca16_csa5_csa_component_fa11_and0 | s_CSAwallace_rca16_csa5_csa_component_fa11_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa12_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa12_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa12_and0 = s_CSAwallace_rca16_csa0_csa_component_fa12_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa12_and1 = s_CSAwallace_rca16_csa5_csa_component_fa12_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa12_or0 = s_CSAwallace_rca16_csa5_csa_component_fa12_and0 | s_CSAwallace_rca16_csa5_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa13_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa13_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa13_and0 = s_CSAwallace_rca16_csa0_csa_component_fa13_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa13_and1 = s_CSAwallace_rca16_csa5_csa_component_fa13_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa13_or0 = s_CSAwallace_rca16_csa5_csa_component_fa13_and0 | s_CSAwallace_rca16_csa5_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa14_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa14_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa14_and0 = s_CSAwallace_rca16_csa0_csa_component_fa14_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa14_and1 = s_CSAwallace_rca16_csa5_csa_component_fa14_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa14_or0 = s_CSAwallace_rca16_csa5_csa_component_fa14_and0 | s_CSAwallace_rca16_csa5_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa15_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa15_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa15_and0 = s_CSAwallace_rca16_csa0_csa_component_fa15_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa15_and1 = s_CSAwallace_rca16_csa5_csa_component_fa15_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa15_or0 = s_CSAwallace_rca16_csa5_csa_component_fa15_and0 | s_CSAwallace_rca16_csa5_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa16_xor0 = s_CSAwallace_rca16_csa0_csa_component_fa16_xor1 ^ s_CSAwallace_rca16_csa0_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa16_and0 = s_CSAwallace_rca16_csa0_csa_component_fa16_xor1 & s_CSAwallace_rca16_csa0_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa16_and1 = s_CSAwallace_rca16_csa5_csa_component_fa16_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa16_or0 = s_CSAwallace_rca16_csa5_csa_component_fa16_and0 | s_CSAwallace_rca16_csa5_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa17_xor0 = s_CSAwallace_rca16_nand_15_2 ^ s_CSAwallace_rca16_csa0_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa17_and0 = s_CSAwallace_rca16_nand_15_2 & s_CSAwallace_rca16_csa0_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa5_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa5_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa17_and1 = s_CSAwallace_rca16_csa5_csa_component_fa17_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa5_csa_component_fa17_or0 = s_CSAwallace_rca16_csa5_csa_component_fa17_and0 | s_CSAwallace_rca16_csa5_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa6_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa5_or0 ^ s_CSAwallace_rca16_and_0_6;
  assign s_CSAwallace_rca16_csa6_csa_component_fa6_and0 = s_CSAwallace_rca16_csa1_csa_component_fa5_or0 & s_CSAwallace_rca16_and_0_6;
  assign s_CSAwallace_rca16_csa6_csa_component_fa7_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa6_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa7_xor0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa7_and0 = s_CSAwallace_rca16_csa1_csa_component_fa6_or0 & s_CSAwallace_rca16_csa2_csa_component_fa7_xor0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa8_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa7_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa8_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa8_and0 = s_CSAwallace_rca16_csa1_csa_component_fa7_or0 & s_CSAwallace_rca16_csa2_csa_component_fa8_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa8_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa8_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa7_and0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa8_and1 = s_CSAwallace_rca16_csa6_csa_component_fa8_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa7_and0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa8_or0 = s_CSAwallace_rca16_csa6_csa_component_fa8_and0 | s_CSAwallace_rca16_csa6_csa_component_fa8_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa9_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa8_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa9_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa9_and0 = s_CSAwallace_rca16_csa1_csa_component_fa8_or0 & s_CSAwallace_rca16_csa2_csa_component_fa9_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa9_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa9_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa9_and1 = s_CSAwallace_rca16_csa6_csa_component_fa9_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa9_or0 = s_CSAwallace_rca16_csa6_csa_component_fa9_and0 | s_CSAwallace_rca16_csa6_csa_component_fa9_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa10_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa9_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa10_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa10_and0 = s_CSAwallace_rca16_csa1_csa_component_fa9_or0 & s_CSAwallace_rca16_csa2_csa_component_fa10_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa10_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa10_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa10_and1 = s_CSAwallace_rca16_csa6_csa_component_fa10_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa10_or0 = s_CSAwallace_rca16_csa6_csa_component_fa10_and0 | s_CSAwallace_rca16_csa6_csa_component_fa10_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa11_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa10_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa11_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa11_and0 = s_CSAwallace_rca16_csa1_csa_component_fa10_or0 & s_CSAwallace_rca16_csa2_csa_component_fa11_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa11_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa11_and1 = s_CSAwallace_rca16_csa6_csa_component_fa11_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa11_or0 = s_CSAwallace_rca16_csa6_csa_component_fa11_and0 | s_CSAwallace_rca16_csa6_csa_component_fa11_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa12_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa11_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa12_and0 = s_CSAwallace_rca16_csa1_csa_component_fa11_or0 & s_CSAwallace_rca16_csa2_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa12_and1 = s_CSAwallace_rca16_csa6_csa_component_fa12_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa12_or0 = s_CSAwallace_rca16_csa6_csa_component_fa12_and0 | s_CSAwallace_rca16_csa6_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa13_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa12_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa13_and0 = s_CSAwallace_rca16_csa1_csa_component_fa12_or0 & s_CSAwallace_rca16_csa2_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa13_and1 = s_CSAwallace_rca16_csa6_csa_component_fa13_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa13_or0 = s_CSAwallace_rca16_csa6_csa_component_fa13_and0 | s_CSAwallace_rca16_csa6_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa14_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa13_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa14_and0 = s_CSAwallace_rca16_csa1_csa_component_fa13_or0 & s_CSAwallace_rca16_csa2_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa14_and1 = s_CSAwallace_rca16_csa6_csa_component_fa14_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa14_or0 = s_CSAwallace_rca16_csa6_csa_component_fa14_and0 | s_CSAwallace_rca16_csa6_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa15_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa14_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa15_and0 = s_CSAwallace_rca16_csa1_csa_component_fa14_or0 & s_CSAwallace_rca16_csa2_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa15_and1 = s_CSAwallace_rca16_csa6_csa_component_fa15_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa15_or0 = s_CSAwallace_rca16_csa6_csa_component_fa15_and0 | s_CSAwallace_rca16_csa6_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa16_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa15_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa16_and0 = s_CSAwallace_rca16_csa1_csa_component_fa15_or0 & s_CSAwallace_rca16_csa2_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa16_and1 = s_CSAwallace_rca16_csa6_csa_component_fa16_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa16_or0 = s_CSAwallace_rca16_csa6_csa_component_fa16_and0 | s_CSAwallace_rca16_csa6_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa17_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa16_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa17_and0 = s_CSAwallace_rca16_csa1_csa_component_fa16_or0 & s_CSAwallace_rca16_csa2_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa17_and1 = s_CSAwallace_rca16_csa6_csa_component_fa17_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa17_or0 = s_CSAwallace_rca16_csa6_csa_component_fa17_and0 | s_CSAwallace_rca16_csa6_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa18_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa17_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa18_and0 = s_CSAwallace_rca16_csa1_csa_component_fa17_or0 & s_CSAwallace_rca16_csa2_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa18_and1 = s_CSAwallace_rca16_csa6_csa_component_fa18_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa18_or0 = s_CSAwallace_rca16_csa6_csa_component_fa18_and0 | s_CSAwallace_rca16_csa6_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa19_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa18_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa19_and0 = s_CSAwallace_rca16_csa1_csa_component_fa18_or0 & s_CSAwallace_rca16_csa2_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa19_and1 = s_CSAwallace_rca16_csa6_csa_component_fa19_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa19_or0 = s_CSAwallace_rca16_csa6_csa_component_fa19_and0 | s_CSAwallace_rca16_csa6_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa20_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa19_or0 ^ s_CSAwallace_rca16_csa2_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa20_and0 = s_CSAwallace_rca16_csa1_csa_component_fa19_or0 & s_CSAwallace_rca16_csa2_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa20_and1 = s_CSAwallace_rca16_csa6_csa_component_fa20_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa20_or0 = s_CSAwallace_rca16_csa6_csa_component_fa20_and0 | s_CSAwallace_rca16_csa6_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa21_xor0 = ~s_CSAwallace_rca16_csa2_csa_component_fa21_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa21_and1 = s_CSAwallace_rca16_csa6_csa_component_fa21_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa21_or0 = s_CSAwallace_rca16_csa2_csa_component_fa21_xor1 | s_CSAwallace_rca16_csa6_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa22_xor0 = ~s_CSAwallace_rca16_csa2_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa22_and1 = s_CSAwallace_rca16_csa6_csa_component_fa22_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa22_or0 = s_CSAwallace_rca16_csa2_csa_component_fa22_xor1 | s_CSAwallace_rca16_csa6_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa6_csa_component_fa23_xor0 = ~s_CSAwallace_rca16_nand_15_8;
  assign s_CSAwallace_rca16_csa6_csa_component_fa23_xor1 = s_CSAwallace_rca16_csa6_csa_component_fa23_xor0 ^ s_CSAwallace_rca16_csa2_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa23_and1 = s_CSAwallace_rca16_csa6_csa_component_fa23_xor0 & s_CSAwallace_rca16_csa2_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa6_csa_component_fa23_or0 = s_CSAwallace_rca16_nand_15_8 | s_CSAwallace_rca16_csa6_csa_component_fa23_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa11_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa11_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa10_and0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa11_and0 = s_CSAwallace_rca16_csa3_csa_component_fa11_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa10_and0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa12_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa12_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa12_and0 = s_CSAwallace_rca16_csa3_csa_component_fa12_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_and_0_12;
  assign s_CSAwallace_rca16_csa7_csa_component_fa12_and1 = s_CSAwallace_rca16_csa7_csa_component_fa12_xor0 & s_CSAwallace_rca16_and_0_12;
  assign s_CSAwallace_rca16_csa7_csa_component_fa12_or0 = s_CSAwallace_rca16_csa7_csa_component_fa12_and0 | s_CSAwallace_rca16_csa7_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa13_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa13_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa13_and0 = s_CSAwallace_rca16_csa3_csa_component_fa13_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa13_xor0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa13_and1 = s_CSAwallace_rca16_csa7_csa_component_fa13_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa13_xor0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa13_or0 = s_CSAwallace_rca16_csa7_csa_component_fa13_and0 | s_CSAwallace_rca16_csa7_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa14_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa14_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa14_and0 = s_CSAwallace_rca16_csa3_csa_component_fa14_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa14_and1 = s_CSAwallace_rca16_csa7_csa_component_fa14_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa14_or0 = s_CSAwallace_rca16_csa7_csa_component_fa14_and0 | s_CSAwallace_rca16_csa7_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa15_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa15_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa15_and0 = s_CSAwallace_rca16_csa3_csa_component_fa15_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa15_and1 = s_CSAwallace_rca16_csa7_csa_component_fa15_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa15_or0 = s_CSAwallace_rca16_csa7_csa_component_fa15_and0 | s_CSAwallace_rca16_csa7_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa16_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa16_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa16_and0 = s_CSAwallace_rca16_csa3_csa_component_fa16_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa16_and1 = s_CSAwallace_rca16_csa7_csa_component_fa16_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa16_or0 = s_CSAwallace_rca16_csa7_csa_component_fa16_and0 | s_CSAwallace_rca16_csa7_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa17_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa17_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa17_and0 = s_CSAwallace_rca16_csa3_csa_component_fa17_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa17_and1 = s_CSAwallace_rca16_csa7_csa_component_fa17_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa17_or0 = s_CSAwallace_rca16_csa7_csa_component_fa17_and0 | s_CSAwallace_rca16_csa7_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa18_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa18_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa18_and0 = s_CSAwallace_rca16_csa3_csa_component_fa18_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa18_and1 = s_CSAwallace_rca16_csa7_csa_component_fa18_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa18_or0 = s_CSAwallace_rca16_csa7_csa_component_fa18_and0 | s_CSAwallace_rca16_csa7_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa19_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa19_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa19_and0 = s_CSAwallace_rca16_csa3_csa_component_fa19_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa19_and1 = s_CSAwallace_rca16_csa7_csa_component_fa19_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa19_or0 = s_CSAwallace_rca16_csa7_csa_component_fa19_and0 | s_CSAwallace_rca16_csa7_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa20_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa20_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa20_and0 = s_CSAwallace_rca16_csa3_csa_component_fa20_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa20_and1 = s_CSAwallace_rca16_csa7_csa_component_fa20_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa20_or0 = s_CSAwallace_rca16_csa7_csa_component_fa20_and0 | s_CSAwallace_rca16_csa7_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa21_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa21_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa21_and0 = s_CSAwallace_rca16_csa3_csa_component_fa21_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa21_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa21_and1 = s_CSAwallace_rca16_csa7_csa_component_fa21_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa21_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa21_or0 = s_CSAwallace_rca16_csa7_csa_component_fa21_and0 | s_CSAwallace_rca16_csa7_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa22_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa22_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa22_and0 = s_CSAwallace_rca16_csa3_csa_component_fa22_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa22_and1 = s_CSAwallace_rca16_csa7_csa_component_fa22_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa22_or0 = s_CSAwallace_rca16_csa7_csa_component_fa22_and0 | s_CSAwallace_rca16_csa7_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa23_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa23_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa23_and0 = s_CSAwallace_rca16_csa3_csa_component_fa23_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa23_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa23_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa23_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa23_and1 = s_CSAwallace_rca16_csa7_csa_component_fa23_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa23_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa23_or0 = s_CSAwallace_rca16_csa7_csa_component_fa23_and0 | s_CSAwallace_rca16_csa7_csa_component_fa23_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa24_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa24_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa24_and0 = s_CSAwallace_rca16_csa3_csa_component_fa24_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa24_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa24_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa24_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa24_and1 = s_CSAwallace_rca16_csa7_csa_component_fa24_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa24_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa24_or0 = s_CSAwallace_rca16_csa7_csa_component_fa24_and0 | s_CSAwallace_rca16_csa7_csa_component_fa24_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa25_xor0 = s_CSAwallace_rca16_csa3_csa_component_fa25_xor1 ^ s_CSAwallace_rca16_csa3_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa25_and0 = s_CSAwallace_rca16_csa3_csa_component_fa25_xor1 & s_CSAwallace_rca16_csa3_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa25_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa25_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa25_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa25_and1 = s_CSAwallace_rca16_csa7_csa_component_fa25_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa25_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa25_or0 = s_CSAwallace_rca16_csa7_csa_component_fa25_and0 | s_CSAwallace_rca16_csa7_csa_component_fa25_and1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa26_xor0 = s_CSAwallace_rca16_nand_15_11 ^ s_CSAwallace_rca16_csa3_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa26_and0 = s_CSAwallace_rca16_nand_15_11 & s_CSAwallace_rca16_csa3_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa7_csa_component_fa26_xor1 = s_CSAwallace_rca16_csa7_csa_component_fa26_xor0 ^ s_CSAwallace_rca16_csa4_csa_component_fa26_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa26_and1 = s_CSAwallace_rca16_csa7_csa_component_fa26_xor0 & s_CSAwallace_rca16_csa4_csa_component_fa26_xor1;
  assign s_CSAwallace_rca16_csa7_csa_component_fa26_or0 = s_CSAwallace_rca16_csa7_csa_component_fa26_and0 | s_CSAwallace_rca16_csa7_csa_component_fa26_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa3_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa3_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa2_and0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa3_and0 = s_CSAwallace_rca16_csa5_csa_component_fa3_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa2_and0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa4_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa4_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa3_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa4_and0 = s_CSAwallace_rca16_csa5_csa_component_fa4_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa3_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa5_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa5_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa4_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa5_and0 = s_CSAwallace_rca16_csa5_csa_component_fa5_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa4_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa5_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa5_xor0 ^ s_CSAwallace_rca16_csa1_csa_component_fa4_and0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa5_and1 = s_CSAwallace_rca16_csa8_csa_component_fa5_xor0 & s_CSAwallace_rca16_csa1_csa_component_fa4_and0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa5_or0 = s_CSAwallace_rca16_csa8_csa_component_fa5_and0 | s_CSAwallace_rca16_csa8_csa_component_fa5_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa6_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa6_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa5_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa6_and0 = s_CSAwallace_rca16_csa5_csa_component_fa6_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa5_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa6_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa6_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa6_xor0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa6_and1 = s_CSAwallace_rca16_csa8_csa_component_fa6_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa6_xor0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa6_or0 = s_CSAwallace_rca16_csa8_csa_component_fa6_and0 | s_CSAwallace_rca16_csa8_csa_component_fa6_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa7_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa7_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa6_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa7_and0 = s_CSAwallace_rca16_csa5_csa_component_fa7_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa6_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa7_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa7_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa7_xor0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa7_and1 = s_CSAwallace_rca16_csa8_csa_component_fa7_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa7_xor0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa7_or0 = s_CSAwallace_rca16_csa8_csa_component_fa7_and0 | s_CSAwallace_rca16_csa8_csa_component_fa7_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa8_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa8_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa7_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa8_and0 = s_CSAwallace_rca16_csa5_csa_component_fa8_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa7_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa8_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa8_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa8_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa8_and1 = s_CSAwallace_rca16_csa8_csa_component_fa8_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa8_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa8_or0 = s_CSAwallace_rca16_csa8_csa_component_fa8_and0 | s_CSAwallace_rca16_csa8_csa_component_fa8_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa9_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa9_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa9_and0 = s_CSAwallace_rca16_csa5_csa_component_fa9_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa9_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa9_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa9_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa9_and1 = s_CSAwallace_rca16_csa8_csa_component_fa9_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa9_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa9_or0 = s_CSAwallace_rca16_csa8_csa_component_fa9_and0 | s_CSAwallace_rca16_csa8_csa_component_fa9_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa10_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa10_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa10_and0 = s_CSAwallace_rca16_csa5_csa_component_fa10_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa10_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa10_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa10_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa10_and1 = s_CSAwallace_rca16_csa8_csa_component_fa10_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa10_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa10_or0 = s_CSAwallace_rca16_csa8_csa_component_fa10_and0 | s_CSAwallace_rca16_csa8_csa_component_fa10_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa11_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa11_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa11_and0 = s_CSAwallace_rca16_csa5_csa_component_fa11_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa11_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa11_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa11_and1 = s_CSAwallace_rca16_csa8_csa_component_fa11_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa11_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa11_or0 = s_CSAwallace_rca16_csa8_csa_component_fa11_and0 | s_CSAwallace_rca16_csa8_csa_component_fa11_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa12_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa12_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa12_and0 = s_CSAwallace_rca16_csa5_csa_component_fa12_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa12_and1 = s_CSAwallace_rca16_csa8_csa_component_fa12_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa12_or0 = s_CSAwallace_rca16_csa8_csa_component_fa12_and0 | s_CSAwallace_rca16_csa8_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa13_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa13_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa13_and0 = s_CSAwallace_rca16_csa5_csa_component_fa13_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa13_and1 = s_CSAwallace_rca16_csa8_csa_component_fa13_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa13_or0 = s_CSAwallace_rca16_csa8_csa_component_fa13_and0 | s_CSAwallace_rca16_csa8_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa14_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa14_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa14_and0 = s_CSAwallace_rca16_csa5_csa_component_fa14_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa14_and1 = s_CSAwallace_rca16_csa8_csa_component_fa14_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa14_or0 = s_CSAwallace_rca16_csa8_csa_component_fa14_and0 | s_CSAwallace_rca16_csa8_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa15_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa15_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa15_and0 = s_CSAwallace_rca16_csa5_csa_component_fa15_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa15_and1 = s_CSAwallace_rca16_csa8_csa_component_fa15_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa15_or0 = s_CSAwallace_rca16_csa8_csa_component_fa15_and0 | s_CSAwallace_rca16_csa8_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa16_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa16_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa16_and0 = s_CSAwallace_rca16_csa5_csa_component_fa16_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa16_and1 = s_CSAwallace_rca16_csa8_csa_component_fa16_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa16_or0 = s_CSAwallace_rca16_csa8_csa_component_fa16_and0 | s_CSAwallace_rca16_csa8_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa17_xor0 = s_CSAwallace_rca16_csa5_csa_component_fa17_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa17_and0 = s_CSAwallace_rca16_csa5_csa_component_fa17_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa17_and1 = s_CSAwallace_rca16_csa8_csa_component_fa17_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa17_or0 = s_CSAwallace_rca16_csa8_csa_component_fa17_and0 | s_CSAwallace_rca16_csa8_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa18_xor0 = s_CSAwallace_rca16_csa1_csa_component_fa18_xor1 ^ s_CSAwallace_rca16_csa5_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa18_and0 = s_CSAwallace_rca16_csa1_csa_component_fa18_xor1 & s_CSAwallace_rca16_csa5_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa8_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa18_and1 = s_CSAwallace_rca16_csa8_csa_component_fa18_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa18_or0 = s_CSAwallace_rca16_csa8_csa_component_fa18_and0 | s_CSAwallace_rca16_csa8_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa19_xor0 = ~s_CSAwallace_rca16_csa1_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa19_and1 = s_CSAwallace_rca16_csa8_csa_component_fa19_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa19_or0 = s_CSAwallace_rca16_csa1_csa_component_fa19_xor1 | s_CSAwallace_rca16_csa8_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa20_xor0 = ~s_CSAwallace_rca16_nand_15_5;
  assign s_CSAwallace_rca16_csa8_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa8_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa20_and1 = s_CSAwallace_rca16_csa8_csa_component_fa20_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa8_csa_component_fa20_or0 = s_CSAwallace_rca16_nand_15_5 | s_CSAwallace_rca16_csa8_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa9_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa8_or0 ^ s_CSAwallace_rca16_and_0_9;
  assign s_CSAwallace_rca16_csa9_csa_component_fa9_and0 = s_CSAwallace_rca16_csa6_csa_component_fa8_or0 & s_CSAwallace_rca16_and_0_9;
  assign s_CSAwallace_rca16_csa9_csa_component_fa10_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa9_or0 ^ s_CSAwallace_rca16_csa3_csa_component_fa10_xor0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa10_and0 = s_CSAwallace_rca16_csa6_csa_component_fa9_or0 & s_CSAwallace_rca16_csa3_csa_component_fa10_xor0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa11_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa10_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa11_xor0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa11_and0 = s_CSAwallace_rca16_csa6_csa_component_fa10_or0 & s_CSAwallace_rca16_csa7_csa_component_fa11_xor0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa12_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa11_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa12_and0 = s_CSAwallace_rca16_csa6_csa_component_fa11_or0 & s_CSAwallace_rca16_csa7_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa11_and0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa12_and1 = s_CSAwallace_rca16_csa9_csa_component_fa12_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa11_and0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa12_or0 = s_CSAwallace_rca16_csa9_csa_component_fa12_and0 | s_CSAwallace_rca16_csa9_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa13_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa12_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa13_and0 = s_CSAwallace_rca16_csa6_csa_component_fa12_or0 & s_CSAwallace_rca16_csa7_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa13_and1 = s_CSAwallace_rca16_csa9_csa_component_fa13_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa13_or0 = s_CSAwallace_rca16_csa9_csa_component_fa13_and0 | s_CSAwallace_rca16_csa9_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa14_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa13_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa14_and0 = s_CSAwallace_rca16_csa6_csa_component_fa13_or0 & s_CSAwallace_rca16_csa7_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa14_and1 = s_CSAwallace_rca16_csa9_csa_component_fa14_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa14_or0 = s_CSAwallace_rca16_csa9_csa_component_fa14_and0 | s_CSAwallace_rca16_csa9_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa15_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa14_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa15_and0 = s_CSAwallace_rca16_csa6_csa_component_fa14_or0 & s_CSAwallace_rca16_csa7_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa15_and1 = s_CSAwallace_rca16_csa9_csa_component_fa15_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa15_or0 = s_CSAwallace_rca16_csa9_csa_component_fa15_and0 | s_CSAwallace_rca16_csa9_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa16_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa15_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa16_and0 = s_CSAwallace_rca16_csa6_csa_component_fa15_or0 & s_CSAwallace_rca16_csa7_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa16_and1 = s_CSAwallace_rca16_csa9_csa_component_fa16_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa16_or0 = s_CSAwallace_rca16_csa9_csa_component_fa16_and0 | s_CSAwallace_rca16_csa9_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa17_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa16_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa17_and0 = s_CSAwallace_rca16_csa6_csa_component_fa16_or0 & s_CSAwallace_rca16_csa7_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa17_and1 = s_CSAwallace_rca16_csa9_csa_component_fa17_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa17_or0 = s_CSAwallace_rca16_csa9_csa_component_fa17_and0 | s_CSAwallace_rca16_csa9_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa18_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa17_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa18_and0 = s_CSAwallace_rca16_csa6_csa_component_fa17_or0 & s_CSAwallace_rca16_csa7_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa18_and1 = s_CSAwallace_rca16_csa9_csa_component_fa18_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa18_or0 = s_CSAwallace_rca16_csa9_csa_component_fa18_and0 | s_CSAwallace_rca16_csa9_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa19_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa18_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa19_and0 = s_CSAwallace_rca16_csa6_csa_component_fa18_or0 & s_CSAwallace_rca16_csa7_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa19_and1 = s_CSAwallace_rca16_csa9_csa_component_fa19_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa19_or0 = s_CSAwallace_rca16_csa9_csa_component_fa19_and0 | s_CSAwallace_rca16_csa9_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa20_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa19_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa20_and0 = s_CSAwallace_rca16_csa6_csa_component_fa19_or0 & s_CSAwallace_rca16_csa7_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa20_and1 = s_CSAwallace_rca16_csa9_csa_component_fa20_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa20_or0 = s_CSAwallace_rca16_csa9_csa_component_fa20_and0 | s_CSAwallace_rca16_csa9_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa21_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa20_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa21_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa21_and0 = s_CSAwallace_rca16_csa6_csa_component_fa20_or0 & s_CSAwallace_rca16_csa7_csa_component_fa21_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa21_and1 = s_CSAwallace_rca16_csa9_csa_component_fa21_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa21_or0 = s_CSAwallace_rca16_csa9_csa_component_fa21_and0 | s_CSAwallace_rca16_csa9_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa22_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa21_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa22_and0 = s_CSAwallace_rca16_csa6_csa_component_fa21_or0 & s_CSAwallace_rca16_csa7_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa22_and1 = s_CSAwallace_rca16_csa9_csa_component_fa22_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa22_or0 = s_CSAwallace_rca16_csa9_csa_component_fa22_and0 | s_CSAwallace_rca16_csa9_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa23_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa22_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa23_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa23_and0 = s_CSAwallace_rca16_csa6_csa_component_fa22_or0 & s_CSAwallace_rca16_csa7_csa_component_fa23_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa23_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa23_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa23_and1 = s_CSAwallace_rca16_csa9_csa_component_fa23_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa23_or0 = s_CSAwallace_rca16_csa9_csa_component_fa23_and0 | s_CSAwallace_rca16_csa9_csa_component_fa23_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa24_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa23_or0 ^ s_CSAwallace_rca16_csa7_csa_component_fa24_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa24_and0 = s_CSAwallace_rca16_csa6_csa_component_fa23_or0 & s_CSAwallace_rca16_csa7_csa_component_fa24_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa24_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa24_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa24_and1 = s_CSAwallace_rca16_csa9_csa_component_fa24_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa24_or0 = s_CSAwallace_rca16_csa9_csa_component_fa24_and0 | s_CSAwallace_rca16_csa9_csa_component_fa24_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa25_xor0 = ~s_CSAwallace_rca16_csa7_csa_component_fa25_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa25_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa25_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa25_and1 = s_CSAwallace_rca16_csa9_csa_component_fa25_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa25_or0 = s_CSAwallace_rca16_csa7_csa_component_fa25_xor1 | s_CSAwallace_rca16_csa9_csa_component_fa25_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa26_xor0 = ~s_CSAwallace_rca16_csa7_csa_component_fa26_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa26_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa26_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa26_and1 = s_CSAwallace_rca16_csa9_csa_component_fa26_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa26_or0 = s_CSAwallace_rca16_csa7_csa_component_fa26_xor1 | s_CSAwallace_rca16_csa9_csa_component_fa26_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa27_xor0 = ~s_CSAwallace_rca16_csa4_csa_component_fa27_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa27_xor1 = s_CSAwallace_rca16_csa9_csa_component_fa27_xor0 ^ s_CSAwallace_rca16_csa7_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa27_and1 = s_CSAwallace_rca16_csa9_csa_component_fa27_xor0 & s_CSAwallace_rca16_csa7_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa27_or0 = s_CSAwallace_rca16_csa4_csa_component_fa27_xor1 | s_CSAwallace_rca16_csa9_csa_component_fa27_and1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa28_xor0 = ~s_CSAwallace_rca16_csa4_csa_component_fa28_xor1;
  assign s_CSAwallace_rca16_csa9_csa_component_fa28_xor1 = ~s_CSAwallace_rca16_csa9_csa_component_fa28_xor0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa28_or0 = s_CSAwallace_rca16_csa4_csa_component_fa28_xor1 | s_CSAwallace_rca16_csa9_csa_component_fa28_xor0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa29_xor0 = ~s_CSAwallace_rca16_nand_15_14;
  assign s_CSAwallace_rca16_csa9_csa_component_fa29_xor1 = ~s_CSAwallace_rca16_csa9_csa_component_fa29_xor0;
  assign s_CSAwallace_rca16_csa9_csa_component_fa29_or0 = s_CSAwallace_rca16_nand_15_14 | s_CSAwallace_rca16_csa9_csa_component_fa29_xor0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa4_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa4_xor0 ^ s_CSAwallace_rca16_csa8_csa_component_fa3_and0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa4_and0 = s_CSAwallace_rca16_csa8_csa_component_fa4_xor0 & s_CSAwallace_rca16_csa8_csa_component_fa3_and0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa5_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa5_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa4_and0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa5_and0 = s_CSAwallace_rca16_csa8_csa_component_fa5_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa4_and0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa6_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa6_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa5_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa6_and0 = s_CSAwallace_rca16_csa8_csa_component_fa6_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa5_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa7_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa7_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa6_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa7_and0 = s_CSAwallace_rca16_csa8_csa_component_fa7_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa6_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa7_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa7_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa6_and0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa7_and1 = s_CSAwallace_rca16_csa10_csa_component_fa7_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa6_and0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa7_or0 = s_CSAwallace_rca16_csa10_csa_component_fa7_and0 | s_CSAwallace_rca16_csa10_csa_component_fa7_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa8_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa8_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa7_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa8_and0 = s_CSAwallace_rca16_csa8_csa_component_fa8_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa7_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa8_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa8_xor0 ^ s_CSAwallace_rca16_csa6_csa_component_fa7_and0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa8_and1 = s_CSAwallace_rca16_csa10_csa_component_fa8_xor0 & s_CSAwallace_rca16_csa6_csa_component_fa7_and0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa8_or0 = s_CSAwallace_rca16_csa10_csa_component_fa8_and0 | s_CSAwallace_rca16_csa10_csa_component_fa8_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa9_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa9_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa9_and0 = s_CSAwallace_rca16_csa8_csa_component_fa9_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa9_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa9_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa9_xor0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa9_and1 = s_CSAwallace_rca16_csa10_csa_component_fa9_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa9_xor0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa9_or0 = s_CSAwallace_rca16_csa10_csa_component_fa9_and0 | s_CSAwallace_rca16_csa10_csa_component_fa9_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa10_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa10_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa10_and0 = s_CSAwallace_rca16_csa8_csa_component_fa10_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa10_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa10_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa10_xor0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa10_and1 = s_CSAwallace_rca16_csa10_csa_component_fa10_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa10_xor0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa10_or0 = s_CSAwallace_rca16_csa10_csa_component_fa10_and0 | s_CSAwallace_rca16_csa10_csa_component_fa10_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa11_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa11_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa11_and0 = s_CSAwallace_rca16_csa8_csa_component_fa11_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa11_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa11_xor0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa11_and1 = s_CSAwallace_rca16_csa10_csa_component_fa11_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa11_xor0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa11_or0 = s_CSAwallace_rca16_csa10_csa_component_fa11_and0 | s_CSAwallace_rca16_csa10_csa_component_fa11_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa12_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa12_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa12_and0 = s_CSAwallace_rca16_csa8_csa_component_fa12_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa12_and1 = s_CSAwallace_rca16_csa10_csa_component_fa12_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa12_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa12_or0 = s_CSAwallace_rca16_csa10_csa_component_fa12_and0 | s_CSAwallace_rca16_csa10_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa13_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa13_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa13_and0 = s_CSAwallace_rca16_csa8_csa_component_fa13_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa13_and1 = s_CSAwallace_rca16_csa10_csa_component_fa13_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa13_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa13_or0 = s_CSAwallace_rca16_csa10_csa_component_fa13_and0 | s_CSAwallace_rca16_csa10_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa14_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa14_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa14_and0 = s_CSAwallace_rca16_csa8_csa_component_fa14_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa14_and1 = s_CSAwallace_rca16_csa10_csa_component_fa14_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa14_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa14_or0 = s_CSAwallace_rca16_csa10_csa_component_fa14_and0 | s_CSAwallace_rca16_csa10_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa15_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa15_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa15_and0 = s_CSAwallace_rca16_csa8_csa_component_fa15_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa15_and1 = s_CSAwallace_rca16_csa10_csa_component_fa15_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa15_or0 = s_CSAwallace_rca16_csa10_csa_component_fa15_and0 | s_CSAwallace_rca16_csa10_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa16_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa16_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa16_and0 = s_CSAwallace_rca16_csa8_csa_component_fa16_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa16_and1 = s_CSAwallace_rca16_csa10_csa_component_fa16_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa16_or0 = s_CSAwallace_rca16_csa10_csa_component_fa16_and0 | s_CSAwallace_rca16_csa10_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa17_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa17_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa17_and0 = s_CSAwallace_rca16_csa8_csa_component_fa17_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa17_and1 = s_CSAwallace_rca16_csa10_csa_component_fa17_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa17_or0 = s_CSAwallace_rca16_csa10_csa_component_fa17_and0 | s_CSAwallace_rca16_csa10_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa18_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa18_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa18_and0 = s_CSAwallace_rca16_csa8_csa_component_fa18_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa18_and1 = s_CSAwallace_rca16_csa10_csa_component_fa18_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa18_or0 = s_CSAwallace_rca16_csa10_csa_component_fa18_and0 | s_CSAwallace_rca16_csa10_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa19_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa19_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa19_and0 = s_CSAwallace_rca16_csa8_csa_component_fa19_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa19_and1 = s_CSAwallace_rca16_csa10_csa_component_fa19_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa19_or0 = s_CSAwallace_rca16_csa10_csa_component_fa19_and0 | s_CSAwallace_rca16_csa10_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa20_xor0 = s_CSAwallace_rca16_csa8_csa_component_fa20_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa20_and0 = s_CSAwallace_rca16_csa8_csa_component_fa20_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa20_and1 = s_CSAwallace_rca16_csa10_csa_component_fa20_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa20_or0 = s_CSAwallace_rca16_csa10_csa_component_fa20_and0 | s_CSAwallace_rca16_csa10_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa21_xor0 = s_CSAwallace_rca16_csa6_csa_component_fa21_xor1 ^ s_CSAwallace_rca16_csa8_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa21_and0 = s_CSAwallace_rca16_csa6_csa_component_fa21_xor1 & s_CSAwallace_rca16_csa8_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa10_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa21_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa21_and1 = s_CSAwallace_rca16_csa10_csa_component_fa21_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa21_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa21_or0 = s_CSAwallace_rca16_csa10_csa_component_fa21_and0 | s_CSAwallace_rca16_csa10_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa22_xor0 = ~s_CSAwallace_rca16_csa6_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa22_and1 = s_CSAwallace_rca16_csa10_csa_component_fa22_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa22_or0 = s_CSAwallace_rca16_csa6_csa_component_fa22_xor1 | s_CSAwallace_rca16_csa10_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa23_xor0 = ~s_CSAwallace_rca16_csa6_csa_component_fa23_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa23_xor1 = s_CSAwallace_rca16_csa10_csa_component_fa23_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa23_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa23_and1 = s_CSAwallace_rca16_csa10_csa_component_fa23_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa23_xor1;
  assign s_CSAwallace_rca16_csa10_csa_component_fa23_or0 = s_CSAwallace_rca16_csa6_csa_component_fa23_xor1 | s_CSAwallace_rca16_csa10_csa_component_fa23_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa14_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa13_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa13_and0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa14_and0 = s_CSAwallace_rca16_csa9_csa_component_fa13_or0 & s_CSAwallace_rca16_csa4_csa_component_fa13_and0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa15_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa14_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa15_and0 = s_CSAwallace_rca16_csa9_csa_component_fa14_or0 & s_CSAwallace_rca16_csa4_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_nand_0_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa15_and1 = s_CSAwallace_rca16_csa11_csa_component_fa15_xor0 & s_CSAwallace_rca16_nand_0_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa15_or0 = s_CSAwallace_rca16_csa11_csa_component_fa15_and0 | s_CSAwallace_rca16_csa11_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa16_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa15_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa16_and0 = s_CSAwallace_rca16_csa9_csa_component_fa15_or0 & s_CSAwallace_rca16_csa4_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_nand_1_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa16_and1 = s_CSAwallace_rca16_csa11_csa_component_fa16_xor0 & s_CSAwallace_rca16_nand_1_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa16_or0 = s_CSAwallace_rca16_csa11_csa_component_fa16_and0 | s_CSAwallace_rca16_csa11_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa17_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa16_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa17_and0 = s_CSAwallace_rca16_csa9_csa_component_fa16_or0 & s_CSAwallace_rca16_csa4_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_nand_2_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa17_and1 = s_CSAwallace_rca16_csa11_csa_component_fa17_xor0 & s_CSAwallace_rca16_nand_2_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa17_or0 = s_CSAwallace_rca16_csa11_csa_component_fa17_and0 | s_CSAwallace_rca16_csa11_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa18_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa17_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa18_and0 = s_CSAwallace_rca16_csa9_csa_component_fa17_or0 & s_CSAwallace_rca16_csa4_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_nand_3_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa18_and1 = s_CSAwallace_rca16_csa11_csa_component_fa18_xor0 & s_CSAwallace_rca16_nand_3_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa18_or0 = s_CSAwallace_rca16_csa11_csa_component_fa18_and0 | s_CSAwallace_rca16_csa11_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa19_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa18_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa19_and0 = s_CSAwallace_rca16_csa9_csa_component_fa18_or0 & s_CSAwallace_rca16_csa4_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_nand_4_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa19_and1 = s_CSAwallace_rca16_csa11_csa_component_fa19_xor0 & s_CSAwallace_rca16_nand_4_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa19_or0 = s_CSAwallace_rca16_csa11_csa_component_fa19_and0 | s_CSAwallace_rca16_csa11_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa20_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa19_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa20_and0 = s_CSAwallace_rca16_csa9_csa_component_fa19_or0 & s_CSAwallace_rca16_csa4_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_nand_5_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa20_and1 = s_CSAwallace_rca16_csa11_csa_component_fa20_xor0 & s_CSAwallace_rca16_nand_5_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa20_or0 = s_CSAwallace_rca16_csa11_csa_component_fa20_and0 | s_CSAwallace_rca16_csa11_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa21_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa20_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa21_and0 = s_CSAwallace_rca16_csa9_csa_component_fa20_or0 & s_CSAwallace_rca16_csa4_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_nand_6_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa21_and1 = s_CSAwallace_rca16_csa11_csa_component_fa21_xor0 & s_CSAwallace_rca16_nand_6_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa21_or0 = s_CSAwallace_rca16_csa11_csa_component_fa21_and0 | s_CSAwallace_rca16_csa11_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa22_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa21_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa22_and0 = s_CSAwallace_rca16_csa9_csa_component_fa21_or0 & s_CSAwallace_rca16_csa4_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_nand_7_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa22_and1 = s_CSAwallace_rca16_csa11_csa_component_fa22_xor0 & s_CSAwallace_rca16_nand_7_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa22_or0 = s_CSAwallace_rca16_csa11_csa_component_fa22_and0 | s_CSAwallace_rca16_csa11_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa23_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa22_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa23_and0 = s_CSAwallace_rca16_csa9_csa_component_fa22_or0 & s_CSAwallace_rca16_csa4_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa23_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa23_xor0 ^ s_CSAwallace_rca16_nand_8_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa23_and1 = s_CSAwallace_rca16_csa11_csa_component_fa23_xor0 & s_CSAwallace_rca16_nand_8_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa23_or0 = s_CSAwallace_rca16_csa11_csa_component_fa23_and0 | s_CSAwallace_rca16_csa11_csa_component_fa23_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa24_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa23_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa24_and0 = s_CSAwallace_rca16_csa9_csa_component_fa23_or0 & s_CSAwallace_rca16_csa4_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa24_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa24_xor0 ^ s_CSAwallace_rca16_nand_9_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa24_and1 = s_CSAwallace_rca16_csa11_csa_component_fa24_xor0 & s_CSAwallace_rca16_nand_9_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa24_or0 = s_CSAwallace_rca16_csa11_csa_component_fa24_and0 | s_CSAwallace_rca16_csa11_csa_component_fa24_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa25_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa24_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa25_and0 = s_CSAwallace_rca16_csa9_csa_component_fa24_or0 & s_CSAwallace_rca16_csa4_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa25_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa25_xor0 ^ s_CSAwallace_rca16_nand_10_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa25_and1 = s_CSAwallace_rca16_csa11_csa_component_fa25_xor0 & s_CSAwallace_rca16_nand_10_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa25_or0 = s_CSAwallace_rca16_csa11_csa_component_fa25_and0 | s_CSAwallace_rca16_csa11_csa_component_fa25_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa26_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa25_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa26_and0 = s_CSAwallace_rca16_csa9_csa_component_fa25_or0 & s_CSAwallace_rca16_csa4_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa26_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa26_xor0 ^ s_CSAwallace_rca16_nand_11_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa26_and1 = s_CSAwallace_rca16_csa11_csa_component_fa26_xor0 & s_CSAwallace_rca16_nand_11_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa26_or0 = s_CSAwallace_rca16_csa11_csa_component_fa26_and0 | s_CSAwallace_rca16_csa11_csa_component_fa26_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa27_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa26_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa27_and0 = s_CSAwallace_rca16_csa9_csa_component_fa26_or0 & s_CSAwallace_rca16_csa4_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa27_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa27_xor0 ^ s_CSAwallace_rca16_nand_12_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa27_and1 = s_CSAwallace_rca16_csa11_csa_component_fa27_xor0 & s_CSAwallace_rca16_nand_12_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa27_or0 = s_CSAwallace_rca16_csa11_csa_component_fa27_and0 | s_CSAwallace_rca16_csa11_csa_component_fa27_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa28_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa27_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa27_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa28_and0 = s_CSAwallace_rca16_csa9_csa_component_fa27_or0 & s_CSAwallace_rca16_csa4_csa_component_fa27_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa28_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa28_xor0 ^ s_CSAwallace_rca16_nand_13_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa28_and1 = s_CSAwallace_rca16_csa11_csa_component_fa28_xor0 & s_CSAwallace_rca16_nand_13_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa28_or0 = s_CSAwallace_rca16_csa11_csa_component_fa28_and0 | s_CSAwallace_rca16_csa11_csa_component_fa28_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa29_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa28_or0 ^ s_CSAwallace_rca16_csa4_csa_component_fa28_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa29_and0 = s_CSAwallace_rca16_csa9_csa_component_fa28_or0 & s_CSAwallace_rca16_csa4_csa_component_fa28_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa29_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa29_xor0 ^ s_CSAwallace_rca16_nand_14_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa29_and1 = s_CSAwallace_rca16_csa11_csa_component_fa29_xor0 & s_CSAwallace_rca16_nand_14_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa29_or0 = s_CSAwallace_rca16_csa11_csa_component_fa29_and0 | s_CSAwallace_rca16_csa11_csa_component_fa29_and1;
  assign s_CSAwallace_rca16_csa11_csa_component_fa30_xor0 = ~s_CSAwallace_rca16_csa9_csa_component_fa29_or0;
  assign s_CSAwallace_rca16_csa11_csa_component_fa30_xor1 = s_CSAwallace_rca16_csa11_csa_component_fa30_xor0 ^ s_CSAwallace_rca16_and_15_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa30_and1 = s_CSAwallace_rca16_csa11_csa_component_fa30_xor0 & s_CSAwallace_rca16_and_15_15;
  assign s_CSAwallace_rca16_csa11_csa_component_fa30_or0 = s_CSAwallace_rca16_csa9_csa_component_fa29_or0 | s_CSAwallace_rca16_csa11_csa_component_fa30_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa5_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa5_xor0 ^ s_CSAwallace_rca16_csa10_csa_component_fa4_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa5_and0 = s_CSAwallace_rca16_csa10_csa_component_fa5_xor0 & s_CSAwallace_rca16_csa10_csa_component_fa4_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa6_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa6_xor0 ^ s_CSAwallace_rca16_csa10_csa_component_fa5_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa6_and0 = s_CSAwallace_rca16_csa10_csa_component_fa6_xor0 & s_CSAwallace_rca16_csa10_csa_component_fa5_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa7_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa7_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa6_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa7_and0 = s_CSAwallace_rca16_csa10_csa_component_fa7_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa6_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa8_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa8_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa7_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa8_and0 = s_CSAwallace_rca16_csa10_csa_component_fa8_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa7_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa9_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa9_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa9_and0 = s_CSAwallace_rca16_csa10_csa_component_fa9_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa8_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa10_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa10_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa10_and0 = s_CSAwallace_rca16_csa10_csa_component_fa10_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa9_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa10_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa10_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa9_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa10_and1 = s_CSAwallace_rca16_csa12_csa_component_fa10_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa9_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa10_or0 = s_CSAwallace_rca16_csa12_csa_component_fa10_and0 | s_CSAwallace_rca16_csa12_csa_component_fa10_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa11_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa11_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa11_and0 = s_CSAwallace_rca16_csa10_csa_component_fa11_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa11_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa10_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa11_and1 = s_CSAwallace_rca16_csa12_csa_component_fa11_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa10_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa11_or0 = s_CSAwallace_rca16_csa12_csa_component_fa11_and0 | s_CSAwallace_rca16_csa12_csa_component_fa11_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa12_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa12_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa12_and0 = s_CSAwallace_rca16_csa10_csa_component_fa12_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa12_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa11_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa12_and1 = s_CSAwallace_rca16_csa12_csa_component_fa12_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa11_and0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa12_or0 = s_CSAwallace_rca16_csa12_csa_component_fa12_and0 | s_CSAwallace_rca16_csa12_csa_component_fa12_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa13_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa13_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa13_and0 = s_CSAwallace_rca16_csa10_csa_component_fa13_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa13_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_csa9_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa13_and1 = s_CSAwallace_rca16_csa12_csa_component_fa13_xor0 & s_CSAwallace_rca16_csa9_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa13_or0 = s_CSAwallace_rca16_csa12_csa_component_fa13_and0 | s_CSAwallace_rca16_csa12_csa_component_fa13_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa14_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa14_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa14_and0 = s_CSAwallace_rca16_csa10_csa_component_fa14_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa14_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa14_xor0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa14_and1 = s_CSAwallace_rca16_csa12_csa_component_fa14_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa14_xor0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa14_or0 = s_CSAwallace_rca16_csa12_csa_component_fa14_and0 | s_CSAwallace_rca16_csa12_csa_component_fa14_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa15_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa15_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa15_and0 = s_CSAwallace_rca16_csa10_csa_component_fa15_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa15_and1 = s_CSAwallace_rca16_csa12_csa_component_fa15_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa15_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa15_or0 = s_CSAwallace_rca16_csa12_csa_component_fa15_and0 | s_CSAwallace_rca16_csa12_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa16_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa16_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa16_and0 = s_CSAwallace_rca16_csa10_csa_component_fa16_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa16_and1 = s_CSAwallace_rca16_csa12_csa_component_fa16_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa16_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa16_or0 = s_CSAwallace_rca16_csa12_csa_component_fa16_and0 | s_CSAwallace_rca16_csa12_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa17_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa17_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa17_and0 = s_CSAwallace_rca16_csa10_csa_component_fa17_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa17_and1 = s_CSAwallace_rca16_csa12_csa_component_fa17_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa17_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa17_or0 = s_CSAwallace_rca16_csa12_csa_component_fa17_and0 | s_CSAwallace_rca16_csa12_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa18_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa18_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa18_and0 = s_CSAwallace_rca16_csa10_csa_component_fa18_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa18_and1 = s_CSAwallace_rca16_csa12_csa_component_fa18_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa18_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa18_or0 = s_CSAwallace_rca16_csa12_csa_component_fa18_and0 | s_CSAwallace_rca16_csa12_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa19_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa19_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa19_and0 = s_CSAwallace_rca16_csa10_csa_component_fa19_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa19_and1 = s_CSAwallace_rca16_csa12_csa_component_fa19_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa19_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa19_or0 = s_CSAwallace_rca16_csa12_csa_component_fa19_and0 | s_CSAwallace_rca16_csa12_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa20_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa20_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa20_and0 = s_CSAwallace_rca16_csa10_csa_component_fa20_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa20_and1 = s_CSAwallace_rca16_csa12_csa_component_fa20_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa20_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa20_or0 = s_CSAwallace_rca16_csa12_csa_component_fa20_and0 | s_CSAwallace_rca16_csa12_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa21_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa21_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa21_and0 = s_CSAwallace_rca16_csa10_csa_component_fa21_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa21_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa21_and1 = s_CSAwallace_rca16_csa12_csa_component_fa21_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa21_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa21_or0 = s_CSAwallace_rca16_csa12_csa_component_fa21_and0 | s_CSAwallace_rca16_csa12_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa22_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa22_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa22_and0 = s_CSAwallace_rca16_csa10_csa_component_fa22_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa22_and1 = s_CSAwallace_rca16_csa12_csa_component_fa22_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa22_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa22_or0 = s_CSAwallace_rca16_csa12_csa_component_fa22_and0 | s_CSAwallace_rca16_csa12_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa23_xor0 = s_CSAwallace_rca16_csa10_csa_component_fa23_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa23_and0 = s_CSAwallace_rca16_csa10_csa_component_fa23_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa23_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa23_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa23_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa23_and1 = s_CSAwallace_rca16_csa12_csa_component_fa23_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa23_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa23_or0 = s_CSAwallace_rca16_csa12_csa_component_fa23_and0 | s_CSAwallace_rca16_csa12_csa_component_fa23_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa24_xor0 = s_CSAwallace_rca16_csa9_csa_component_fa24_xor1 ^ s_CSAwallace_rca16_csa10_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa24_and0 = s_CSAwallace_rca16_csa9_csa_component_fa24_xor1 & s_CSAwallace_rca16_csa10_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa12_csa_component_fa24_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa24_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa24_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa24_and1 = s_CSAwallace_rca16_csa12_csa_component_fa24_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa24_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa24_or0 = s_CSAwallace_rca16_csa12_csa_component_fa24_and0 | s_CSAwallace_rca16_csa12_csa_component_fa24_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa25_xor0 = ~s_CSAwallace_rca16_csa9_csa_component_fa25_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa25_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa25_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa25_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa25_and1 = s_CSAwallace_rca16_csa12_csa_component_fa25_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa25_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa25_or0 = s_CSAwallace_rca16_csa9_csa_component_fa25_xor1 | s_CSAwallace_rca16_csa12_csa_component_fa25_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa26_xor0 = ~s_CSAwallace_rca16_csa9_csa_component_fa26_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa26_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa26_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa26_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa26_and1 = s_CSAwallace_rca16_csa12_csa_component_fa26_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa26_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa26_or0 = s_CSAwallace_rca16_csa9_csa_component_fa26_xor1 | s_CSAwallace_rca16_csa12_csa_component_fa26_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa27_xor0 = ~s_CSAwallace_rca16_csa9_csa_component_fa27_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa27_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa27_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa27_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa27_and1 = s_CSAwallace_rca16_csa12_csa_component_fa27_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa27_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa27_or0 = s_CSAwallace_rca16_csa9_csa_component_fa27_xor1 | s_CSAwallace_rca16_csa12_csa_component_fa27_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa28_xor0 = ~s_CSAwallace_rca16_csa9_csa_component_fa28_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa28_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa28_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa28_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa28_and1 = s_CSAwallace_rca16_csa12_csa_component_fa28_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa28_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa28_or0 = s_CSAwallace_rca16_csa9_csa_component_fa28_xor1 | s_CSAwallace_rca16_csa12_csa_component_fa28_and1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa29_xor0 = ~s_CSAwallace_rca16_csa9_csa_component_fa29_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa29_xor1 = s_CSAwallace_rca16_csa12_csa_component_fa29_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa29_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa29_and1 = s_CSAwallace_rca16_csa12_csa_component_fa29_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa29_xor1;
  assign s_CSAwallace_rca16_csa12_csa_component_fa29_or0 = s_CSAwallace_rca16_csa9_csa_component_fa29_xor1 | s_CSAwallace_rca16_csa12_csa_component_fa29_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa6_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa6_xor0 ^ s_CSAwallace_rca16_csa12_csa_component_fa5_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa6_and0 = s_CSAwallace_rca16_csa12_csa_component_fa6_xor0 & s_CSAwallace_rca16_csa12_csa_component_fa5_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa7_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa7_xor0 ^ s_CSAwallace_rca16_csa12_csa_component_fa6_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa7_and0 = s_CSAwallace_rca16_csa12_csa_component_fa7_xor0 & s_CSAwallace_rca16_csa12_csa_component_fa6_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa8_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa8_xor0 ^ s_CSAwallace_rca16_csa12_csa_component_fa7_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa8_and0 = s_CSAwallace_rca16_csa12_csa_component_fa8_xor0 & s_CSAwallace_rca16_csa12_csa_component_fa7_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa9_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa9_xor0 ^ s_CSAwallace_rca16_csa12_csa_component_fa8_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa9_and0 = s_CSAwallace_rca16_csa12_csa_component_fa9_xor0 & s_CSAwallace_rca16_csa12_csa_component_fa8_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa10_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa10_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa9_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa10_and0 = s_CSAwallace_rca16_csa12_csa_component_fa10_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa9_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa11_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa11_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa11_and0 = s_CSAwallace_rca16_csa12_csa_component_fa11_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa10_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa12_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa12_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa12_and0 = s_CSAwallace_rca16_csa12_csa_component_fa12_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa11_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa13_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa13_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa13_and0 = s_CSAwallace_rca16_csa12_csa_component_fa13_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa12_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa14_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa14_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa14_and0 = s_CSAwallace_rca16_csa12_csa_component_fa14_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa13_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa15_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa15_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa15_and0 = s_CSAwallace_rca16_csa12_csa_component_fa15_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa14_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa15_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa15_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa14_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa15_and1 = s_CSAwallace_rca16_csa13_csa_component_fa15_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa14_and0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa15_or0 = s_CSAwallace_rca16_csa13_csa_component_fa15_and0 | s_CSAwallace_rca16_csa13_csa_component_fa15_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa16_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa16_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa16_and0 = s_CSAwallace_rca16_csa12_csa_component_fa16_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa16_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa16_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa16_and1 = s_CSAwallace_rca16_csa13_csa_component_fa16_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa16_or0 = s_CSAwallace_rca16_csa13_csa_component_fa16_and0 | s_CSAwallace_rca16_csa13_csa_component_fa16_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa17_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa17_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa17_and0 = s_CSAwallace_rca16_csa12_csa_component_fa17_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa17_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa17_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa17_and1 = s_CSAwallace_rca16_csa13_csa_component_fa17_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa17_or0 = s_CSAwallace_rca16_csa13_csa_component_fa17_and0 | s_CSAwallace_rca16_csa13_csa_component_fa17_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa18_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa18_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa18_and0 = s_CSAwallace_rca16_csa12_csa_component_fa18_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa18_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa18_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa18_and1 = s_CSAwallace_rca16_csa13_csa_component_fa18_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa18_or0 = s_CSAwallace_rca16_csa13_csa_component_fa18_and0 | s_CSAwallace_rca16_csa13_csa_component_fa18_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa19_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa19_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa19_and0 = s_CSAwallace_rca16_csa12_csa_component_fa19_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa19_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa19_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa19_and1 = s_CSAwallace_rca16_csa13_csa_component_fa19_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa19_or0 = s_CSAwallace_rca16_csa13_csa_component_fa19_and0 | s_CSAwallace_rca16_csa13_csa_component_fa19_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa20_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa20_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa20_and0 = s_CSAwallace_rca16_csa12_csa_component_fa20_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa20_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa20_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa20_and1 = s_CSAwallace_rca16_csa13_csa_component_fa20_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa20_or0 = s_CSAwallace_rca16_csa13_csa_component_fa20_and0 | s_CSAwallace_rca16_csa13_csa_component_fa20_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa21_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa21_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa21_and0 = s_CSAwallace_rca16_csa12_csa_component_fa21_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa21_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa21_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa21_and1 = s_CSAwallace_rca16_csa13_csa_component_fa21_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa21_or0 = s_CSAwallace_rca16_csa13_csa_component_fa21_and0 | s_CSAwallace_rca16_csa13_csa_component_fa21_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa22_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa22_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa22_and0 = s_CSAwallace_rca16_csa12_csa_component_fa22_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa22_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa22_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa22_and1 = s_CSAwallace_rca16_csa13_csa_component_fa22_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa22_or0 = s_CSAwallace_rca16_csa13_csa_component_fa22_and0 | s_CSAwallace_rca16_csa13_csa_component_fa22_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa23_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa23_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa23_and0 = s_CSAwallace_rca16_csa12_csa_component_fa23_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa23_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa23_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa23_and1 = s_CSAwallace_rca16_csa13_csa_component_fa23_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa23_or0 = s_CSAwallace_rca16_csa13_csa_component_fa23_and0 | s_CSAwallace_rca16_csa13_csa_component_fa23_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa24_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa24_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa24_and0 = s_CSAwallace_rca16_csa12_csa_component_fa24_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa24_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa24_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa24_and1 = s_CSAwallace_rca16_csa13_csa_component_fa24_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa24_or0 = s_CSAwallace_rca16_csa13_csa_component_fa24_and0 | s_CSAwallace_rca16_csa13_csa_component_fa24_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa25_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa25_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa25_and0 = s_CSAwallace_rca16_csa12_csa_component_fa25_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa25_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa25_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa25_and1 = s_CSAwallace_rca16_csa13_csa_component_fa25_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa25_or0 = s_CSAwallace_rca16_csa13_csa_component_fa25_and0 | s_CSAwallace_rca16_csa13_csa_component_fa25_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa26_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa26_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa26_and0 = s_CSAwallace_rca16_csa12_csa_component_fa26_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa26_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa26_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa26_and1 = s_CSAwallace_rca16_csa13_csa_component_fa26_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa26_or0 = s_CSAwallace_rca16_csa13_csa_component_fa26_and0 | s_CSAwallace_rca16_csa13_csa_component_fa26_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa27_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa27_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa27_and0 = s_CSAwallace_rca16_csa12_csa_component_fa27_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa27_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa27_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa27_and1 = s_CSAwallace_rca16_csa13_csa_component_fa27_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa27_or0 = s_CSAwallace_rca16_csa13_csa_component_fa27_and0 | s_CSAwallace_rca16_csa13_csa_component_fa27_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa28_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa28_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa27_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa28_and0 = s_CSAwallace_rca16_csa12_csa_component_fa28_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa27_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa28_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa28_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa27_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa28_and1 = s_CSAwallace_rca16_csa13_csa_component_fa28_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa27_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa28_or0 = s_CSAwallace_rca16_csa13_csa_component_fa28_and0 | s_CSAwallace_rca16_csa13_csa_component_fa28_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa29_xor0 = s_CSAwallace_rca16_csa12_csa_component_fa29_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa28_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa29_and0 = s_CSAwallace_rca16_csa12_csa_component_fa29_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa28_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa29_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa29_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa28_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa29_and1 = s_CSAwallace_rca16_csa13_csa_component_fa29_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa28_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa29_or0 = s_CSAwallace_rca16_csa13_csa_component_fa29_and0 | s_CSAwallace_rca16_csa13_csa_component_fa29_and1;
  assign s_CSAwallace_rca16_csa13_csa_component_fa30_xor0 = s_CSAwallace_rca16_csa11_csa_component_fa30_xor1 ^ s_CSAwallace_rca16_csa12_csa_component_fa29_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa30_and0 = s_CSAwallace_rca16_csa11_csa_component_fa30_xor1 & s_CSAwallace_rca16_csa12_csa_component_fa29_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa30_xor1 = s_CSAwallace_rca16_csa13_csa_component_fa30_xor0 ^ s_CSAwallace_rca16_csa11_csa_component_fa29_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa30_and1 = s_CSAwallace_rca16_csa13_csa_component_fa30_xor0 & s_CSAwallace_rca16_csa11_csa_component_fa29_or0;
  assign s_CSAwallace_rca16_csa13_csa_component_fa30_or0 = s_CSAwallace_rca16_csa13_csa_component_fa30_and0 | s_CSAwallace_rca16_csa13_csa_component_fa30_and1;
  assign s_CSAwallace_rca16_u_rca32_fa7_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa7_xor0 ^ s_CSAwallace_rca16_csa13_csa_component_fa6_and0;
  assign s_CSAwallace_rca16_u_rca32_fa7_and0 = s_CSAwallace_rca16_csa13_csa_component_fa7_xor0 & s_CSAwallace_rca16_csa13_csa_component_fa6_and0;
  assign s_CSAwallace_rca16_u_rca32_fa8_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa8_xor0 ^ s_CSAwallace_rca16_csa13_csa_component_fa7_and0;
  assign s_CSAwallace_rca16_u_rca32_fa8_and0 = s_CSAwallace_rca16_csa13_csa_component_fa8_xor0 & s_CSAwallace_rca16_csa13_csa_component_fa7_and0;
  assign s_CSAwallace_rca16_u_rca32_fa8_xor1 = s_CSAwallace_rca16_u_rca32_fa8_xor0 ^ s_CSAwallace_rca16_u_rca32_fa7_and0;
  assign s_CSAwallace_rca16_u_rca32_fa8_and1 = s_CSAwallace_rca16_u_rca32_fa8_xor0 & s_CSAwallace_rca16_u_rca32_fa7_and0;
  assign s_CSAwallace_rca16_u_rca32_fa8_or0 = s_CSAwallace_rca16_u_rca32_fa8_and0 | s_CSAwallace_rca16_u_rca32_fa8_and1;
  assign s_CSAwallace_rca16_u_rca32_fa9_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa9_xor0 ^ s_CSAwallace_rca16_csa13_csa_component_fa8_and0;
  assign s_CSAwallace_rca16_u_rca32_fa9_and0 = s_CSAwallace_rca16_csa13_csa_component_fa9_xor0 & s_CSAwallace_rca16_csa13_csa_component_fa8_and0;
  assign s_CSAwallace_rca16_u_rca32_fa9_xor1 = s_CSAwallace_rca16_u_rca32_fa9_xor0 ^ s_CSAwallace_rca16_u_rca32_fa8_or0;
  assign s_CSAwallace_rca16_u_rca32_fa9_and1 = s_CSAwallace_rca16_u_rca32_fa9_xor0 & s_CSAwallace_rca16_u_rca32_fa8_or0;
  assign s_CSAwallace_rca16_u_rca32_fa9_or0 = s_CSAwallace_rca16_u_rca32_fa9_and0 | s_CSAwallace_rca16_u_rca32_fa9_and1;
  assign s_CSAwallace_rca16_u_rca32_fa10_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa10_xor0 ^ s_CSAwallace_rca16_csa13_csa_component_fa9_and0;
  assign s_CSAwallace_rca16_u_rca32_fa10_and0 = s_CSAwallace_rca16_csa13_csa_component_fa10_xor0 & s_CSAwallace_rca16_csa13_csa_component_fa9_and0;
  assign s_CSAwallace_rca16_u_rca32_fa10_xor1 = s_CSAwallace_rca16_u_rca32_fa10_xor0 ^ s_CSAwallace_rca16_u_rca32_fa9_or0;
  assign s_CSAwallace_rca16_u_rca32_fa10_and1 = s_CSAwallace_rca16_u_rca32_fa10_xor0 & s_CSAwallace_rca16_u_rca32_fa9_or0;
  assign s_CSAwallace_rca16_u_rca32_fa10_or0 = s_CSAwallace_rca16_u_rca32_fa10_and0 | s_CSAwallace_rca16_u_rca32_fa10_and1;
  assign s_CSAwallace_rca16_u_rca32_fa11_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa11_xor0 ^ s_CSAwallace_rca16_csa13_csa_component_fa10_and0;
  assign s_CSAwallace_rca16_u_rca32_fa11_and0 = s_CSAwallace_rca16_csa13_csa_component_fa11_xor0 & s_CSAwallace_rca16_csa13_csa_component_fa10_and0;
  assign s_CSAwallace_rca16_u_rca32_fa11_xor1 = s_CSAwallace_rca16_u_rca32_fa11_xor0 ^ s_CSAwallace_rca16_u_rca32_fa10_or0;
  assign s_CSAwallace_rca16_u_rca32_fa11_and1 = s_CSAwallace_rca16_u_rca32_fa11_xor0 & s_CSAwallace_rca16_u_rca32_fa10_or0;
  assign s_CSAwallace_rca16_u_rca32_fa11_or0 = s_CSAwallace_rca16_u_rca32_fa11_and0 | s_CSAwallace_rca16_u_rca32_fa11_and1;
  assign s_CSAwallace_rca16_u_rca32_fa12_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa12_xor0 ^ s_CSAwallace_rca16_csa13_csa_component_fa11_and0;
  assign s_CSAwallace_rca16_u_rca32_fa12_and0 = s_CSAwallace_rca16_csa13_csa_component_fa12_xor0 & s_CSAwallace_rca16_csa13_csa_component_fa11_and0;
  assign s_CSAwallace_rca16_u_rca32_fa12_xor1 = s_CSAwallace_rca16_u_rca32_fa12_xor0 ^ s_CSAwallace_rca16_u_rca32_fa11_or0;
  assign s_CSAwallace_rca16_u_rca32_fa12_and1 = s_CSAwallace_rca16_u_rca32_fa12_xor0 & s_CSAwallace_rca16_u_rca32_fa11_or0;
  assign s_CSAwallace_rca16_u_rca32_fa12_or0 = s_CSAwallace_rca16_u_rca32_fa12_and0 | s_CSAwallace_rca16_u_rca32_fa12_and1;
  assign s_CSAwallace_rca16_u_rca32_fa13_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa13_xor0 ^ s_CSAwallace_rca16_csa13_csa_component_fa12_and0;
  assign s_CSAwallace_rca16_u_rca32_fa13_and0 = s_CSAwallace_rca16_csa13_csa_component_fa13_xor0 & s_CSAwallace_rca16_csa13_csa_component_fa12_and0;
  assign s_CSAwallace_rca16_u_rca32_fa13_xor1 = s_CSAwallace_rca16_u_rca32_fa13_xor0 ^ s_CSAwallace_rca16_u_rca32_fa12_or0;
  assign s_CSAwallace_rca16_u_rca32_fa13_and1 = s_CSAwallace_rca16_u_rca32_fa13_xor0 & s_CSAwallace_rca16_u_rca32_fa12_or0;
  assign s_CSAwallace_rca16_u_rca32_fa13_or0 = s_CSAwallace_rca16_u_rca32_fa13_and0 | s_CSAwallace_rca16_u_rca32_fa13_and1;
  assign s_CSAwallace_rca16_u_rca32_fa14_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa14_xor0 ^ s_CSAwallace_rca16_csa13_csa_component_fa13_and0;
  assign s_CSAwallace_rca16_u_rca32_fa14_and0 = s_CSAwallace_rca16_csa13_csa_component_fa14_xor0 & s_CSAwallace_rca16_csa13_csa_component_fa13_and0;
  assign s_CSAwallace_rca16_u_rca32_fa14_xor1 = s_CSAwallace_rca16_u_rca32_fa14_xor0 ^ s_CSAwallace_rca16_u_rca32_fa13_or0;
  assign s_CSAwallace_rca16_u_rca32_fa14_and1 = s_CSAwallace_rca16_u_rca32_fa14_xor0 & s_CSAwallace_rca16_u_rca32_fa13_or0;
  assign s_CSAwallace_rca16_u_rca32_fa14_or0 = s_CSAwallace_rca16_u_rca32_fa14_and0 | s_CSAwallace_rca16_u_rca32_fa14_and1;
  assign s_CSAwallace_rca16_u_rca32_fa15_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa15_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa14_and0;
  assign s_CSAwallace_rca16_u_rca32_fa15_and0 = s_CSAwallace_rca16_csa13_csa_component_fa15_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa14_and0;
  assign s_CSAwallace_rca16_u_rca32_fa15_xor1 = s_CSAwallace_rca16_u_rca32_fa15_xor0 ^ s_CSAwallace_rca16_u_rca32_fa14_or0;
  assign s_CSAwallace_rca16_u_rca32_fa15_and1 = s_CSAwallace_rca16_u_rca32_fa15_xor0 & s_CSAwallace_rca16_u_rca32_fa14_or0;
  assign s_CSAwallace_rca16_u_rca32_fa15_or0 = s_CSAwallace_rca16_u_rca32_fa15_and0 | s_CSAwallace_rca16_u_rca32_fa15_and1;
  assign s_CSAwallace_rca16_u_rca32_fa16_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa16_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_u_rca32_fa16_and0 = s_CSAwallace_rca16_csa13_csa_component_fa16_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa15_or0;
  assign s_CSAwallace_rca16_u_rca32_fa16_xor1 = s_CSAwallace_rca16_u_rca32_fa16_xor0 ^ s_CSAwallace_rca16_u_rca32_fa15_or0;
  assign s_CSAwallace_rca16_u_rca32_fa16_and1 = s_CSAwallace_rca16_u_rca32_fa16_xor0 & s_CSAwallace_rca16_u_rca32_fa15_or0;
  assign s_CSAwallace_rca16_u_rca32_fa16_or0 = s_CSAwallace_rca16_u_rca32_fa16_and0 | s_CSAwallace_rca16_u_rca32_fa16_and1;
  assign s_CSAwallace_rca16_u_rca32_fa17_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa17_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_u_rca32_fa17_and0 = s_CSAwallace_rca16_csa13_csa_component_fa17_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa16_or0;
  assign s_CSAwallace_rca16_u_rca32_fa17_xor1 = s_CSAwallace_rca16_u_rca32_fa17_xor0 ^ s_CSAwallace_rca16_u_rca32_fa16_or0;
  assign s_CSAwallace_rca16_u_rca32_fa17_and1 = s_CSAwallace_rca16_u_rca32_fa17_xor0 & s_CSAwallace_rca16_u_rca32_fa16_or0;
  assign s_CSAwallace_rca16_u_rca32_fa17_or0 = s_CSAwallace_rca16_u_rca32_fa17_and0 | s_CSAwallace_rca16_u_rca32_fa17_and1;
  assign s_CSAwallace_rca16_u_rca32_fa18_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa18_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_u_rca32_fa18_and0 = s_CSAwallace_rca16_csa13_csa_component_fa18_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa17_or0;
  assign s_CSAwallace_rca16_u_rca32_fa18_xor1 = s_CSAwallace_rca16_u_rca32_fa18_xor0 ^ s_CSAwallace_rca16_u_rca32_fa17_or0;
  assign s_CSAwallace_rca16_u_rca32_fa18_and1 = s_CSAwallace_rca16_u_rca32_fa18_xor0 & s_CSAwallace_rca16_u_rca32_fa17_or0;
  assign s_CSAwallace_rca16_u_rca32_fa18_or0 = s_CSAwallace_rca16_u_rca32_fa18_and0 | s_CSAwallace_rca16_u_rca32_fa18_and1;
  assign s_CSAwallace_rca16_u_rca32_fa19_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa19_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_u_rca32_fa19_and0 = s_CSAwallace_rca16_csa13_csa_component_fa19_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa18_or0;
  assign s_CSAwallace_rca16_u_rca32_fa19_xor1 = s_CSAwallace_rca16_u_rca32_fa19_xor0 ^ s_CSAwallace_rca16_u_rca32_fa18_or0;
  assign s_CSAwallace_rca16_u_rca32_fa19_and1 = s_CSAwallace_rca16_u_rca32_fa19_xor0 & s_CSAwallace_rca16_u_rca32_fa18_or0;
  assign s_CSAwallace_rca16_u_rca32_fa19_or0 = s_CSAwallace_rca16_u_rca32_fa19_and0 | s_CSAwallace_rca16_u_rca32_fa19_and1;
  assign s_CSAwallace_rca16_u_rca32_fa20_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa20_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_u_rca32_fa20_and0 = s_CSAwallace_rca16_csa13_csa_component_fa20_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa19_or0;
  assign s_CSAwallace_rca16_u_rca32_fa20_xor1 = s_CSAwallace_rca16_u_rca32_fa20_xor0 ^ s_CSAwallace_rca16_u_rca32_fa19_or0;
  assign s_CSAwallace_rca16_u_rca32_fa20_and1 = s_CSAwallace_rca16_u_rca32_fa20_xor0 & s_CSAwallace_rca16_u_rca32_fa19_or0;
  assign s_CSAwallace_rca16_u_rca32_fa20_or0 = s_CSAwallace_rca16_u_rca32_fa20_and0 | s_CSAwallace_rca16_u_rca32_fa20_and1;
  assign s_CSAwallace_rca16_u_rca32_fa21_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa21_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_u_rca32_fa21_and0 = s_CSAwallace_rca16_csa13_csa_component_fa21_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa20_or0;
  assign s_CSAwallace_rca16_u_rca32_fa21_xor1 = s_CSAwallace_rca16_u_rca32_fa21_xor0 ^ s_CSAwallace_rca16_u_rca32_fa20_or0;
  assign s_CSAwallace_rca16_u_rca32_fa21_and1 = s_CSAwallace_rca16_u_rca32_fa21_xor0 & s_CSAwallace_rca16_u_rca32_fa20_or0;
  assign s_CSAwallace_rca16_u_rca32_fa21_or0 = s_CSAwallace_rca16_u_rca32_fa21_and0 | s_CSAwallace_rca16_u_rca32_fa21_and1;
  assign s_CSAwallace_rca16_u_rca32_fa22_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa22_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_u_rca32_fa22_and0 = s_CSAwallace_rca16_csa13_csa_component_fa22_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa21_or0;
  assign s_CSAwallace_rca16_u_rca32_fa22_xor1 = s_CSAwallace_rca16_u_rca32_fa22_xor0 ^ s_CSAwallace_rca16_u_rca32_fa21_or0;
  assign s_CSAwallace_rca16_u_rca32_fa22_and1 = s_CSAwallace_rca16_u_rca32_fa22_xor0 & s_CSAwallace_rca16_u_rca32_fa21_or0;
  assign s_CSAwallace_rca16_u_rca32_fa22_or0 = s_CSAwallace_rca16_u_rca32_fa22_and0 | s_CSAwallace_rca16_u_rca32_fa22_and1;
  assign s_CSAwallace_rca16_u_rca32_fa23_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa23_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_u_rca32_fa23_and0 = s_CSAwallace_rca16_csa13_csa_component_fa23_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa22_or0;
  assign s_CSAwallace_rca16_u_rca32_fa23_xor1 = s_CSAwallace_rca16_u_rca32_fa23_xor0 ^ s_CSAwallace_rca16_u_rca32_fa22_or0;
  assign s_CSAwallace_rca16_u_rca32_fa23_and1 = s_CSAwallace_rca16_u_rca32_fa23_xor0 & s_CSAwallace_rca16_u_rca32_fa22_or0;
  assign s_CSAwallace_rca16_u_rca32_fa23_or0 = s_CSAwallace_rca16_u_rca32_fa23_and0 | s_CSAwallace_rca16_u_rca32_fa23_and1;
  assign s_CSAwallace_rca16_u_rca32_fa24_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa24_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_u_rca32_fa24_and0 = s_CSAwallace_rca16_csa13_csa_component_fa24_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa23_or0;
  assign s_CSAwallace_rca16_u_rca32_fa24_xor1 = s_CSAwallace_rca16_u_rca32_fa24_xor0 ^ s_CSAwallace_rca16_u_rca32_fa23_or0;
  assign s_CSAwallace_rca16_u_rca32_fa24_and1 = s_CSAwallace_rca16_u_rca32_fa24_xor0 & s_CSAwallace_rca16_u_rca32_fa23_or0;
  assign s_CSAwallace_rca16_u_rca32_fa24_or0 = s_CSAwallace_rca16_u_rca32_fa24_and0 | s_CSAwallace_rca16_u_rca32_fa24_and1;
  assign s_CSAwallace_rca16_u_rca32_fa25_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa25_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_u_rca32_fa25_and0 = s_CSAwallace_rca16_csa13_csa_component_fa25_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa24_or0;
  assign s_CSAwallace_rca16_u_rca32_fa25_xor1 = s_CSAwallace_rca16_u_rca32_fa25_xor0 ^ s_CSAwallace_rca16_u_rca32_fa24_or0;
  assign s_CSAwallace_rca16_u_rca32_fa25_and1 = s_CSAwallace_rca16_u_rca32_fa25_xor0 & s_CSAwallace_rca16_u_rca32_fa24_or0;
  assign s_CSAwallace_rca16_u_rca32_fa25_or0 = s_CSAwallace_rca16_u_rca32_fa25_and0 | s_CSAwallace_rca16_u_rca32_fa25_and1;
  assign s_CSAwallace_rca16_u_rca32_fa26_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa26_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_u_rca32_fa26_and0 = s_CSAwallace_rca16_csa13_csa_component_fa26_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa25_or0;
  assign s_CSAwallace_rca16_u_rca32_fa26_xor1 = s_CSAwallace_rca16_u_rca32_fa26_xor0 ^ s_CSAwallace_rca16_u_rca32_fa25_or0;
  assign s_CSAwallace_rca16_u_rca32_fa26_and1 = s_CSAwallace_rca16_u_rca32_fa26_xor0 & s_CSAwallace_rca16_u_rca32_fa25_or0;
  assign s_CSAwallace_rca16_u_rca32_fa26_or0 = s_CSAwallace_rca16_u_rca32_fa26_and0 | s_CSAwallace_rca16_u_rca32_fa26_and1;
  assign s_CSAwallace_rca16_u_rca32_fa27_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa27_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_u_rca32_fa27_and0 = s_CSAwallace_rca16_csa13_csa_component_fa27_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa26_or0;
  assign s_CSAwallace_rca16_u_rca32_fa27_xor1 = s_CSAwallace_rca16_u_rca32_fa27_xor0 ^ s_CSAwallace_rca16_u_rca32_fa26_or0;
  assign s_CSAwallace_rca16_u_rca32_fa27_and1 = s_CSAwallace_rca16_u_rca32_fa27_xor0 & s_CSAwallace_rca16_u_rca32_fa26_or0;
  assign s_CSAwallace_rca16_u_rca32_fa27_or0 = s_CSAwallace_rca16_u_rca32_fa27_and0 | s_CSAwallace_rca16_u_rca32_fa27_and1;
  assign s_CSAwallace_rca16_u_rca32_fa28_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa28_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa27_or0;
  assign s_CSAwallace_rca16_u_rca32_fa28_and0 = s_CSAwallace_rca16_csa13_csa_component_fa28_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa27_or0;
  assign s_CSAwallace_rca16_u_rca32_fa28_xor1 = s_CSAwallace_rca16_u_rca32_fa28_xor0 ^ s_CSAwallace_rca16_u_rca32_fa27_or0;
  assign s_CSAwallace_rca16_u_rca32_fa28_and1 = s_CSAwallace_rca16_u_rca32_fa28_xor0 & s_CSAwallace_rca16_u_rca32_fa27_or0;
  assign s_CSAwallace_rca16_u_rca32_fa28_or0 = s_CSAwallace_rca16_u_rca32_fa28_and0 | s_CSAwallace_rca16_u_rca32_fa28_and1;
  assign s_CSAwallace_rca16_u_rca32_fa29_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa29_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa28_or0;
  assign s_CSAwallace_rca16_u_rca32_fa29_and0 = s_CSAwallace_rca16_csa13_csa_component_fa29_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa28_or0;
  assign s_CSAwallace_rca16_u_rca32_fa29_xor1 = s_CSAwallace_rca16_u_rca32_fa29_xor0 ^ s_CSAwallace_rca16_u_rca32_fa28_or0;
  assign s_CSAwallace_rca16_u_rca32_fa29_and1 = s_CSAwallace_rca16_u_rca32_fa29_xor0 & s_CSAwallace_rca16_u_rca32_fa28_or0;
  assign s_CSAwallace_rca16_u_rca32_fa29_or0 = s_CSAwallace_rca16_u_rca32_fa29_and0 | s_CSAwallace_rca16_u_rca32_fa29_and1;
  assign s_CSAwallace_rca16_u_rca32_fa30_xor0 = s_CSAwallace_rca16_csa13_csa_component_fa30_xor1 ^ s_CSAwallace_rca16_csa13_csa_component_fa29_or0;
  assign s_CSAwallace_rca16_u_rca32_fa30_and0 = s_CSAwallace_rca16_csa13_csa_component_fa30_xor1 & s_CSAwallace_rca16_csa13_csa_component_fa29_or0;
  assign s_CSAwallace_rca16_u_rca32_fa30_xor1 = s_CSAwallace_rca16_u_rca32_fa30_xor0 ^ s_CSAwallace_rca16_u_rca32_fa29_or0;
  assign s_CSAwallace_rca16_u_rca32_fa30_and1 = s_CSAwallace_rca16_u_rca32_fa30_xor0 & s_CSAwallace_rca16_u_rca32_fa29_or0;
  assign s_CSAwallace_rca16_u_rca32_fa30_or0 = s_CSAwallace_rca16_u_rca32_fa30_and0 | s_CSAwallace_rca16_u_rca32_fa30_and1;
  assign s_CSAwallace_rca16_u_rca32_fa31_xor0 = s_CSAwallace_rca16_csa11_csa_component_fa30_or0 ^ s_CSAwallace_rca16_csa13_csa_component_fa30_or0;
  assign s_CSAwallace_rca16_u_rca32_fa31_and0 = s_CSAwallace_rca16_csa11_csa_component_fa30_or0 & s_CSAwallace_rca16_csa13_csa_component_fa30_or0;
  assign s_CSAwallace_rca16_u_rca32_fa31_xor1 = s_CSAwallace_rca16_u_rca32_fa31_xor0 ^ s_CSAwallace_rca16_u_rca32_fa30_or0;
  assign s_CSAwallace_rca16_u_rca32_fa31_and1 = s_CSAwallace_rca16_u_rca32_fa31_xor0 & s_CSAwallace_rca16_u_rca32_fa30_or0;
  assign s_CSAwallace_rca16_u_rca32_fa31_or0 = s_CSAwallace_rca16_u_rca32_fa31_and0 | s_CSAwallace_rca16_u_rca32_fa31_and1;
  assign s_CSAwallace_rca16_xor0 = ~s_CSAwallace_rca16_u_rca32_fa31_xor1;

  assign s_CSAwallace_rca16_out[0] = s_CSAwallace_rca16_and_0_0;
  assign s_CSAwallace_rca16_out[1] = s_CSAwallace_rca16_csa0_csa_component_fa1_xor0;
  assign s_CSAwallace_rca16_out[2] = s_CSAwallace_rca16_csa5_csa_component_fa2_xor0;
  assign s_CSAwallace_rca16_out[3] = s_CSAwallace_rca16_csa8_csa_component_fa3_xor0;
  assign s_CSAwallace_rca16_out[4] = s_CSAwallace_rca16_csa10_csa_component_fa4_xor0;
  assign s_CSAwallace_rca16_out[5] = s_CSAwallace_rca16_csa12_csa_component_fa5_xor0;
  assign s_CSAwallace_rca16_out[6] = s_CSAwallace_rca16_csa13_csa_component_fa6_xor0;
  assign s_CSAwallace_rca16_out[7] = s_CSAwallace_rca16_u_rca32_fa7_xor0;
  assign s_CSAwallace_rca16_out[8] = s_CSAwallace_rca16_u_rca32_fa8_xor1;
  assign s_CSAwallace_rca16_out[9] = s_CSAwallace_rca16_u_rca32_fa9_xor1;
  assign s_CSAwallace_rca16_out[10] = s_CSAwallace_rca16_u_rca32_fa10_xor1;
  assign s_CSAwallace_rca16_out[11] = s_CSAwallace_rca16_u_rca32_fa11_xor1;
  assign s_CSAwallace_rca16_out[12] = s_CSAwallace_rca16_u_rca32_fa12_xor1;
  assign s_CSAwallace_rca16_out[13] = s_CSAwallace_rca16_u_rca32_fa13_xor1;
  assign s_CSAwallace_rca16_out[14] = s_CSAwallace_rca16_u_rca32_fa14_xor1;
  assign s_CSAwallace_rca16_out[15] = s_CSAwallace_rca16_u_rca32_fa15_xor1;
  assign s_CSAwallace_rca16_out[16] = s_CSAwallace_rca16_u_rca32_fa16_xor1;
  assign s_CSAwallace_rca16_out[17] = s_CSAwallace_rca16_u_rca32_fa17_xor1;
  assign s_CSAwallace_rca16_out[18] = s_CSAwallace_rca16_u_rca32_fa18_xor1;
  assign s_CSAwallace_rca16_out[19] = s_CSAwallace_rca16_u_rca32_fa19_xor1;
  assign s_CSAwallace_rca16_out[20] = s_CSAwallace_rca16_u_rca32_fa20_xor1;
  assign s_CSAwallace_rca16_out[21] = s_CSAwallace_rca16_u_rca32_fa21_xor1;
  assign s_CSAwallace_rca16_out[22] = s_CSAwallace_rca16_u_rca32_fa22_xor1;
  assign s_CSAwallace_rca16_out[23] = s_CSAwallace_rca16_u_rca32_fa23_xor1;
  assign s_CSAwallace_rca16_out[24] = s_CSAwallace_rca16_u_rca32_fa24_xor1;
  assign s_CSAwallace_rca16_out[25] = s_CSAwallace_rca16_u_rca32_fa25_xor1;
  assign s_CSAwallace_rca16_out[26] = s_CSAwallace_rca16_u_rca32_fa26_xor1;
  assign s_CSAwallace_rca16_out[27] = s_CSAwallace_rca16_u_rca32_fa27_xor1;
  assign s_CSAwallace_rca16_out[28] = s_CSAwallace_rca16_u_rca32_fa28_xor1;
  assign s_CSAwallace_rca16_out[29] = s_CSAwallace_rca16_u_rca32_fa29_xor1;
  assign s_CSAwallace_rca16_out[30] = s_CSAwallace_rca16_u_rca32_fa30_xor1;
  assign s_CSAwallace_rca16_out[31] = s_CSAwallace_rca16_xor0;
endmodule