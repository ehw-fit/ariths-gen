module not_gate(input a, output not_gate);
  assign not_gate = ~a;
endmodule