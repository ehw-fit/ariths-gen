module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(.a(a[0]), .b(b[0]), .out(pg_logic_or0));
  and_gate and_gate_pg_logic_and0(.a(a[0]), .b(b[0]), .out(pg_logic_and0));
  xor_gate xor_gate_pg_logic_xor0(.a(a[0]), .b(b[0]), .out(pg_logic_xor0));
endmodule

module u_cla30(input [29:0] a, input [29:0] b, output [30:0] u_cla30_out);
  wire [0:0] u_cla30_pg_logic0_or0;
  wire [0:0] u_cla30_pg_logic0_and0;
  wire [0:0] u_cla30_pg_logic0_xor0;
  wire [0:0] u_cla30_pg_logic1_or0;
  wire [0:0] u_cla30_pg_logic1_and0;
  wire [0:0] u_cla30_pg_logic1_xor0;
  wire [0:0] u_cla30_xor1;
  wire [0:0] u_cla30_and0;
  wire [0:0] u_cla30_or0;
  wire [0:0] u_cla30_pg_logic2_or0;
  wire [0:0] u_cla30_pg_logic2_and0;
  wire [0:0] u_cla30_pg_logic2_xor0;
  wire [0:0] u_cla30_xor2;
  wire [0:0] u_cla30_and1;
  wire [0:0] u_cla30_and2;
  wire [0:0] u_cla30_and3;
  wire [0:0] u_cla30_and4;
  wire [0:0] u_cla30_or1;
  wire [0:0] u_cla30_or2;
  wire [0:0] u_cla30_pg_logic3_or0;
  wire [0:0] u_cla30_pg_logic3_and0;
  wire [0:0] u_cla30_pg_logic3_xor0;
  wire [0:0] u_cla30_xor3;
  wire [0:0] u_cla30_and5;
  wire [0:0] u_cla30_and6;
  wire [0:0] u_cla30_and7;
  wire [0:0] u_cla30_and8;
  wire [0:0] u_cla30_and9;
  wire [0:0] u_cla30_and10;
  wire [0:0] u_cla30_and11;
  wire [0:0] u_cla30_or3;
  wire [0:0] u_cla30_or4;
  wire [0:0] u_cla30_or5;
  wire [0:0] u_cla30_pg_logic4_or0;
  wire [0:0] u_cla30_pg_logic4_and0;
  wire [0:0] u_cla30_pg_logic4_xor0;
  wire [0:0] u_cla30_xor4;
  wire [0:0] u_cla30_and12;
  wire [0:0] u_cla30_or6;
  wire [0:0] u_cla30_pg_logic5_or0;
  wire [0:0] u_cla30_pg_logic5_and0;
  wire [0:0] u_cla30_pg_logic5_xor0;
  wire [0:0] u_cla30_xor5;
  wire [0:0] u_cla30_and13;
  wire [0:0] u_cla30_and14;
  wire [0:0] u_cla30_and15;
  wire [0:0] u_cla30_or7;
  wire [0:0] u_cla30_or8;
  wire [0:0] u_cla30_pg_logic6_or0;
  wire [0:0] u_cla30_pg_logic6_and0;
  wire [0:0] u_cla30_pg_logic6_xor0;
  wire [0:0] u_cla30_xor6;
  wire [0:0] u_cla30_and16;
  wire [0:0] u_cla30_and17;
  wire [0:0] u_cla30_and18;
  wire [0:0] u_cla30_and19;
  wire [0:0] u_cla30_and20;
  wire [0:0] u_cla30_and21;
  wire [0:0] u_cla30_or9;
  wire [0:0] u_cla30_or10;
  wire [0:0] u_cla30_or11;
  wire [0:0] u_cla30_pg_logic7_or0;
  wire [0:0] u_cla30_pg_logic7_and0;
  wire [0:0] u_cla30_pg_logic7_xor0;
  wire [0:0] u_cla30_xor7;
  wire [0:0] u_cla30_and22;
  wire [0:0] u_cla30_and23;
  wire [0:0] u_cla30_and24;
  wire [0:0] u_cla30_and25;
  wire [0:0] u_cla30_and26;
  wire [0:0] u_cla30_and27;
  wire [0:0] u_cla30_and28;
  wire [0:0] u_cla30_and29;
  wire [0:0] u_cla30_and30;
  wire [0:0] u_cla30_and31;
  wire [0:0] u_cla30_or12;
  wire [0:0] u_cla30_or13;
  wire [0:0] u_cla30_or14;
  wire [0:0] u_cla30_or15;
  wire [0:0] u_cla30_pg_logic8_or0;
  wire [0:0] u_cla30_pg_logic8_and0;
  wire [0:0] u_cla30_pg_logic8_xor0;
  wire [0:0] u_cla30_xor8;
  wire [0:0] u_cla30_and32;
  wire [0:0] u_cla30_or16;
  wire [0:0] u_cla30_pg_logic9_or0;
  wire [0:0] u_cla30_pg_logic9_and0;
  wire [0:0] u_cla30_pg_logic9_xor0;
  wire [0:0] u_cla30_xor9;
  wire [0:0] u_cla30_and33;
  wire [0:0] u_cla30_and34;
  wire [0:0] u_cla30_and35;
  wire [0:0] u_cla30_or17;
  wire [0:0] u_cla30_or18;
  wire [0:0] u_cla30_pg_logic10_or0;
  wire [0:0] u_cla30_pg_logic10_and0;
  wire [0:0] u_cla30_pg_logic10_xor0;
  wire [0:0] u_cla30_xor10;
  wire [0:0] u_cla30_and36;
  wire [0:0] u_cla30_and37;
  wire [0:0] u_cla30_and38;
  wire [0:0] u_cla30_and39;
  wire [0:0] u_cla30_and40;
  wire [0:0] u_cla30_and41;
  wire [0:0] u_cla30_or19;
  wire [0:0] u_cla30_or20;
  wire [0:0] u_cla30_or21;
  wire [0:0] u_cla30_pg_logic11_or0;
  wire [0:0] u_cla30_pg_logic11_and0;
  wire [0:0] u_cla30_pg_logic11_xor0;
  wire [0:0] u_cla30_xor11;
  wire [0:0] u_cla30_and42;
  wire [0:0] u_cla30_and43;
  wire [0:0] u_cla30_and44;
  wire [0:0] u_cla30_and45;
  wire [0:0] u_cla30_and46;
  wire [0:0] u_cla30_and47;
  wire [0:0] u_cla30_and48;
  wire [0:0] u_cla30_and49;
  wire [0:0] u_cla30_and50;
  wire [0:0] u_cla30_and51;
  wire [0:0] u_cla30_or22;
  wire [0:0] u_cla30_or23;
  wire [0:0] u_cla30_or24;
  wire [0:0] u_cla30_or25;
  wire [0:0] u_cla30_pg_logic12_or0;
  wire [0:0] u_cla30_pg_logic12_and0;
  wire [0:0] u_cla30_pg_logic12_xor0;
  wire [0:0] u_cla30_xor12;
  wire [0:0] u_cla30_and52;
  wire [0:0] u_cla30_or26;
  wire [0:0] u_cla30_pg_logic13_or0;
  wire [0:0] u_cla30_pg_logic13_and0;
  wire [0:0] u_cla30_pg_logic13_xor0;
  wire [0:0] u_cla30_xor13;
  wire [0:0] u_cla30_and53;
  wire [0:0] u_cla30_and54;
  wire [0:0] u_cla30_and55;
  wire [0:0] u_cla30_or27;
  wire [0:0] u_cla30_or28;
  wire [0:0] u_cla30_pg_logic14_or0;
  wire [0:0] u_cla30_pg_logic14_and0;
  wire [0:0] u_cla30_pg_logic14_xor0;
  wire [0:0] u_cla30_xor14;
  wire [0:0] u_cla30_and56;
  wire [0:0] u_cla30_and57;
  wire [0:0] u_cla30_and58;
  wire [0:0] u_cla30_and59;
  wire [0:0] u_cla30_and60;
  wire [0:0] u_cla30_and61;
  wire [0:0] u_cla30_or29;
  wire [0:0] u_cla30_or30;
  wire [0:0] u_cla30_or31;
  wire [0:0] u_cla30_pg_logic15_or0;
  wire [0:0] u_cla30_pg_logic15_and0;
  wire [0:0] u_cla30_pg_logic15_xor0;
  wire [0:0] u_cla30_xor15;
  wire [0:0] u_cla30_and62;
  wire [0:0] u_cla30_and63;
  wire [0:0] u_cla30_and64;
  wire [0:0] u_cla30_and65;
  wire [0:0] u_cla30_and66;
  wire [0:0] u_cla30_and67;
  wire [0:0] u_cla30_and68;
  wire [0:0] u_cla30_and69;
  wire [0:0] u_cla30_and70;
  wire [0:0] u_cla30_and71;
  wire [0:0] u_cla30_or32;
  wire [0:0] u_cla30_or33;
  wire [0:0] u_cla30_or34;
  wire [0:0] u_cla30_or35;
  wire [0:0] u_cla30_pg_logic16_or0;
  wire [0:0] u_cla30_pg_logic16_and0;
  wire [0:0] u_cla30_pg_logic16_xor0;
  wire [0:0] u_cla30_xor16;
  wire [0:0] u_cla30_and72;
  wire [0:0] u_cla30_or36;
  wire [0:0] u_cla30_pg_logic17_or0;
  wire [0:0] u_cla30_pg_logic17_and0;
  wire [0:0] u_cla30_pg_logic17_xor0;
  wire [0:0] u_cla30_xor17;
  wire [0:0] u_cla30_and73;
  wire [0:0] u_cla30_and74;
  wire [0:0] u_cla30_and75;
  wire [0:0] u_cla30_or37;
  wire [0:0] u_cla30_or38;
  wire [0:0] u_cla30_pg_logic18_or0;
  wire [0:0] u_cla30_pg_logic18_and0;
  wire [0:0] u_cla30_pg_logic18_xor0;
  wire [0:0] u_cla30_xor18;
  wire [0:0] u_cla30_and76;
  wire [0:0] u_cla30_and77;
  wire [0:0] u_cla30_and78;
  wire [0:0] u_cla30_and79;
  wire [0:0] u_cla30_and80;
  wire [0:0] u_cla30_and81;
  wire [0:0] u_cla30_or39;
  wire [0:0] u_cla30_or40;
  wire [0:0] u_cla30_or41;
  wire [0:0] u_cla30_pg_logic19_or0;
  wire [0:0] u_cla30_pg_logic19_and0;
  wire [0:0] u_cla30_pg_logic19_xor0;
  wire [0:0] u_cla30_xor19;
  wire [0:0] u_cla30_and82;
  wire [0:0] u_cla30_and83;
  wire [0:0] u_cla30_and84;
  wire [0:0] u_cla30_and85;
  wire [0:0] u_cla30_and86;
  wire [0:0] u_cla30_and87;
  wire [0:0] u_cla30_and88;
  wire [0:0] u_cla30_and89;
  wire [0:0] u_cla30_and90;
  wire [0:0] u_cla30_and91;
  wire [0:0] u_cla30_or42;
  wire [0:0] u_cla30_or43;
  wire [0:0] u_cla30_or44;
  wire [0:0] u_cla30_or45;
  wire [0:0] u_cla30_pg_logic20_or0;
  wire [0:0] u_cla30_pg_logic20_and0;
  wire [0:0] u_cla30_pg_logic20_xor0;
  wire [0:0] u_cla30_xor20;
  wire [0:0] u_cla30_and92;
  wire [0:0] u_cla30_or46;
  wire [0:0] u_cla30_pg_logic21_or0;
  wire [0:0] u_cla30_pg_logic21_and0;
  wire [0:0] u_cla30_pg_logic21_xor0;
  wire [0:0] u_cla30_xor21;
  wire [0:0] u_cla30_and93;
  wire [0:0] u_cla30_and94;
  wire [0:0] u_cla30_and95;
  wire [0:0] u_cla30_or47;
  wire [0:0] u_cla30_or48;
  wire [0:0] u_cla30_pg_logic22_or0;
  wire [0:0] u_cla30_pg_logic22_and0;
  wire [0:0] u_cla30_pg_logic22_xor0;
  wire [0:0] u_cla30_xor22;
  wire [0:0] u_cla30_and96;
  wire [0:0] u_cla30_and97;
  wire [0:0] u_cla30_and98;
  wire [0:0] u_cla30_and99;
  wire [0:0] u_cla30_and100;
  wire [0:0] u_cla30_and101;
  wire [0:0] u_cla30_or49;
  wire [0:0] u_cla30_or50;
  wire [0:0] u_cla30_or51;
  wire [0:0] u_cla30_pg_logic23_or0;
  wire [0:0] u_cla30_pg_logic23_and0;
  wire [0:0] u_cla30_pg_logic23_xor0;
  wire [0:0] u_cla30_xor23;
  wire [0:0] u_cla30_and102;
  wire [0:0] u_cla30_and103;
  wire [0:0] u_cla30_and104;
  wire [0:0] u_cla30_and105;
  wire [0:0] u_cla30_and106;
  wire [0:0] u_cla30_and107;
  wire [0:0] u_cla30_and108;
  wire [0:0] u_cla30_and109;
  wire [0:0] u_cla30_and110;
  wire [0:0] u_cla30_and111;
  wire [0:0] u_cla30_or52;
  wire [0:0] u_cla30_or53;
  wire [0:0] u_cla30_or54;
  wire [0:0] u_cla30_or55;
  wire [0:0] u_cla30_pg_logic24_or0;
  wire [0:0] u_cla30_pg_logic24_and0;
  wire [0:0] u_cla30_pg_logic24_xor0;
  wire [0:0] u_cla30_xor24;
  wire [0:0] u_cla30_and112;
  wire [0:0] u_cla30_or56;
  wire [0:0] u_cla30_pg_logic25_or0;
  wire [0:0] u_cla30_pg_logic25_and0;
  wire [0:0] u_cla30_pg_logic25_xor0;
  wire [0:0] u_cla30_xor25;
  wire [0:0] u_cla30_and113;
  wire [0:0] u_cla30_and114;
  wire [0:0] u_cla30_and115;
  wire [0:0] u_cla30_or57;
  wire [0:0] u_cla30_or58;
  wire [0:0] u_cla30_pg_logic26_or0;
  wire [0:0] u_cla30_pg_logic26_and0;
  wire [0:0] u_cla30_pg_logic26_xor0;
  wire [0:0] u_cla30_xor26;
  wire [0:0] u_cla30_and116;
  wire [0:0] u_cla30_and117;
  wire [0:0] u_cla30_and118;
  wire [0:0] u_cla30_and119;
  wire [0:0] u_cla30_and120;
  wire [0:0] u_cla30_and121;
  wire [0:0] u_cla30_or59;
  wire [0:0] u_cla30_or60;
  wire [0:0] u_cla30_or61;
  wire [0:0] u_cla30_pg_logic27_or0;
  wire [0:0] u_cla30_pg_logic27_and0;
  wire [0:0] u_cla30_pg_logic27_xor0;
  wire [0:0] u_cla30_xor27;
  wire [0:0] u_cla30_and122;
  wire [0:0] u_cla30_and123;
  wire [0:0] u_cla30_and124;
  wire [0:0] u_cla30_and125;
  wire [0:0] u_cla30_and126;
  wire [0:0] u_cla30_and127;
  wire [0:0] u_cla30_and128;
  wire [0:0] u_cla30_and129;
  wire [0:0] u_cla30_and130;
  wire [0:0] u_cla30_and131;
  wire [0:0] u_cla30_or62;
  wire [0:0] u_cla30_or63;
  wire [0:0] u_cla30_or64;
  wire [0:0] u_cla30_or65;
  wire [0:0] u_cla30_pg_logic28_or0;
  wire [0:0] u_cla30_pg_logic28_and0;
  wire [0:0] u_cla30_pg_logic28_xor0;
  wire [0:0] u_cla30_xor28;
  wire [0:0] u_cla30_and132;
  wire [0:0] u_cla30_or66;
  wire [0:0] u_cla30_pg_logic29_or0;
  wire [0:0] u_cla30_pg_logic29_and0;
  wire [0:0] u_cla30_pg_logic29_xor0;
  wire [0:0] u_cla30_xor29;
  wire [0:0] u_cla30_and133;
  wire [0:0] u_cla30_and134;
  wire [0:0] u_cla30_and135;
  wire [0:0] u_cla30_or67;
  wire [0:0] u_cla30_or68;

  pg_logic pg_logic_u_cla30_pg_logic0_out(.a(a[0]), .b(b[0]), .pg_logic_or0(u_cla30_pg_logic0_or0), .pg_logic_and0(u_cla30_pg_logic0_and0), .pg_logic_xor0(u_cla30_pg_logic0_xor0));
  pg_logic pg_logic_u_cla30_pg_logic1_out(.a(a[1]), .b(b[1]), .pg_logic_or0(u_cla30_pg_logic1_or0), .pg_logic_and0(u_cla30_pg_logic1_and0), .pg_logic_xor0(u_cla30_pg_logic1_xor0));
  xor_gate xor_gate_u_cla30_xor1(.a(u_cla30_pg_logic1_xor0[0]), .b(u_cla30_pg_logic0_and0[0]), .out(u_cla30_xor1));
  and_gate and_gate_u_cla30_and0(.a(u_cla30_pg_logic0_and0[0]), .b(u_cla30_pg_logic1_or0[0]), .out(u_cla30_and0));
  or_gate or_gate_u_cla30_or0(.a(u_cla30_pg_logic1_and0[0]), .b(u_cla30_and0[0]), .out(u_cla30_or0));
  pg_logic pg_logic_u_cla30_pg_logic2_out(.a(a[2]), .b(b[2]), .pg_logic_or0(u_cla30_pg_logic2_or0), .pg_logic_and0(u_cla30_pg_logic2_and0), .pg_logic_xor0(u_cla30_pg_logic2_xor0));
  xor_gate xor_gate_u_cla30_xor2(.a(u_cla30_pg_logic2_xor0[0]), .b(u_cla30_or0[0]), .out(u_cla30_xor2));
  and_gate and_gate_u_cla30_and1(.a(u_cla30_pg_logic2_or0[0]), .b(u_cla30_pg_logic0_or0[0]), .out(u_cla30_and1));
  and_gate and_gate_u_cla30_and2(.a(u_cla30_pg_logic0_and0[0]), .b(u_cla30_pg_logic2_or0[0]), .out(u_cla30_and2));
  and_gate and_gate_u_cla30_and3(.a(u_cla30_and2[0]), .b(u_cla30_pg_logic1_or0[0]), .out(u_cla30_and3));
  and_gate and_gate_u_cla30_and4(.a(u_cla30_pg_logic1_and0[0]), .b(u_cla30_pg_logic2_or0[0]), .out(u_cla30_and4));
  or_gate or_gate_u_cla30_or1(.a(u_cla30_and3[0]), .b(u_cla30_and4[0]), .out(u_cla30_or1));
  or_gate or_gate_u_cla30_or2(.a(u_cla30_pg_logic2_and0[0]), .b(u_cla30_or1[0]), .out(u_cla30_or2));
  pg_logic pg_logic_u_cla30_pg_logic3_out(.a(a[3]), .b(b[3]), .pg_logic_or0(u_cla30_pg_logic3_or0), .pg_logic_and0(u_cla30_pg_logic3_and0), .pg_logic_xor0(u_cla30_pg_logic3_xor0));
  xor_gate xor_gate_u_cla30_xor3(.a(u_cla30_pg_logic3_xor0[0]), .b(u_cla30_or2[0]), .out(u_cla30_xor3));
  and_gate and_gate_u_cla30_and5(.a(u_cla30_pg_logic3_or0[0]), .b(u_cla30_pg_logic1_or0[0]), .out(u_cla30_and5));
  and_gate and_gate_u_cla30_and6(.a(u_cla30_pg_logic0_and0[0]), .b(u_cla30_pg_logic2_or0[0]), .out(u_cla30_and6));
  and_gate and_gate_u_cla30_and7(.a(u_cla30_pg_logic3_or0[0]), .b(u_cla30_pg_logic1_or0[0]), .out(u_cla30_and7));
  and_gate and_gate_u_cla30_and8(.a(u_cla30_and6[0]), .b(u_cla30_and7[0]), .out(u_cla30_and8));
  and_gate and_gate_u_cla30_and9(.a(u_cla30_pg_logic1_and0[0]), .b(u_cla30_pg_logic3_or0[0]), .out(u_cla30_and9));
  and_gate and_gate_u_cla30_and10(.a(u_cla30_and9[0]), .b(u_cla30_pg_logic2_or0[0]), .out(u_cla30_and10));
  and_gate and_gate_u_cla30_and11(.a(u_cla30_pg_logic2_and0[0]), .b(u_cla30_pg_logic3_or0[0]), .out(u_cla30_and11));
  or_gate or_gate_u_cla30_or3(.a(u_cla30_and8[0]), .b(u_cla30_and11[0]), .out(u_cla30_or3));
  or_gate or_gate_u_cla30_or4(.a(u_cla30_and10[0]), .b(u_cla30_or3[0]), .out(u_cla30_or4));
  or_gate or_gate_u_cla30_or5(.a(u_cla30_pg_logic3_and0[0]), .b(u_cla30_or4[0]), .out(u_cla30_or5));
  pg_logic pg_logic_u_cla30_pg_logic4_out(.a(a[4]), .b(b[4]), .pg_logic_or0(u_cla30_pg_logic4_or0), .pg_logic_and0(u_cla30_pg_logic4_and0), .pg_logic_xor0(u_cla30_pg_logic4_xor0));
  xor_gate xor_gate_u_cla30_xor4(.a(u_cla30_pg_logic4_xor0[0]), .b(u_cla30_or5[0]), .out(u_cla30_xor4));
  and_gate and_gate_u_cla30_and12(.a(u_cla30_or5[0]), .b(u_cla30_pg_logic4_or0[0]), .out(u_cla30_and12));
  or_gate or_gate_u_cla30_or6(.a(u_cla30_pg_logic4_and0[0]), .b(u_cla30_and12[0]), .out(u_cla30_or6));
  pg_logic pg_logic_u_cla30_pg_logic5_out(.a(a[5]), .b(b[5]), .pg_logic_or0(u_cla30_pg_logic5_or0), .pg_logic_and0(u_cla30_pg_logic5_and0), .pg_logic_xor0(u_cla30_pg_logic5_xor0));
  xor_gate xor_gate_u_cla30_xor5(.a(u_cla30_pg_logic5_xor0[0]), .b(u_cla30_or6[0]), .out(u_cla30_xor5));
  and_gate and_gate_u_cla30_and13(.a(u_cla30_or5[0]), .b(u_cla30_pg_logic5_or0[0]), .out(u_cla30_and13));
  and_gate and_gate_u_cla30_and14(.a(u_cla30_and13[0]), .b(u_cla30_pg_logic4_or0[0]), .out(u_cla30_and14));
  and_gate and_gate_u_cla30_and15(.a(u_cla30_pg_logic4_and0[0]), .b(u_cla30_pg_logic5_or0[0]), .out(u_cla30_and15));
  or_gate or_gate_u_cla30_or7(.a(u_cla30_and14[0]), .b(u_cla30_and15[0]), .out(u_cla30_or7));
  or_gate or_gate_u_cla30_or8(.a(u_cla30_pg_logic5_and0[0]), .b(u_cla30_or7[0]), .out(u_cla30_or8));
  pg_logic pg_logic_u_cla30_pg_logic6_out(.a(a[6]), .b(b[6]), .pg_logic_or0(u_cla30_pg_logic6_or0), .pg_logic_and0(u_cla30_pg_logic6_and0), .pg_logic_xor0(u_cla30_pg_logic6_xor0));
  xor_gate xor_gate_u_cla30_xor6(.a(u_cla30_pg_logic6_xor0[0]), .b(u_cla30_or8[0]), .out(u_cla30_xor6));
  and_gate and_gate_u_cla30_and16(.a(u_cla30_or5[0]), .b(u_cla30_pg_logic5_or0[0]), .out(u_cla30_and16));
  and_gate and_gate_u_cla30_and17(.a(u_cla30_pg_logic6_or0[0]), .b(u_cla30_pg_logic4_or0[0]), .out(u_cla30_and17));
  and_gate and_gate_u_cla30_and18(.a(u_cla30_and16[0]), .b(u_cla30_and17[0]), .out(u_cla30_and18));
  and_gate and_gate_u_cla30_and19(.a(u_cla30_pg_logic4_and0[0]), .b(u_cla30_pg_logic6_or0[0]), .out(u_cla30_and19));
  and_gate and_gate_u_cla30_and20(.a(u_cla30_and19[0]), .b(u_cla30_pg_logic5_or0[0]), .out(u_cla30_and20));
  and_gate and_gate_u_cla30_and21(.a(u_cla30_pg_logic5_and0[0]), .b(u_cla30_pg_logic6_or0[0]), .out(u_cla30_and21));
  or_gate or_gate_u_cla30_or9(.a(u_cla30_and18[0]), .b(u_cla30_and20[0]), .out(u_cla30_or9));
  or_gate or_gate_u_cla30_or10(.a(u_cla30_or9[0]), .b(u_cla30_and21[0]), .out(u_cla30_or10));
  or_gate or_gate_u_cla30_or11(.a(u_cla30_pg_logic6_and0[0]), .b(u_cla30_or10[0]), .out(u_cla30_or11));
  pg_logic pg_logic_u_cla30_pg_logic7_out(.a(a[7]), .b(b[7]), .pg_logic_or0(u_cla30_pg_logic7_or0), .pg_logic_and0(u_cla30_pg_logic7_and0), .pg_logic_xor0(u_cla30_pg_logic7_xor0));
  xor_gate xor_gate_u_cla30_xor7(.a(u_cla30_pg_logic7_xor0[0]), .b(u_cla30_or11[0]), .out(u_cla30_xor7));
  and_gate and_gate_u_cla30_and22(.a(u_cla30_or5[0]), .b(u_cla30_pg_logic6_or0[0]), .out(u_cla30_and22));
  and_gate and_gate_u_cla30_and23(.a(u_cla30_pg_logic7_or0[0]), .b(u_cla30_pg_logic5_or0[0]), .out(u_cla30_and23));
  and_gate and_gate_u_cla30_and24(.a(u_cla30_and22[0]), .b(u_cla30_and23[0]), .out(u_cla30_and24));
  and_gate and_gate_u_cla30_and25(.a(u_cla30_and24[0]), .b(u_cla30_pg_logic4_or0[0]), .out(u_cla30_and25));
  and_gate and_gate_u_cla30_and26(.a(u_cla30_pg_logic4_and0[0]), .b(u_cla30_pg_logic6_or0[0]), .out(u_cla30_and26));
  and_gate and_gate_u_cla30_and27(.a(u_cla30_pg_logic7_or0[0]), .b(u_cla30_pg_logic5_or0[0]), .out(u_cla30_and27));
  and_gate and_gate_u_cla30_and28(.a(u_cla30_and26[0]), .b(u_cla30_and27[0]), .out(u_cla30_and28));
  and_gate and_gate_u_cla30_and29(.a(u_cla30_pg_logic5_and0[0]), .b(u_cla30_pg_logic7_or0[0]), .out(u_cla30_and29));
  and_gate and_gate_u_cla30_and30(.a(u_cla30_and29[0]), .b(u_cla30_pg_logic6_or0[0]), .out(u_cla30_and30));
  and_gate and_gate_u_cla30_and31(.a(u_cla30_pg_logic6_and0[0]), .b(u_cla30_pg_logic7_or0[0]), .out(u_cla30_and31));
  or_gate or_gate_u_cla30_or12(.a(u_cla30_and25[0]), .b(u_cla30_and30[0]), .out(u_cla30_or12));
  or_gate or_gate_u_cla30_or13(.a(u_cla30_and28[0]), .b(u_cla30_and31[0]), .out(u_cla30_or13));
  or_gate or_gate_u_cla30_or14(.a(u_cla30_or12[0]), .b(u_cla30_or13[0]), .out(u_cla30_or14));
  or_gate or_gate_u_cla30_or15(.a(u_cla30_pg_logic7_and0[0]), .b(u_cla30_or14[0]), .out(u_cla30_or15));
  pg_logic pg_logic_u_cla30_pg_logic8_out(.a(a[8]), .b(b[8]), .pg_logic_or0(u_cla30_pg_logic8_or0), .pg_logic_and0(u_cla30_pg_logic8_and0), .pg_logic_xor0(u_cla30_pg_logic8_xor0));
  xor_gate xor_gate_u_cla30_xor8(.a(u_cla30_pg_logic8_xor0[0]), .b(u_cla30_or15[0]), .out(u_cla30_xor8));
  and_gate and_gate_u_cla30_and32(.a(u_cla30_or15[0]), .b(u_cla30_pg_logic8_or0[0]), .out(u_cla30_and32));
  or_gate or_gate_u_cla30_or16(.a(u_cla30_pg_logic8_and0[0]), .b(u_cla30_and32[0]), .out(u_cla30_or16));
  pg_logic pg_logic_u_cla30_pg_logic9_out(.a(a[9]), .b(b[9]), .pg_logic_or0(u_cla30_pg_logic9_or0), .pg_logic_and0(u_cla30_pg_logic9_and0), .pg_logic_xor0(u_cla30_pg_logic9_xor0));
  xor_gate xor_gate_u_cla30_xor9(.a(u_cla30_pg_logic9_xor0[0]), .b(u_cla30_or16[0]), .out(u_cla30_xor9));
  and_gate and_gate_u_cla30_and33(.a(u_cla30_or15[0]), .b(u_cla30_pg_logic9_or0[0]), .out(u_cla30_and33));
  and_gate and_gate_u_cla30_and34(.a(u_cla30_and33[0]), .b(u_cla30_pg_logic8_or0[0]), .out(u_cla30_and34));
  and_gate and_gate_u_cla30_and35(.a(u_cla30_pg_logic8_and0[0]), .b(u_cla30_pg_logic9_or0[0]), .out(u_cla30_and35));
  or_gate or_gate_u_cla30_or17(.a(u_cla30_and34[0]), .b(u_cla30_and35[0]), .out(u_cla30_or17));
  or_gate or_gate_u_cla30_or18(.a(u_cla30_pg_logic9_and0[0]), .b(u_cla30_or17[0]), .out(u_cla30_or18));
  pg_logic pg_logic_u_cla30_pg_logic10_out(.a(a[10]), .b(b[10]), .pg_logic_or0(u_cla30_pg_logic10_or0), .pg_logic_and0(u_cla30_pg_logic10_and0), .pg_logic_xor0(u_cla30_pg_logic10_xor0));
  xor_gate xor_gate_u_cla30_xor10(.a(u_cla30_pg_logic10_xor0[0]), .b(u_cla30_or18[0]), .out(u_cla30_xor10));
  and_gate and_gate_u_cla30_and36(.a(u_cla30_or15[0]), .b(u_cla30_pg_logic9_or0[0]), .out(u_cla30_and36));
  and_gate and_gate_u_cla30_and37(.a(u_cla30_pg_logic10_or0[0]), .b(u_cla30_pg_logic8_or0[0]), .out(u_cla30_and37));
  and_gate and_gate_u_cla30_and38(.a(u_cla30_and36[0]), .b(u_cla30_and37[0]), .out(u_cla30_and38));
  and_gate and_gate_u_cla30_and39(.a(u_cla30_pg_logic8_and0[0]), .b(u_cla30_pg_logic10_or0[0]), .out(u_cla30_and39));
  and_gate and_gate_u_cla30_and40(.a(u_cla30_and39[0]), .b(u_cla30_pg_logic9_or0[0]), .out(u_cla30_and40));
  and_gate and_gate_u_cla30_and41(.a(u_cla30_pg_logic9_and0[0]), .b(u_cla30_pg_logic10_or0[0]), .out(u_cla30_and41));
  or_gate or_gate_u_cla30_or19(.a(u_cla30_and38[0]), .b(u_cla30_and40[0]), .out(u_cla30_or19));
  or_gate or_gate_u_cla30_or20(.a(u_cla30_or19[0]), .b(u_cla30_and41[0]), .out(u_cla30_or20));
  or_gate or_gate_u_cla30_or21(.a(u_cla30_pg_logic10_and0[0]), .b(u_cla30_or20[0]), .out(u_cla30_or21));
  pg_logic pg_logic_u_cla30_pg_logic11_out(.a(a[11]), .b(b[11]), .pg_logic_or0(u_cla30_pg_logic11_or0), .pg_logic_and0(u_cla30_pg_logic11_and0), .pg_logic_xor0(u_cla30_pg_logic11_xor0));
  xor_gate xor_gate_u_cla30_xor11(.a(u_cla30_pg_logic11_xor0[0]), .b(u_cla30_or21[0]), .out(u_cla30_xor11));
  and_gate and_gate_u_cla30_and42(.a(u_cla30_or15[0]), .b(u_cla30_pg_logic10_or0[0]), .out(u_cla30_and42));
  and_gate and_gate_u_cla30_and43(.a(u_cla30_pg_logic11_or0[0]), .b(u_cla30_pg_logic9_or0[0]), .out(u_cla30_and43));
  and_gate and_gate_u_cla30_and44(.a(u_cla30_and42[0]), .b(u_cla30_and43[0]), .out(u_cla30_and44));
  and_gate and_gate_u_cla30_and45(.a(u_cla30_and44[0]), .b(u_cla30_pg_logic8_or0[0]), .out(u_cla30_and45));
  and_gate and_gate_u_cla30_and46(.a(u_cla30_pg_logic8_and0[0]), .b(u_cla30_pg_logic10_or0[0]), .out(u_cla30_and46));
  and_gate and_gate_u_cla30_and47(.a(u_cla30_pg_logic11_or0[0]), .b(u_cla30_pg_logic9_or0[0]), .out(u_cla30_and47));
  and_gate and_gate_u_cla30_and48(.a(u_cla30_and46[0]), .b(u_cla30_and47[0]), .out(u_cla30_and48));
  and_gate and_gate_u_cla30_and49(.a(u_cla30_pg_logic9_and0[0]), .b(u_cla30_pg_logic11_or0[0]), .out(u_cla30_and49));
  and_gate and_gate_u_cla30_and50(.a(u_cla30_and49[0]), .b(u_cla30_pg_logic10_or0[0]), .out(u_cla30_and50));
  and_gate and_gate_u_cla30_and51(.a(u_cla30_pg_logic10_and0[0]), .b(u_cla30_pg_logic11_or0[0]), .out(u_cla30_and51));
  or_gate or_gate_u_cla30_or22(.a(u_cla30_and45[0]), .b(u_cla30_and50[0]), .out(u_cla30_or22));
  or_gate or_gate_u_cla30_or23(.a(u_cla30_and48[0]), .b(u_cla30_and51[0]), .out(u_cla30_or23));
  or_gate or_gate_u_cla30_or24(.a(u_cla30_or22[0]), .b(u_cla30_or23[0]), .out(u_cla30_or24));
  or_gate or_gate_u_cla30_or25(.a(u_cla30_pg_logic11_and0[0]), .b(u_cla30_or24[0]), .out(u_cla30_or25));
  pg_logic pg_logic_u_cla30_pg_logic12_out(.a(a[12]), .b(b[12]), .pg_logic_or0(u_cla30_pg_logic12_or0), .pg_logic_and0(u_cla30_pg_logic12_and0), .pg_logic_xor0(u_cla30_pg_logic12_xor0));
  xor_gate xor_gate_u_cla30_xor12(.a(u_cla30_pg_logic12_xor0[0]), .b(u_cla30_or25[0]), .out(u_cla30_xor12));
  and_gate and_gate_u_cla30_and52(.a(u_cla30_or25[0]), .b(u_cla30_pg_logic12_or0[0]), .out(u_cla30_and52));
  or_gate or_gate_u_cla30_or26(.a(u_cla30_pg_logic12_and0[0]), .b(u_cla30_and52[0]), .out(u_cla30_or26));
  pg_logic pg_logic_u_cla30_pg_logic13_out(.a(a[13]), .b(b[13]), .pg_logic_or0(u_cla30_pg_logic13_or0), .pg_logic_and0(u_cla30_pg_logic13_and0), .pg_logic_xor0(u_cla30_pg_logic13_xor0));
  xor_gate xor_gate_u_cla30_xor13(.a(u_cla30_pg_logic13_xor0[0]), .b(u_cla30_or26[0]), .out(u_cla30_xor13));
  and_gate and_gate_u_cla30_and53(.a(u_cla30_or25[0]), .b(u_cla30_pg_logic13_or0[0]), .out(u_cla30_and53));
  and_gate and_gate_u_cla30_and54(.a(u_cla30_and53[0]), .b(u_cla30_pg_logic12_or0[0]), .out(u_cla30_and54));
  and_gate and_gate_u_cla30_and55(.a(u_cla30_pg_logic12_and0[0]), .b(u_cla30_pg_logic13_or0[0]), .out(u_cla30_and55));
  or_gate or_gate_u_cla30_or27(.a(u_cla30_and54[0]), .b(u_cla30_and55[0]), .out(u_cla30_or27));
  or_gate or_gate_u_cla30_or28(.a(u_cla30_pg_logic13_and0[0]), .b(u_cla30_or27[0]), .out(u_cla30_or28));
  pg_logic pg_logic_u_cla30_pg_logic14_out(.a(a[14]), .b(b[14]), .pg_logic_or0(u_cla30_pg_logic14_or0), .pg_logic_and0(u_cla30_pg_logic14_and0), .pg_logic_xor0(u_cla30_pg_logic14_xor0));
  xor_gate xor_gate_u_cla30_xor14(.a(u_cla30_pg_logic14_xor0[0]), .b(u_cla30_or28[0]), .out(u_cla30_xor14));
  and_gate and_gate_u_cla30_and56(.a(u_cla30_or25[0]), .b(u_cla30_pg_logic13_or0[0]), .out(u_cla30_and56));
  and_gate and_gate_u_cla30_and57(.a(u_cla30_pg_logic14_or0[0]), .b(u_cla30_pg_logic12_or0[0]), .out(u_cla30_and57));
  and_gate and_gate_u_cla30_and58(.a(u_cla30_and56[0]), .b(u_cla30_and57[0]), .out(u_cla30_and58));
  and_gate and_gate_u_cla30_and59(.a(u_cla30_pg_logic12_and0[0]), .b(u_cla30_pg_logic14_or0[0]), .out(u_cla30_and59));
  and_gate and_gate_u_cla30_and60(.a(u_cla30_and59[0]), .b(u_cla30_pg_logic13_or0[0]), .out(u_cla30_and60));
  and_gate and_gate_u_cla30_and61(.a(u_cla30_pg_logic13_and0[0]), .b(u_cla30_pg_logic14_or0[0]), .out(u_cla30_and61));
  or_gate or_gate_u_cla30_or29(.a(u_cla30_and58[0]), .b(u_cla30_and60[0]), .out(u_cla30_or29));
  or_gate or_gate_u_cla30_or30(.a(u_cla30_or29[0]), .b(u_cla30_and61[0]), .out(u_cla30_or30));
  or_gate or_gate_u_cla30_or31(.a(u_cla30_pg_logic14_and0[0]), .b(u_cla30_or30[0]), .out(u_cla30_or31));
  pg_logic pg_logic_u_cla30_pg_logic15_out(.a(a[15]), .b(b[15]), .pg_logic_or0(u_cla30_pg_logic15_or0), .pg_logic_and0(u_cla30_pg_logic15_and0), .pg_logic_xor0(u_cla30_pg_logic15_xor0));
  xor_gate xor_gate_u_cla30_xor15(.a(u_cla30_pg_logic15_xor0[0]), .b(u_cla30_or31[0]), .out(u_cla30_xor15));
  and_gate and_gate_u_cla30_and62(.a(u_cla30_or25[0]), .b(u_cla30_pg_logic14_or0[0]), .out(u_cla30_and62));
  and_gate and_gate_u_cla30_and63(.a(u_cla30_pg_logic15_or0[0]), .b(u_cla30_pg_logic13_or0[0]), .out(u_cla30_and63));
  and_gate and_gate_u_cla30_and64(.a(u_cla30_and62[0]), .b(u_cla30_and63[0]), .out(u_cla30_and64));
  and_gate and_gate_u_cla30_and65(.a(u_cla30_and64[0]), .b(u_cla30_pg_logic12_or0[0]), .out(u_cla30_and65));
  and_gate and_gate_u_cla30_and66(.a(u_cla30_pg_logic12_and0[0]), .b(u_cla30_pg_logic14_or0[0]), .out(u_cla30_and66));
  and_gate and_gate_u_cla30_and67(.a(u_cla30_pg_logic15_or0[0]), .b(u_cla30_pg_logic13_or0[0]), .out(u_cla30_and67));
  and_gate and_gate_u_cla30_and68(.a(u_cla30_and66[0]), .b(u_cla30_and67[0]), .out(u_cla30_and68));
  and_gate and_gate_u_cla30_and69(.a(u_cla30_pg_logic13_and0[0]), .b(u_cla30_pg_logic15_or0[0]), .out(u_cla30_and69));
  and_gate and_gate_u_cla30_and70(.a(u_cla30_and69[0]), .b(u_cla30_pg_logic14_or0[0]), .out(u_cla30_and70));
  and_gate and_gate_u_cla30_and71(.a(u_cla30_pg_logic14_and0[0]), .b(u_cla30_pg_logic15_or0[0]), .out(u_cla30_and71));
  or_gate or_gate_u_cla30_or32(.a(u_cla30_and65[0]), .b(u_cla30_and70[0]), .out(u_cla30_or32));
  or_gate or_gate_u_cla30_or33(.a(u_cla30_and68[0]), .b(u_cla30_and71[0]), .out(u_cla30_or33));
  or_gate or_gate_u_cla30_or34(.a(u_cla30_or32[0]), .b(u_cla30_or33[0]), .out(u_cla30_or34));
  or_gate or_gate_u_cla30_or35(.a(u_cla30_pg_logic15_and0[0]), .b(u_cla30_or34[0]), .out(u_cla30_or35));
  pg_logic pg_logic_u_cla30_pg_logic16_out(.a(a[16]), .b(b[16]), .pg_logic_or0(u_cla30_pg_logic16_or0), .pg_logic_and0(u_cla30_pg_logic16_and0), .pg_logic_xor0(u_cla30_pg_logic16_xor0));
  xor_gate xor_gate_u_cla30_xor16(.a(u_cla30_pg_logic16_xor0[0]), .b(u_cla30_or35[0]), .out(u_cla30_xor16));
  and_gate and_gate_u_cla30_and72(.a(u_cla30_or35[0]), .b(u_cla30_pg_logic16_or0[0]), .out(u_cla30_and72));
  or_gate or_gate_u_cla30_or36(.a(u_cla30_pg_logic16_and0[0]), .b(u_cla30_and72[0]), .out(u_cla30_or36));
  pg_logic pg_logic_u_cla30_pg_logic17_out(.a(a[17]), .b(b[17]), .pg_logic_or0(u_cla30_pg_logic17_or0), .pg_logic_and0(u_cla30_pg_logic17_and0), .pg_logic_xor0(u_cla30_pg_logic17_xor0));
  xor_gate xor_gate_u_cla30_xor17(.a(u_cla30_pg_logic17_xor0[0]), .b(u_cla30_or36[0]), .out(u_cla30_xor17));
  and_gate and_gate_u_cla30_and73(.a(u_cla30_or35[0]), .b(u_cla30_pg_logic17_or0[0]), .out(u_cla30_and73));
  and_gate and_gate_u_cla30_and74(.a(u_cla30_and73[0]), .b(u_cla30_pg_logic16_or0[0]), .out(u_cla30_and74));
  and_gate and_gate_u_cla30_and75(.a(u_cla30_pg_logic16_and0[0]), .b(u_cla30_pg_logic17_or0[0]), .out(u_cla30_and75));
  or_gate or_gate_u_cla30_or37(.a(u_cla30_and74[0]), .b(u_cla30_and75[0]), .out(u_cla30_or37));
  or_gate or_gate_u_cla30_or38(.a(u_cla30_pg_logic17_and0[0]), .b(u_cla30_or37[0]), .out(u_cla30_or38));
  pg_logic pg_logic_u_cla30_pg_logic18_out(.a(a[18]), .b(b[18]), .pg_logic_or0(u_cla30_pg_logic18_or0), .pg_logic_and0(u_cla30_pg_logic18_and0), .pg_logic_xor0(u_cla30_pg_logic18_xor0));
  xor_gate xor_gate_u_cla30_xor18(.a(u_cla30_pg_logic18_xor0[0]), .b(u_cla30_or38[0]), .out(u_cla30_xor18));
  and_gate and_gate_u_cla30_and76(.a(u_cla30_or35[0]), .b(u_cla30_pg_logic17_or0[0]), .out(u_cla30_and76));
  and_gate and_gate_u_cla30_and77(.a(u_cla30_pg_logic18_or0[0]), .b(u_cla30_pg_logic16_or0[0]), .out(u_cla30_and77));
  and_gate and_gate_u_cla30_and78(.a(u_cla30_and76[0]), .b(u_cla30_and77[0]), .out(u_cla30_and78));
  and_gate and_gate_u_cla30_and79(.a(u_cla30_pg_logic16_and0[0]), .b(u_cla30_pg_logic18_or0[0]), .out(u_cla30_and79));
  and_gate and_gate_u_cla30_and80(.a(u_cla30_and79[0]), .b(u_cla30_pg_logic17_or0[0]), .out(u_cla30_and80));
  and_gate and_gate_u_cla30_and81(.a(u_cla30_pg_logic17_and0[0]), .b(u_cla30_pg_logic18_or0[0]), .out(u_cla30_and81));
  or_gate or_gate_u_cla30_or39(.a(u_cla30_and78[0]), .b(u_cla30_and80[0]), .out(u_cla30_or39));
  or_gate or_gate_u_cla30_or40(.a(u_cla30_or39[0]), .b(u_cla30_and81[0]), .out(u_cla30_or40));
  or_gate or_gate_u_cla30_or41(.a(u_cla30_pg_logic18_and0[0]), .b(u_cla30_or40[0]), .out(u_cla30_or41));
  pg_logic pg_logic_u_cla30_pg_logic19_out(.a(a[19]), .b(b[19]), .pg_logic_or0(u_cla30_pg_logic19_or0), .pg_logic_and0(u_cla30_pg_logic19_and0), .pg_logic_xor0(u_cla30_pg_logic19_xor0));
  xor_gate xor_gate_u_cla30_xor19(.a(u_cla30_pg_logic19_xor0[0]), .b(u_cla30_or41[0]), .out(u_cla30_xor19));
  and_gate and_gate_u_cla30_and82(.a(u_cla30_or35[0]), .b(u_cla30_pg_logic18_or0[0]), .out(u_cla30_and82));
  and_gate and_gate_u_cla30_and83(.a(u_cla30_pg_logic19_or0[0]), .b(u_cla30_pg_logic17_or0[0]), .out(u_cla30_and83));
  and_gate and_gate_u_cla30_and84(.a(u_cla30_and82[0]), .b(u_cla30_and83[0]), .out(u_cla30_and84));
  and_gate and_gate_u_cla30_and85(.a(u_cla30_and84[0]), .b(u_cla30_pg_logic16_or0[0]), .out(u_cla30_and85));
  and_gate and_gate_u_cla30_and86(.a(u_cla30_pg_logic16_and0[0]), .b(u_cla30_pg_logic18_or0[0]), .out(u_cla30_and86));
  and_gate and_gate_u_cla30_and87(.a(u_cla30_pg_logic19_or0[0]), .b(u_cla30_pg_logic17_or0[0]), .out(u_cla30_and87));
  and_gate and_gate_u_cla30_and88(.a(u_cla30_and86[0]), .b(u_cla30_and87[0]), .out(u_cla30_and88));
  and_gate and_gate_u_cla30_and89(.a(u_cla30_pg_logic17_and0[0]), .b(u_cla30_pg_logic19_or0[0]), .out(u_cla30_and89));
  and_gate and_gate_u_cla30_and90(.a(u_cla30_and89[0]), .b(u_cla30_pg_logic18_or0[0]), .out(u_cla30_and90));
  and_gate and_gate_u_cla30_and91(.a(u_cla30_pg_logic18_and0[0]), .b(u_cla30_pg_logic19_or0[0]), .out(u_cla30_and91));
  or_gate or_gate_u_cla30_or42(.a(u_cla30_and85[0]), .b(u_cla30_and90[0]), .out(u_cla30_or42));
  or_gate or_gate_u_cla30_or43(.a(u_cla30_and88[0]), .b(u_cla30_and91[0]), .out(u_cla30_or43));
  or_gate or_gate_u_cla30_or44(.a(u_cla30_or42[0]), .b(u_cla30_or43[0]), .out(u_cla30_or44));
  or_gate or_gate_u_cla30_or45(.a(u_cla30_pg_logic19_and0[0]), .b(u_cla30_or44[0]), .out(u_cla30_or45));
  pg_logic pg_logic_u_cla30_pg_logic20_out(.a(a[20]), .b(b[20]), .pg_logic_or0(u_cla30_pg_logic20_or0), .pg_logic_and0(u_cla30_pg_logic20_and0), .pg_logic_xor0(u_cla30_pg_logic20_xor0));
  xor_gate xor_gate_u_cla30_xor20(.a(u_cla30_pg_logic20_xor0[0]), .b(u_cla30_or45[0]), .out(u_cla30_xor20));
  and_gate and_gate_u_cla30_and92(.a(u_cla30_or45[0]), .b(u_cla30_pg_logic20_or0[0]), .out(u_cla30_and92));
  or_gate or_gate_u_cla30_or46(.a(u_cla30_pg_logic20_and0[0]), .b(u_cla30_and92[0]), .out(u_cla30_or46));
  pg_logic pg_logic_u_cla30_pg_logic21_out(.a(a[21]), .b(b[21]), .pg_logic_or0(u_cla30_pg_logic21_or0), .pg_logic_and0(u_cla30_pg_logic21_and0), .pg_logic_xor0(u_cla30_pg_logic21_xor0));
  xor_gate xor_gate_u_cla30_xor21(.a(u_cla30_pg_logic21_xor0[0]), .b(u_cla30_or46[0]), .out(u_cla30_xor21));
  and_gate and_gate_u_cla30_and93(.a(u_cla30_or45[0]), .b(u_cla30_pg_logic21_or0[0]), .out(u_cla30_and93));
  and_gate and_gate_u_cla30_and94(.a(u_cla30_and93[0]), .b(u_cla30_pg_logic20_or0[0]), .out(u_cla30_and94));
  and_gate and_gate_u_cla30_and95(.a(u_cla30_pg_logic20_and0[0]), .b(u_cla30_pg_logic21_or0[0]), .out(u_cla30_and95));
  or_gate or_gate_u_cla30_or47(.a(u_cla30_and94[0]), .b(u_cla30_and95[0]), .out(u_cla30_or47));
  or_gate or_gate_u_cla30_or48(.a(u_cla30_pg_logic21_and0[0]), .b(u_cla30_or47[0]), .out(u_cla30_or48));
  pg_logic pg_logic_u_cla30_pg_logic22_out(.a(a[22]), .b(b[22]), .pg_logic_or0(u_cla30_pg_logic22_or0), .pg_logic_and0(u_cla30_pg_logic22_and0), .pg_logic_xor0(u_cla30_pg_logic22_xor0));
  xor_gate xor_gate_u_cla30_xor22(.a(u_cla30_pg_logic22_xor0[0]), .b(u_cla30_or48[0]), .out(u_cla30_xor22));
  and_gate and_gate_u_cla30_and96(.a(u_cla30_or45[0]), .b(u_cla30_pg_logic21_or0[0]), .out(u_cla30_and96));
  and_gate and_gate_u_cla30_and97(.a(u_cla30_pg_logic22_or0[0]), .b(u_cla30_pg_logic20_or0[0]), .out(u_cla30_and97));
  and_gate and_gate_u_cla30_and98(.a(u_cla30_and96[0]), .b(u_cla30_and97[0]), .out(u_cla30_and98));
  and_gate and_gate_u_cla30_and99(.a(u_cla30_pg_logic20_and0[0]), .b(u_cla30_pg_logic22_or0[0]), .out(u_cla30_and99));
  and_gate and_gate_u_cla30_and100(.a(u_cla30_and99[0]), .b(u_cla30_pg_logic21_or0[0]), .out(u_cla30_and100));
  and_gate and_gate_u_cla30_and101(.a(u_cla30_pg_logic21_and0[0]), .b(u_cla30_pg_logic22_or0[0]), .out(u_cla30_and101));
  or_gate or_gate_u_cla30_or49(.a(u_cla30_and98[0]), .b(u_cla30_and100[0]), .out(u_cla30_or49));
  or_gate or_gate_u_cla30_or50(.a(u_cla30_or49[0]), .b(u_cla30_and101[0]), .out(u_cla30_or50));
  or_gate or_gate_u_cla30_or51(.a(u_cla30_pg_logic22_and0[0]), .b(u_cla30_or50[0]), .out(u_cla30_or51));
  pg_logic pg_logic_u_cla30_pg_logic23_out(.a(a[23]), .b(b[23]), .pg_logic_or0(u_cla30_pg_logic23_or0), .pg_logic_and0(u_cla30_pg_logic23_and0), .pg_logic_xor0(u_cla30_pg_logic23_xor0));
  xor_gate xor_gate_u_cla30_xor23(.a(u_cla30_pg_logic23_xor0[0]), .b(u_cla30_or51[0]), .out(u_cla30_xor23));
  and_gate and_gate_u_cla30_and102(.a(u_cla30_or45[0]), .b(u_cla30_pg_logic22_or0[0]), .out(u_cla30_and102));
  and_gate and_gate_u_cla30_and103(.a(u_cla30_pg_logic23_or0[0]), .b(u_cla30_pg_logic21_or0[0]), .out(u_cla30_and103));
  and_gate and_gate_u_cla30_and104(.a(u_cla30_and102[0]), .b(u_cla30_and103[0]), .out(u_cla30_and104));
  and_gate and_gate_u_cla30_and105(.a(u_cla30_and104[0]), .b(u_cla30_pg_logic20_or0[0]), .out(u_cla30_and105));
  and_gate and_gate_u_cla30_and106(.a(u_cla30_pg_logic20_and0[0]), .b(u_cla30_pg_logic22_or0[0]), .out(u_cla30_and106));
  and_gate and_gate_u_cla30_and107(.a(u_cla30_pg_logic23_or0[0]), .b(u_cla30_pg_logic21_or0[0]), .out(u_cla30_and107));
  and_gate and_gate_u_cla30_and108(.a(u_cla30_and106[0]), .b(u_cla30_and107[0]), .out(u_cla30_and108));
  and_gate and_gate_u_cla30_and109(.a(u_cla30_pg_logic21_and0[0]), .b(u_cla30_pg_logic23_or0[0]), .out(u_cla30_and109));
  and_gate and_gate_u_cla30_and110(.a(u_cla30_and109[0]), .b(u_cla30_pg_logic22_or0[0]), .out(u_cla30_and110));
  and_gate and_gate_u_cla30_and111(.a(u_cla30_pg_logic22_and0[0]), .b(u_cla30_pg_logic23_or0[0]), .out(u_cla30_and111));
  or_gate or_gate_u_cla30_or52(.a(u_cla30_and105[0]), .b(u_cla30_and110[0]), .out(u_cla30_or52));
  or_gate or_gate_u_cla30_or53(.a(u_cla30_and108[0]), .b(u_cla30_and111[0]), .out(u_cla30_or53));
  or_gate or_gate_u_cla30_or54(.a(u_cla30_or52[0]), .b(u_cla30_or53[0]), .out(u_cla30_or54));
  or_gate or_gate_u_cla30_or55(.a(u_cla30_pg_logic23_and0[0]), .b(u_cla30_or54[0]), .out(u_cla30_or55));
  pg_logic pg_logic_u_cla30_pg_logic24_out(.a(a[24]), .b(b[24]), .pg_logic_or0(u_cla30_pg_logic24_or0), .pg_logic_and0(u_cla30_pg_logic24_and0), .pg_logic_xor0(u_cla30_pg_logic24_xor0));
  xor_gate xor_gate_u_cla30_xor24(.a(u_cla30_pg_logic24_xor0[0]), .b(u_cla30_or55[0]), .out(u_cla30_xor24));
  and_gate and_gate_u_cla30_and112(.a(u_cla30_or55[0]), .b(u_cla30_pg_logic24_or0[0]), .out(u_cla30_and112));
  or_gate or_gate_u_cla30_or56(.a(u_cla30_pg_logic24_and0[0]), .b(u_cla30_and112[0]), .out(u_cla30_or56));
  pg_logic pg_logic_u_cla30_pg_logic25_out(.a(a[25]), .b(b[25]), .pg_logic_or0(u_cla30_pg_logic25_or0), .pg_logic_and0(u_cla30_pg_logic25_and0), .pg_logic_xor0(u_cla30_pg_logic25_xor0));
  xor_gate xor_gate_u_cla30_xor25(.a(u_cla30_pg_logic25_xor0[0]), .b(u_cla30_or56[0]), .out(u_cla30_xor25));
  and_gate and_gate_u_cla30_and113(.a(u_cla30_or55[0]), .b(u_cla30_pg_logic25_or0[0]), .out(u_cla30_and113));
  and_gate and_gate_u_cla30_and114(.a(u_cla30_and113[0]), .b(u_cla30_pg_logic24_or0[0]), .out(u_cla30_and114));
  and_gate and_gate_u_cla30_and115(.a(u_cla30_pg_logic24_and0[0]), .b(u_cla30_pg_logic25_or0[0]), .out(u_cla30_and115));
  or_gate or_gate_u_cla30_or57(.a(u_cla30_and114[0]), .b(u_cla30_and115[0]), .out(u_cla30_or57));
  or_gate or_gate_u_cla30_or58(.a(u_cla30_pg_logic25_and0[0]), .b(u_cla30_or57[0]), .out(u_cla30_or58));
  pg_logic pg_logic_u_cla30_pg_logic26_out(.a(a[26]), .b(b[26]), .pg_logic_or0(u_cla30_pg_logic26_or0), .pg_logic_and0(u_cla30_pg_logic26_and0), .pg_logic_xor0(u_cla30_pg_logic26_xor0));
  xor_gate xor_gate_u_cla30_xor26(.a(u_cla30_pg_logic26_xor0[0]), .b(u_cla30_or58[0]), .out(u_cla30_xor26));
  and_gate and_gate_u_cla30_and116(.a(u_cla30_or55[0]), .b(u_cla30_pg_logic25_or0[0]), .out(u_cla30_and116));
  and_gate and_gate_u_cla30_and117(.a(u_cla30_pg_logic26_or0[0]), .b(u_cla30_pg_logic24_or0[0]), .out(u_cla30_and117));
  and_gate and_gate_u_cla30_and118(.a(u_cla30_and116[0]), .b(u_cla30_and117[0]), .out(u_cla30_and118));
  and_gate and_gate_u_cla30_and119(.a(u_cla30_pg_logic24_and0[0]), .b(u_cla30_pg_logic26_or0[0]), .out(u_cla30_and119));
  and_gate and_gate_u_cla30_and120(.a(u_cla30_and119[0]), .b(u_cla30_pg_logic25_or0[0]), .out(u_cla30_and120));
  and_gate and_gate_u_cla30_and121(.a(u_cla30_pg_logic25_and0[0]), .b(u_cla30_pg_logic26_or0[0]), .out(u_cla30_and121));
  or_gate or_gate_u_cla30_or59(.a(u_cla30_and118[0]), .b(u_cla30_and120[0]), .out(u_cla30_or59));
  or_gate or_gate_u_cla30_or60(.a(u_cla30_or59[0]), .b(u_cla30_and121[0]), .out(u_cla30_or60));
  or_gate or_gate_u_cla30_or61(.a(u_cla30_pg_logic26_and0[0]), .b(u_cla30_or60[0]), .out(u_cla30_or61));
  pg_logic pg_logic_u_cla30_pg_logic27_out(.a(a[27]), .b(b[27]), .pg_logic_or0(u_cla30_pg_logic27_or0), .pg_logic_and0(u_cla30_pg_logic27_and0), .pg_logic_xor0(u_cla30_pg_logic27_xor0));
  xor_gate xor_gate_u_cla30_xor27(.a(u_cla30_pg_logic27_xor0[0]), .b(u_cla30_or61[0]), .out(u_cla30_xor27));
  and_gate and_gate_u_cla30_and122(.a(u_cla30_or55[0]), .b(u_cla30_pg_logic26_or0[0]), .out(u_cla30_and122));
  and_gate and_gate_u_cla30_and123(.a(u_cla30_pg_logic27_or0[0]), .b(u_cla30_pg_logic25_or0[0]), .out(u_cla30_and123));
  and_gate and_gate_u_cla30_and124(.a(u_cla30_and122[0]), .b(u_cla30_and123[0]), .out(u_cla30_and124));
  and_gate and_gate_u_cla30_and125(.a(u_cla30_and124[0]), .b(u_cla30_pg_logic24_or0[0]), .out(u_cla30_and125));
  and_gate and_gate_u_cla30_and126(.a(u_cla30_pg_logic24_and0[0]), .b(u_cla30_pg_logic26_or0[0]), .out(u_cla30_and126));
  and_gate and_gate_u_cla30_and127(.a(u_cla30_pg_logic27_or0[0]), .b(u_cla30_pg_logic25_or0[0]), .out(u_cla30_and127));
  and_gate and_gate_u_cla30_and128(.a(u_cla30_and126[0]), .b(u_cla30_and127[0]), .out(u_cla30_and128));
  and_gate and_gate_u_cla30_and129(.a(u_cla30_pg_logic25_and0[0]), .b(u_cla30_pg_logic27_or0[0]), .out(u_cla30_and129));
  and_gate and_gate_u_cla30_and130(.a(u_cla30_and129[0]), .b(u_cla30_pg_logic26_or0[0]), .out(u_cla30_and130));
  and_gate and_gate_u_cla30_and131(.a(u_cla30_pg_logic26_and0[0]), .b(u_cla30_pg_logic27_or0[0]), .out(u_cla30_and131));
  or_gate or_gate_u_cla30_or62(.a(u_cla30_and125[0]), .b(u_cla30_and130[0]), .out(u_cla30_or62));
  or_gate or_gate_u_cla30_or63(.a(u_cla30_and128[0]), .b(u_cla30_and131[0]), .out(u_cla30_or63));
  or_gate or_gate_u_cla30_or64(.a(u_cla30_or62[0]), .b(u_cla30_or63[0]), .out(u_cla30_or64));
  or_gate or_gate_u_cla30_or65(.a(u_cla30_pg_logic27_and0[0]), .b(u_cla30_or64[0]), .out(u_cla30_or65));
  pg_logic pg_logic_u_cla30_pg_logic28_out(.a(a[28]), .b(b[28]), .pg_logic_or0(u_cla30_pg_logic28_or0), .pg_logic_and0(u_cla30_pg_logic28_and0), .pg_logic_xor0(u_cla30_pg_logic28_xor0));
  xor_gate xor_gate_u_cla30_xor28(.a(u_cla30_pg_logic28_xor0[0]), .b(u_cla30_or65[0]), .out(u_cla30_xor28));
  and_gate and_gate_u_cla30_and132(.a(u_cla30_or65[0]), .b(u_cla30_pg_logic28_or0[0]), .out(u_cla30_and132));
  or_gate or_gate_u_cla30_or66(.a(u_cla30_pg_logic28_and0[0]), .b(u_cla30_and132[0]), .out(u_cla30_or66));
  pg_logic pg_logic_u_cla30_pg_logic29_out(.a(a[29]), .b(b[29]), .pg_logic_or0(u_cla30_pg_logic29_or0), .pg_logic_and0(u_cla30_pg_logic29_and0), .pg_logic_xor0(u_cla30_pg_logic29_xor0));
  xor_gate xor_gate_u_cla30_xor29(.a(u_cla30_pg_logic29_xor0[0]), .b(u_cla30_or66[0]), .out(u_cla30_xor29));
  and_gate and_gate_u_cla30_and133(.a(u_cla30_or65[0]), .b(u_cla30_pg_logic29_or0[0]), .out(u_cla30_and133));
  and_gate and_gate_u_cla30_and134(.a(u_cla30_and133[0]), .b(u_cla30_pg_logic28_or0[0]), .out(u_cla30_and134));
  and_gate and_gate_u_cla30_and135(.a(u_cla30_pg_logic28_and0[0]), .b(u_cla30_pg_logic29_or0[0]), .out(u_cla30_and135));
  or_gate or_gate_u_cla30_or67(.a(u_cla30_and134[0]), .b(u_cla30_and135[0]), .out(u_cla30_or67));
  or_gate or_gate_u_cla30_or68(.a(u_cla30_pg_logic29_and0[0]), .b(u_cla30_or67[0]), .out(u_cla30_or68));

  assign u_cla30_out[0] = u_cla30_pg_logic0_xor0[0];
  assign u_cla30_out[1] = u_cla30_xor1[0];
  assign u_cla30_out[2] = u_cla30_xor2[0];
  assign u_cla30_out[3] = u_cla30_xor3[0];
  assign u_cla30_out[4] = u_cla30_xor4[0];
  assign u_cla30_out[5] = u_cla30_xor5[0];
  assign u_cla30_out[6] = u_cla30_xor6[0];
  assign u_cla30_out[7] = u_cla30_xor7[0];
  assign u_cla30_out[8] = u_cla30_xor8[0];
  assign u_cla30_out[9] = u_cla30_xor9[0];
  assign u_cla30_out[10] = u_cla30_xor10[0];
  assign u_cla30_out[11] = u_cla30_xor11[0];
  assign u_cla30_out[12] = u_cla30_xor12[0];
  assign u_cla30_out[13] = u_cla30_xor13[0];
  assign u_cla30_out[14] = u_cla30_xor14[0];
  assign u_cla30_out[15] = u_cla30_xor15[0];
  assign u_cla30_out[16] = u_cla30_xor16[0];
  assign u_cla30_out[17] = u_cla30_xor17[0];
  assign u_cla30_out[18] = u_cla30_xor18[0];
  assign u_cla30_out[19] = u_cla30_xor19[0];
  assign u_cla30_out[20] = u_cla30_xor20[0];
  assign u_cla30_out[21] = u_cla30_xor21[0];
  assign u_cla30_out[22] = u_cla30_xor22[0];
  assign u_cla30_out[23] = u_cla30_xor23[0];
  assign u_cla30_out[24] = u_cla30_xor24[0];
  assign u_cla30_out[25] = u_cla30_xor25[0];
  assign u_cla30_out[26] = u_cla30_xor26[0];
  assign u_cla30_out[27] = u_cla30_xor27[0];
  assign u_cla30_out[28] = u_cla30_xor28[0];
  assign u_cla30_out[29] = u_cla30_xor29[0];
  assign u_cla30_out[30] = u_cla30_or68[0];
endmodule

module h_u_wallace_cla16(input [15:0] a, input [15:0] b, output [31:0] h_u_wallace_cla16_out);
  wire [0:0] h_u_wallace_cla16_and_2_0;
  wire [0:0] h_u_wallace_cla16_and_1_1;
  wire [0:0] h_u_wallace_cla16_ha0_xor0;
  wire [0:0] h_u_wallace_cla16_ha0_and0;
  wire [0:0] h_u_wallace_cla16_and_3_0;
  wire [0:0] h_u_wallace_cla16_and_2_1;
  wire [0:0] h_u_wallace_cla16_fa0_xor1;
  wire [0:0] h_u_wallace_cla16_fa0_or0;
  wire [0:0] h_u_wallace_cla16_and_4_0;
  wire [0:0] h_u_wallace_cla16_and_3_1;
  wire [0:0] h_u_wallace_cla16_fa1_xor1;
  wire [0:0] h_u_wallace_cla16_fa1_or0;
  wire [0:0] h_u_wallace_cla16_and_5_0;
  wire [0:0] h_u_wallace_cla16_and_4_1;
  wire [0:0] h_u_wallace_cla16_fa2_xor1;
  wire [0:0] h_u_wallace_cla16_fa2_or0;
  wire [0:0] h_u_wallace_cla16_and_6_0;
  wire [0:0] h_u_wallace_cla16_and_5_1;
  wire [0:0] h_u_wallace_cla16_fa3_xor1;
  wire [0:0] h_u_wallace_cla16_fa3_or0;
  wire [0:0] h_u_wallace_cla16_and_7_0;
  wire [0:0] h_u_wallace_cla16_and_6_1;
  wire [0:0] h_u_wallace_cla16_fa4_xor1;
  wire [0:0] h_u_wallace_cla16_fa4_or0;
  wire [0:0] h_u_wallace_cla16_and_8_0;
  wire [0:0] h_u_wallace_cla16_and_7_1;
  wire [0:0] h_u_wallace_cla16_fa5_xor1;
  wire [0:0] h_u_wallace_cla16_fa5_or0;
  wire [0:0] h_u_wallace_cla16_and_9_0;
  wire [0:0] h_u_wallace_cla16_and_8_1;
  wire [0:0] h_u_wallace_cla16_fa6_xor1;
  wire [0:0] h_u_wallace_cla16_fa6_or0;
  wire [0:0] h_u_wallace_cla16_and_10_0;
  wire [0:0] h_u_wallace_cla16_and_9_1;
  wire [0:0] h_u_wallace_cla16_fa7_xor1;
  wire [0:0] h_u_wallace_cla16_fa7_or0;
  wire [0:0] h_u_wallace_cla16_and_11_0;
  wire [0:0] h_u_wallace_cla16_and_10_1;
  wire [0:0] h_u_wallace_cla16_fa8_xor1;
  wire [0:0] h_u_wallace_cla16_fa8_or0;
  wire [0:0] h_u_wallace_cla16_and_12_0;
  wire [0:0] h_u_wallace_cla16_and_11_1;
  wire [0:0] h_u_wallace_cla16_fa9_xor1;
  wire [0:0] h_u_wallace_cla16_fa9_or0;
  wire [0:0] h_u_wallace_cla16_and_13_0;
  wire [0:0] h_u_wallace_cla16_and_12_1;
  wire [0:0] h_u_wallace_cla16_fa10_xor1;
  wire [0:0] h_u_wallace_cla16_fa10_or0;
  wire [0:0] h_u_wallace_cla16_and_14_0;
  wire [0:0] h_u_wallace_cla16_and_13_1;
  wire [0:0] h_u_wallace_cla16_fa11_xor1;
  wire [0:0] h_u_wallace_cla16_fa11_or0;
  wire [0:0] h_u_wallace_cla16_and_15_0;
  wire [0:0] h_u_wallace_cla16_and_14_1;
  wire [0:0] h_u_wallace_cla16_fa12_xor1;
  wire [0:0] h_u_wallace_cla16_fa12_or0;
  wire [0:0] h_u_wallace_cla16_and_15_1;
  wire [0:0] h_u_wallace_cla16_and_14_2;
  wire [0:0] h_u_wallace_cla16_fa13_xor1;
  wire [0:0] h_u_wallace_cla16_fa13_or0;
  wire [0:0] h_u_wallace_cla16_and_15_2;
  wire [0:0] h_u_wallace_cla16_and_14_3;
  wire [0:0] h_u_wallace_cla16_fa14_xor1;
  wire [0:0] h_u_wallace_cla16_fa14_or0;
  wire [0:0] h_u_wallace_cla16_and_15_3;
  wire [0:0] h_u_wallace_cla16_and_14_4;
  wire [0:0] h_u_wallace_cla16_fa15_xor1;
  wire [0:0] h_u_wallace_cla16_fa15_or0;
  wire [0:0] h_u_wallace_cla16_and_15_4;
  wire [0:0] h_u_wallace_cla16_and_14_5;
  wire [0:0] h_u_wallace_cla16_fa16_xor1;
  wire [0:0] h_u_wallace_cla16_fa16_or0;
  wire [0:0] h_u_wallace_cla16_and_15_5;
  wire [0:0] h_u_wallace_cla16_and_14_6;
  wire [0:0] h_u_wallace_cla16_fa17_xor1;
  wire [0:0] h_u_wallace_cla16_fa17_or0;
  wire [0:0] h_u_wallace_cla16_and_15_6;
  wire [0:0] h_u_wallace_cla16_and_14_7;
  wire [0:0] h_u_wallace_cla16_fa18_xor1;
  wire [0:0] h_u_wallace_cla16_fa18_or0;
  wire [0:0] h_u_wallace_cla16_and_15_7;
  wire [0:0] h_u_wallace_cla16_and_14_8;
  wire [0:0] h_u_wallace_cla16_fa19_xor1;
  wire [0:0] h_u_wallace_cla16_fa19_or0;
  wire [0:0] h_u_wallace_cla16_and_15_8;
  wire [0:0] h_u_wallace_cla16_and_14_9;
  wire [0:0] h_u_wallace_cla16_fa20_xor1;
  wire [0:0] h_u_wallace_cla16_fa20_or0;
  wire [0:0] h_u_wallace_cla16_and_15_9;
  wire [0:0] h_u_wallace_cla16_and_14_10;
  wire [0:0] h_u_wallace_cla16_fa21_xor1;
  wire [0:0] h_u_wallace_cla16_fa21_or0;
  wire [0:0] h_u_wallace_cla16_and_15_10;
  wire [0:0] h_u_wallace_cla16_and_14_11;
  wire [0:0] h_u_wallace_cla16_fa22_xor1;
  wire [0:0] h_u_wallace_cla16_fa22_or0;
  wire [0:0] h_u_wallace_cla16_and_15_11;
  wire [0:0] h_u_wallace_cla16_and_14_12;
  wire [0:0] h_u_wallace_cla16_fa23_xor1;
  wire [0:0] h_u_wallace_cla16_fa23_or0;
  wire [0:0] h_u_wallace_cla16_and_15_12;
  wire [0:0] h_u_wallace_cla16_and_14_13;
  wire [0:0] h_u_wallace_cla16_fa24_xor1;
  wire [0:0] h_u_wallace_cla16_fa24_or0;
  wire [0:0] h_u_wallace_cla16_and_15_13;
  wire [0:0] h_u_wallace_cla16_and_14_14;
  wire [0:0] h_u_wallace_cla16_fa25_xor1;
  wire [0:0] h_u_wallace_cla16_fa25_or0;
  wire [0:0] h_u_wallace_cla16_and_1_2;
  wire [0:0] h_u_wallace_cla16_and_0_3;
  wire [0:0] h_u_wallace_cla16_ha1_xor0;
  wire [0:0] h_u_wallace_cla16_ha1_and0;
  wire [0:0] h_u_wallace_cla16_and_2_2;
  wire [0:0] h_u_wallace_cla16_and_1_3;
  wire [0:0] h_u_wallace_cla16_fa26_xor1;
  wire [0:0] h_u_wallace_cla16_fa26_or0;
  wire [0:0] h_u_wallace_cla16_and_3_2;
  wire [0:0] h_u_wallace_cla16_and_2_3;
  wire [0:0] h_u_wallace_cla16_fa27_xor1;
  wire [0:0] h_u_wallace_cla16_fa27_or0;
  wire [0:0] h_u_wallace_cla16_and_4_2;
  wire [0:0] h_u_wallace_cla16_and_3_3;
  wire [0:0] h_u_wallace_cla16_fa28_xor1;
  wire [0:0] h_u_wallace_cla16_fa28_or0;
  wire [0:0] h_u_wallace_cla16_and_5_2;
  wire [0:0] h_u_wallace_cla16_and_4_3;
  wire [0:0] h_u_wallace_cla16_fa29_xor1;
  wire [0:0] h_u_wallace_cla16_fa29_or0;
  wire [0:0] h_u_wallace_cla16_and_6_2;
  wire [0:0] h_u_wallace_cla16_and_5_3;
  wire [0:0] h_u_wallace_cla16_fa30_xor1;
  wire [0:0] h_u_wallace_cla16_fa30_or0;
  wire [0:0] h_u_wallace_cla16_and_7_2;
  wire [0:0] h_u_wallace_cla16_and_6_3;
  wire [0:0] h_u_wallace_cla16_fa31_xor1;
  wire [0:0] h_u_wallace_cla16_fa31_or0;
  wire [0:0] h_u_wallace_cla16_and_8_2;
  wire [0:0] h_u_wallace_cla16_and_7_3;
  wire [0:0] h_u_wallace_cla16_fa32_xor1;
  wire [0:0] h_u_wallace_cla16_fa32_or0;
  wire [0:0] h_u_wallace_cla16_and_9_2;
  wire [0:0] h_u_wallace_cla16_and_8_3;
  wire [0:0] h_u_wallace_cla16_fa33_xor1;
  wire [0:0] h_u_wallace_cla16_fa33_or0;
  wire [0:0] h_u_wallace_cla16_and_10_2;
  wire [0:0] h_u_wallace_cla16_and_9_3;
  wire [0:0] h_u_wallace_cla16_fa34_xor1;
  wire [0:0] h_u_wallace_cla16_fa34_or0;
  wire [0:0] h_u_wallace_cla16_and_11_2;
  wire [0:0] h_u_wallace_cla16_and_10_3;
  wire [0:0] h_u_wallace_cla16_fa35_xor1;
  wire [0:0] h_u_wallace_cla16_fa35_or0;
  wire [0:0] h_u_wallace_cla16_and_12_2;
  wire [0:0] h_u_wallace_cla16_and_11_3;
  wire [0:0] h_u_wallace_cla16_fa36_xor1;
  wire [0:0] h_u_wallace_cla16_fa36_or0;
  wire [0:0] h_u_wallace_cla16_and_13_2;
  wire [0:0] h_u_wallace_cla16_and_12_3;
  wire [0:0] h_u_wallace_cla16_fa37_xor1;
  wire [0:0] h_u_wallace_cla16_fa37_or0;
  wire [0:0] h_u_wallace_cla16_and_13_3;
  wire [0:0] h_u_wallace_cla16_and_12_4;
  wire [0:0] h_u_wallace_cla16_fa38_xor1;
  wire [0:0] h_u_wallace_cla16_fa38_or0;
  wire [0:0] h_u_wallace_cla16_and_13_4;
  wire [0:0] h_u_wallace_cla16_and_12_5;
  wire [0:0] h_u_wallace_cla16_fa39_xor1;
  wire [0:0] h_u_wallace_cla16_fa39_or0;
  wire [0:0] h_u_wallace_cla16_and_13_5;
  wire [0:0] h_u_wallace_cla16_and_12_6;
  wire [0:0] h_u_wallace_cla16_fa40_xor1;
  wire [0:0] h_u_wallace_cla16_fa40_or0;
  wire [0:0] h_u_wallace_cla16_and_13_6;
  wire [0:0] h_u_wallace_cla16_and_12_7;
  wire [0:0] h_u_wallace_cla16_fa41_xor1;
  wire [0:0] h_u_wallace_cla16_fa41_or0;
  wire [0:0] h_u_wallace_cla16_and_13_7;
  wire [0:0] h_u_wallace_cla16_and_12_8;
  wire [0:0] h_u_wallace_cla16_fa42_xor1;
  wire [0:0] h_u_wallace_cla16_fa42_or0;
  wire [0:0] h_u_wallace_cla16_and_13_8;
  wire [0:0] h_u_wallace_cla16_and_12_9;
  wire [0:0] h_u_wallace_cla16_fa43_xor1;
  wire [0:0] h_u_wallace_cla16_fa43_or0;
  wire [0:0] h_u_wallace_cla16_and_13_9;
  wire [0:0] h_u_wallace_cla16_and_12_10;
  wire [0:0] h_u_wallace_cla16_fa44_xor1;
  wire [0:0] h_u_wallace_cla16_fa44_or0;
  wire [0:0] h_u_wallace_cla16_and_13_10;
  wire [0:0] h_u_wallace_cla16_and_12_11;
  wire [0:0] h_u_wallace_cla16_fa45_xor1;
  wire [0:0] h_u_wallace_cla16_fa45_or0;
  wire [0:0] h_u_wallace_cla16_and_13_11;
  wire [0:0] h_u_wallace_cla16_and_12_12;
  wire [0:0] h_u_wallace_cla16_fa46_xor1;
  wire [0:0] h_u_wallace_cla16_fa46_or0;
  wire [0:0] h_u_wallace_cla16_and_13_12;
  wire [0:0] h_u_wallace_cla16_and_12_13;
  wire [0:0] h_u_wallace_cla16_fa47_xor1;
  wire [0:0] h_u_wallace_cla16_fa47_or0;
  wire [0:0] h_u_wallace_cla16_and_13_13;
  wire [0:0] h_u_wallace_cla16_and_12_14;
  wire [0:0] h_u_wallace_cla16_fa48_xor1;
  wire [0:0] h_u_wallace_cla16_fa48_or0;
  wire [0:0] h_u_wallace_cla16_and_13_14;
  wire [0:0] h_u_wallace_cla16_and_12_15;
  wire [0:0] h_u_wallace_cla16_fa49_xor1;
  wire [0:0] h_u_wallace_cla16_fa49_or0;
  wire [0:0] h_u_wallace_cla16_and_0_4;
  wire [0:0] h_u_wallace_cla16_ha2_xor0;
  wire [0:0] h_u_wallace_cla16_ha2_and0;
  wire [0:0] h_u_wallace_cla16_and_1_4;
  wire [0:0] h_u_wallace_cla16_and_0_5;
  wire [0:0] h_u_wallace_cla16_fa50_xor1;
  wire [0:0] h_u_wallace_cla16_fa50_or0;
  wire [0:0] h_u_wallace_cla16_and_2_4;
  wire [0:0] h_u_wallace_cla16_and_1_5;
  wire [0:0] h_u_wallace_cla16_fa51_xor1;
  wire [0:0] h_u_wallace_cla16_fa51_or0;
  wire [0:0] h_u_wallace_cla16_and_3_4;
  wire [0:0] h_u_wallace_cla16_and_2_5;
  wire [0:0] h_u_wallace_cla16_fa52_xor1;
  wire [0:0] h_u_wallace_cla16_fa52_or0;
  wire [0:0] h_u_wallace_cla16_and_4_4;
  wire [0:0] h_u_wallace_cla16_and_3_5;
  wire [0:0] h_u_wallace_cla16_fa53_xor1;
  wire [0:0] h_u_wallace_cla16_fa53_or0;
  wire [0:0] h_u_wallace_cla16_and_5_4;
  wire [0:0] h_u_wallace_cla16_and_4_5;
  wire [0:0] h_u_wallace_cla16_fa54_xor1;
  wire [0:0] h_u_wallace_cla16_fa54_or0;
  wire [0:0] h_u_wallace_cla16_and_6_4;
  wire [0:0] h_u_wallace_cla16_and_5_5;
  wire [0:0] h_u_wallace_cla16_fa55_xor1;
  wire [0:0] h_u_wallace_cla16_fa55_or0;
  wire [0:0] h_u_wallace_cla16_and_7_4;
  wire [0:0] h_u_wallace_cla16_and_6_5;
  wire [0:0] h_u_wallace_cla16_fa56_xor1;
  wire [0:0] h_u_wallace_cla16_fa56_or0;
  wire [0:0] h_u_wallace_cla16_and_8_4;
  wire [0:0] h_u_wallace_cla16_and_7_5;
  wire [0:0] h_u_wallace_cla16_fa57_xor1;
  wire [0:0] h_u_wallace_cla16_fa57_or0;
  wire [0:0] h_u_wallace_cla16_and_9_4;
  wire [0:0] h_u_wallace_cla16_and_8_5;
  wire [0:0] h_u_wallace_cla16_fa58_xor1;
  wire [0:0] h_u_wallace_cla16_fa58_or0;
  wire [0:0] h_u_wallace_cla16_and_10_4;
  wire [0:0] h_u_wallace_cla16_and_9_5;
  wire [0:0] h_u_wallace_cla16_fa59_xor1;
  wire [0:0] h_u_wallace_cla16_fa59_or0;
  wire [0:0] h_u_wallace_cla16_and_11_4;
  wire [0:0] h_u_wallace_cla16_and_10_5;
  wire [0:0] h_u_wallace_cla16_fa60_xor1;
  wire [0:0] h_u_wallace_cla16_fa60_or0;
  wire [0:0] h_u_wallace_cla16_and_11_5;
  wire [0:0] h_u_wallace_cla16_and_10_6;
  wire [0:0] h_u_wallace_cla16_fa61_xor1;
  wire [0:0] h_u_wallace_cla16_fa61_or0;
  wire [0:0] h_u_wallace_cla16_and_11_6;
  wire [0:0] h_u_wallace_cla16_and_10_7;
  wire [0:0] h_u_wallace_cla16_fa62_xor1;
  wire [0:0] h_u_wallace_cla16_fa62_or0;
  wire [0:0] h_u_wallace_cla16_and_11_7;
  wire [0:0] h_u_wallace_cla16_and_10_8;
  wire [0:0] h_u_wallace_cla16_fa63_xor1;
  wire [0:0] h_u_wallace_cla16_fa63_or0;
  wire [0:0] h_u_wallace_cla16_and_11_8;
  wire [0:0] h_u_wallace_cla16_and_10_9;
  wire [0:0] h_u_wallace_cla16_fa64_xor1;
  wire [0:0] h_u_wallace_cla16_fa64_or0;
  wire [0:0] h_u_wallace_cla16_and_11_9;
  wire [0:0] h_u_wallace_cla16_and_10_10;
  wire [0:0] h_u_wallace_cla16_fa65_xor1;
  wire [0:0] h_u_wallace_cla16_fa65_or0;
  wire [0:0] h_u_wallace_cla16_and_11_10;
  wire [0:0] h_u_wallace_cla16_and_10_11;
  wire [0:0] h_u_wallace_cla16_fa66_xor1;
  wire [0:0] h_u_wallace_cla16_fa66_or0;
  wire [0:0] h_u_wallace_cla16_and_11_11;
  wire [0:0] h_u_wallace_cla16_and_10_12;
  wire [0:0] h_u_wallace_cla16_fa67_xor1;
  wire [0:0] h_u_wallace_cla16_fa67_or0;
  wire [0:0] h_u_wallace_cla16_and_11_12;
  wire [0:0] h_u_wallace_cla16_and_10_13;
  wire [0:0] h_u_wallace_cla16_fa68_xor1;
  wire [0:0] h_u_wallace_cla16_fa68_or0;
  wire [0:0] h_u_wallace_cla16_and_11_13;
  wire [0:0] h_u_wallace_cla16_and_10_14;
  wire [0:0] h_u_wallace_cla16_fa69_xor1;
  wire [0:0] h_u_wallace_cla16_fa69_or0;
  wire [0:0] h_u_wallace_cla16_and_11_14;
  wire [0:0] h_u_wallace_cla16_and_10_15;
  wire [0:0] h_u_wallace_cla16_fa70_xor1;
  wire [0:0] h_u_wallace_cla16_fa70_or0;
  wire [0:0] h_u_wallace_cla16_and_11_15;
  wire [0:0] h_u_wallace_cla16_fa71_xor1;
  wire [0:0] h_u_wallace_cla16_fa71_or0;
  wire [0:0] h_u_wallace_cla16_ha3_xor0;
  wire [0:0] h_u_wallace_cla16_ha3_and0;
  wire [0:0] h_u_wallace_cla16_and_0_6;
  wire [0:0] h_u_wallace_cla16_fa72_xor1;
  wire [0:0] h_u_wallace_cla16_fa72_or0;
  wire [0:0] h_u_wallace_cla16_and_1_6;
  wire [0:0] h_u_wallace_cla16_and_0_7;
  wire [0:0] h_u_wallace_cla16_fa73_xor1;
  wire [0:0] h_u_wallace_cla16_fa73_or0;
  wire [0:0] h_u_wallace_cla16_and_2_6;
  wire [0:0] h_u_wallace_cla16_and_1_7;
  wire [0:0] h_u_wallace_cla16_fa74_xor1;
  wire [0:0] h_u_wallace_cla16_fa74_or0;
  wire [0:0] h_u_wallace_cla16_and_3_6;
  wire [0:0] h_u_wallace_cla16_and_2_7;
  wire [0:0] h_u_wallace_cla16_fa75_xor1;
  wire [0:0] h_u_wallace_cla16_fa75_or0;
  wire [0:0] h_u_wallace_cla16_and_4_6;
  wire [0:0] h_u_wallace_cla16_and_3_7;
  wire [0:0] h_u_wallace_cla16_fa76_xor1;
  wire [0:0] h_u_wallace_cla16_fa76_or0;
  wire [0:0] h_u_wallace_cla16_and_5_6;
  wire [0:0] h_u_wallace_cla16_and_4_7;
  wire [0:0] h_u_wallace_cla16_fa77_xor1;
  wire [0:0] h_u_wallace_cla16_fa77_or0;
  wire [0:0] h_u_wallace_cla16_and_6_6;
  wire [0:0] h_u_wallace_cla16_and_5_7;
  wire [0:0] h_u_wallace_cla16_fa78_xor1;
  wire [0:0] h_u_wallace_cla16_fa78_or0;
  wire [0:0] h_u_wallace_cla16_and_7_6;
  wire [0:0] h_u_wallace_cla16_and_6_7;
  wire [0:0] h_u_wallace_cla16_fa79_xor1;
  wire [0:0] h_u_wallace_cla16_fa79_or0;
  wire [0:0] h_u_wallace_cla16_and_8_6;
  wire [0:0] h_u_wallace_cla16_and_7_7;
  wire [0:0] h_u_wallace_cla16_fa80_xor1;
  wire [0:0] h_u_wallace_cla16_fa80_or0;
  wire [0:0] h_u_wallace_cla16_and_9_6;
  wire [0:0] h_u_wallace_cla16_and_8_7;
  wire [0:0] h_u_wallace_cla16_fa81_xor1;
  wire [0:0] h_u_wallace_cla16_fa81_or0;
  wire [0:0] h_u_wallace_cla16_and_9_7;
  wire [0:0] h_u_wallace_cla16_and_8_8;
  wire [0:0] h_u_wallace_cla16_fa82_xor1;
  wire [0:0] h_u_wallace_cla16_fa82_or0;
  wire [0:0] h_u_wallace_cla16_and_9_8;
  wire [0:0] h_u_wallace_cla16_and_8_9;
  wire [0:0] h_u_wallace_cla16_fa83_xor1;
  wire [0:0] h_u_wallace_cla16_fa83_or0;
  wire [0:0] h_u_wallace_cla16_and_9_9;
  wire [0:0] h_u_wallace_cla16_and_8_10;
  wire [0:0] h_u_wallace_cla16_fa84_xor1;
  wire [0:0] h_u_wallace_cla16_fa84_or0;
  wire [0:0] h_u_wallace_cla16_and_9_10;
  wire [0:0] h_u_wallace_cla16_and_8_11;
  wire [0:0] h_u_wallace_cla16_fa85_xor1;
  wire [0:0] h_u_wallace_cla16_fa85_or0;
  wire [0:0] h_u_wallace_cla16_and_9_11;
  wire [0:0] h_u_wallace_cla16_and_8_12;
  wire [0:0] h_u_wallace_cla16_fa86_xor1;
  wire [0:0] h_u_wallace_cla16_fa86_or0;
  wire [0:0] h_u_wallace_cla16_and_9_12;
  wire [0:0] h_u_wallace_cla16_and_8_13;
  wire [0:0] h_u_wallace_cla16_fa87_xor1;
  wire [0:0] h_u_wallace_cla16_fa87_or0;
  wire [0:0] h_u_wallace_cla16_and_9_13;
  wire [0:0] h_u_wallace_cla16_and_8_14;
  wire [0:0] h_u_wallace_cla16_fa88_xor1;
  wire [0:0] h_u_wallace_cla16_fa88_or0;
  wire [0:0] h_u_wallace_cla16_and_9_14;
  wire [0:0] h_u_wallace_cla16_and_8_15;
  wire [0:0] h_u_wallace_cla16_fa89_xor1;
  wire [0:0] h_u_wallace_cla16_fa89_or0;
  wire [0:0] h_u_wallace_cla16_and_9_15;
  wire [0:0] h_u_wallace_cla16_fa90_xor1;
  wire [0:0] h_u_wallace_cla16_fa90_or0;
  wire [0:0] h_u_wallace_cla16_fa91_xor1;
  wire [0:0] h_u_wallace_cla16_fa91_or0;
  wire [0:0] h_u_wallace_cla16_ha4_xor0;
  wire [0:0] h_u_wallace_cla16_ha4_and0;
  wire [0:0] h_u_wallace_cla16_fa92_xor1;
  wire [0:0] h_u_wallace_cla16_fa92_or0;
  wire [0:0] h_u_wallace_cla16_and_0_8;
  wire [0:0] h_u_wallace_cla16_fa93_xor1;
  wire [0:0] h_u_wallace_cla16_fa93_or0;
  wire [0:0] h_u_wallace_cla16_and_1_8;
  wire [0:0] h_u_wallace_cla16_and_0_9;
  wire [0:0] h_u_wallace_cla16_fa94_xor1;
  wire [0:0] h_u_wallace_cla16_fa94_or0;
  wire [0:0] h_u_wallace_cla16_and_2_8;
  wire [0:0] h_u_wallace_cla16_and_1_9;
  wire [0:0] h_u_wallace_cla16_fa95_xor1;
  wire [0:0] h_u_wallace_cla16_fa95_or0;
  wire [0:0] h_u_wallace_cla16_and_3_8;
  wire [0:0] h_u_wallace_cla16_and_2_9;
  wire [0:0] h_u_wallace_cla16_fa96_xor1;
  wire [0:0] h_u_wallace_cla16_fa96_or0;
  wire [0:0] h_u_wallace_cla16_and_4_8;
  wire [0:0] h_u_wallace_cla16_and_3_9;
  wire [0:0] h_u_wallace_cla16_fa97_xor1;
  wire [0:0] h_u_wallace_cla16_fa97_or0;
  wire [0:0] h_u_wallace_cla16_and_5_8;
  wire [0:0] h_u_wallace_cla16_and_4_9;
  wire [0:0] h_u_wallace_cla16_fa98_xor1;
  wire [0:0] h_u_wallace_cla16_fa98_or0;
  wire [0:0] h_u_wallace_cla16_and_6_8;
  wire [0:0] h_u_wallace_cla16_and_5_9;
  wire [0:0] h_u_wallace_cla16_fa99_xor1;
  wire [0:0] h_u_wallace_cla16_fa99_or0;
  wire [0:0] h_u_wallace_cla16_and_7_8;
  wire [0:0] h_u_wallace_cla16_and_6_9;
  wire [0:0] h_u_wallace_cla16_fa100_xor1;
  wire [0:0] h_u_wallace_cla16_fa100_or0;
  wire [0:0] h_u_wallace_cla16_and_7_9;
  wire [0:0] h_u_wallace_cla16_and_6_10;
  wire [0:0] h_u_wallace_cla16_fa101_xor1;
  wire [0:0] h_u_wallace_cla16_fa101_or0;
  wire [0:0] h_u_wallace_cla16_and_7_10;
  wire [0:0] h_u_wallace_cla16_and_6_11;
  wire [0:0] h_u_wallace_cla16_fa102_xor1;
  wire [0:0] h_u_wallace_cla16_fa102_or0;
  wire [0:0] h_u_wallace_cla16_and_7_11;
  wire [0:0] h_u_wallace_cla16_and_6_12;
  wire [0:0] h_u_wallace_cla16_fa103_xor1;
  wire [0:0] h_u_wallace_cla16_fa103_or0;
  wire [0:0] h_u_wallace_cla16_and_7_12;
  wire [0:0] h_u_wallace_cla16_and_6_13;
  wire [0:0] h_u_wallace_cla16_fa104_xor1;
  wire [0:0] h_u_wallace_cla16_fa104_or0;
  wire [0:0] h_u_wallace_cla16_and_7_13;
  wire [0:0] h_u_wallace_cla16_and_6_14;
  wire [0:0] h_u_wallace_cla16_fa105_xor1;
  wire [0:0] h_u_wallace_cla16_fa105_or0;
  wire [0:0] h_u_wallace_cla16_and_7_14;
  wire [0:0] h_u_wallace_cla16_and_6_15;
  wire [0:0] h_u_wallace_cla16_fa106_xor1;
  wire [0:0] h_u_wallace_cla16_fa106_or0;
  wire [0:0] h_u_wallace_cla16_and_7_15;
  wire [0:0] h_u_wallace_cla16_fa107_xor1;
  wire [0:0] h_u_wallace_cla16_fa107_or0;
  wire [0:0] h_u_wallace_cla16_fa108_xor1;
  wire [0:0] h_u_wallace_cla16_fa108_or0;
  wire [0:0] h_u_wallace_cla16_fa109_xor1;
  wire [0:0] h_u_wallace_cla16_fa109_or0;
  wire [0:0] h_u_wallace_cla16_ha5_xor0;
  wire [0:0] h_u_wallace_cla16_ha5_and0;
  wire [0:0] h_u_wallace_cla16_fa110_xor1;
  wire [0:0] h_u_wallace_cla16_fa110_or0;
  wire [0:0] h_u_wallace_cla16_fa111_xor1;
  wire [0:0] h_u_wallace_cla16_fa111_or0;
  wire [0:0] h_u_wallace_cla16_and_0_10;
  wire [0:0] h_u_wallace_cla16_fa112_xor1;
  wire [0:0] h_u_wallace_cla16_fa112_or0;
  wire [0:0] h_u_wallace_cla16_and_1_10;
  wire [0:0] h_u_wallace_cla16_and_0_11;
  wire [0:0] h_u_wallace_cla16_fa113_xor1;
  wire [0:0] h_u_wallace_cla16_fa113_or0;
  wire [0:0] h_u_wallace_cla16_and_2_10;
  wire [0:0] h_u_wallace_cla16_and_1_11;
  wire [0:0] h_u_wallace_cla16_fa114_xor1;
  wire [0:0] h_u_wallace_cla16_fa114_or0;
  wire [0:0] h_u_wallace_cla16_and_3_10;
  wire [0:0] h_u_wallace_cla16_and_2_11;
  wire [0:0] h_u_wallace_cla16_fa115_xor1;
  wire [0:0] h_u_wallace_cla16_fa115_or0;
  wire [0:0] h_u_wallace_cla16_and_4_10;
  wire [0:0] h_u_wallace_cla16_and_3_11;
  wire [0:0] h_u_wallace_cla16_fa116_xor1;
  wire [0:0] h_u_wallace_cla16_fa116_or0;
  wire [0:0] h_u_wallace_cla16_and_5_10;
  wire [0:0] h_u_wallace_cla16_and_4_11;
  wire [0:0] h_u_wallace_cla16_fa117_xor1;
  wire [0:0] h_u_wallace_cla16_fa117_or0;
  wire [0:0] h_u_wallace_cla16_and_5_11;
  wire [0:0] h_u_wallace_cla16_and_4_12;
  wire [0:0] h_u_wallace_cla16_fa118_xor1;
  wire [0:0] h_u_wallace_cla16_fa118_or0;
  wire [0:0] h_u_wallace_cla16_and_5_12;
  wire [0:0] h_u_wallace_cla16_and_4_13;
  wire [0:0] h_u_wallace_cla16_fa119_xor1;
  wire [0:0] h_u_wallace_cla16_fa119_or0;
  wire [0:0] h_u_wallace_cla16_and_5_13;
  wire [0:0] h_u_wallace_cla16_and_4_14;
  wire [0:0] h_u_wallace_cla16_fa120_xor1;
  wire [0:0] h_u_wallace_cla16_fa120_or0;
  wire [0:0] h_u_wallace_cla16_and_5_14;
  wire [0:0] h_u_wallace_cla16_and_4_15;
  wire [0:0] h_u_wallace_cla16_fa121_xor1;
  wire [0:0] h_u_wallace_cla16_fa121_or0;
  wire [0:0] h_u_wallace_cla16_and_5_15;
  wire [0:0] h_u_wallace_cla16_fa122_xor1;
  wire [0:0] h_u_wallace_cla16_fa122_or0;
  wire [0:0] h_u_wallace_cla16_fa123_xor1;
  wire [0:0] h_u_wallace_cla16_fa123_or0;
  wire [0:0] h_u_wallace_cla16_fa124_xor1;
  wire [0:0] h_u_wallace_cla16_fa124_or0;
  wire [0:0] h_u_wallace_cla16_fa125_xor1;
  wire [0:0] h_u_wallace_cla16_fa125_or0;
  wire [0:0] h_u_wallace_cla16_ha6_xor0;
  wire [0:0] h_u_wallace_cla16_ha6_and0;
  wire [0:0] h_u_wallace_cla16_fa126_xor1;
  wire [0:0] h_u_wallace_cla16_fa126_or0;
  wire [0:0] h_u_wallace_cla16_fa127_xor1;
  wire [0:0] h_u_wallace_cla16_fa127_or0;
  wire [0:0] h_u_wallace_cla16_fa128_xor1;
  wire [0:0] h_u_wallace_cla16_fa128_or0;
  wire [0:0] h_u_wallace_cla16_and_0_12;
  wire [0:0] h_u_wallace_cla16_fa129_xor1;
  wire [0:0] h_u_wallace_cla16_fa129_or0;
  wire [0:0] h_u_wallace_cla16_and_1_12;
  wire [0:0] h_u_wallace_cla16_and_0_13;
  wire [0:0] h_u_wallace_cla16_fa130_xor1;
  wire [0:0] h_u_wallace_cla16_fa130_or0;
  wire [0:0] h_u_wallace_cla16_and_2_12;
  wire [0:0] h_u_wallace_cla16_and_1_13;
  wire [0:0] h_u_wallace_cla16_fa131_xor1;
  wire [0:0] h_u_wallace_cla16_fa131_or0;
  wire [0:0] h_u_wallace_cla16_and_3_12;
  wire [0:0] h_u_wallace_cla16_and_2_13;
  wire [0:0] h_u_wallace_cla16_fa132_xor1;
  wire [0:0] h_u_wallace_cla16_fa132_or0;
  wire [0:0] h_u_wallace_cla16_and_3_13;
  wire [0:0] h_u_wallace_cla16_and_2_14;
  wire [0:0] h_u_wallace_cla16_fa133_xor1;
  wire [0:0] h_u_wallace_cla16_fa133_or0;
  wire [0:0] h_u_wallace_cla16_and_3_14;
  wire [0:0] h_u_wallace_cla16_and_2_15;
  wire [0:0] h_u_wallace_cla16_fa134_xor1;
  wire [0:0] h_u_wallace_cla16_fa134_or0;
  wire [0:0] h_u_wallace_cla16_and_3_15;
  wire [0:0] h_u_wallace_cla16_fa135_xor1;
  wire [0:0] h_u_wallace_cla16_fa135_or0;
  wire [0:0] h_u_wallace_cla16_fa136_xor1;
  wire [0:0] h_u_wallace_cla16_fa136_or0;
  wire [0:0] h_u_wallace_cla16_fa137_xor1;
  wire [0:0] h_u_wallace_cla16_fa137_or0;
  wire [0:0] h_u_wallace_cla16_fa138_xor1;
  wire [0:0] h_u_wallace_cla16_fa138_or0;
  wire [0:0] h_u_wallace_cla16_fa139_xor1;
  wire [0:0] h_u_wallace_cla16_fa139_or0;
  wire [0:0] h_u_wallace_cla16_ha7_xor0;
  wire [0:0] h_u_wallace_cla16_ha7_and0;
  wire [0:0] h_u_wallace_cla16_fa140_xor1;
  wire [0:0] h_u_wallace_cla16_fa140_or0;
  wire [0:0] h_u_wallace_cla16_fa141_xor1;
  wire [0:0] h_u_wallace_cla16_fa141_or0;
  wire [0:0] h_u_wallace_cla16_fa142_xor1;
  wire [0:0] h_u_wallace_cla16_fa142_or0;
  wire [0:0] h_u_wallace_cla16_fa143_xor1;
  wire [0:0] h_u_wallace_cla16_fa143_or0;
  wire [0:0] h_u_wallace_cla16_and_0_14;
  wire [0:0] h_u_wallace_cla16_fa144_xor1;
  wire [0:0] h_u_wallace_cla16_fa144_or0;
  wire [0:0] h_u_wallace_cla16_and_1_14;
  wire [0:0] h_u_wallace_cla16_and_0_15;
  wire [0:0] h_u_wallace_cla16_fa145_xor1;
  wire [0:0] h_u_wallace_cla16_fa145_or0;
  wire [0:0] h_u_wallace_cla16_and_1_15;
  wire [0:0] h_u_wallace_cla16_fa146_xor1;
  wire [0:0] h_u_wallace_cla16_fa146_or0;
  wire [0:0] h_u_wallace_cla16_fa147_xor1;
  wire [0:0] h_u_wallace_cla16_fa147_or0;
  wire [0:0] h_u_wallace_cla16_fa148_xor1;
  wire [0:0] h_u_wallace_cla16_fa148_or0;
  wire [0:0] h_u_wallace_cla16_fa149_xor1;
  wire [0:0] h_u_wallace_cla16_fa149_or0;
  wire [0:0] h_u_wallace_cla16_fa150_xor1;
  wire [0:0] h_u_wallace_cla16_fa150_or0;
  wire [0:0] h_u_wallace_cla16_fa151_xor1;
  wire [0:0] h_u_wallace_cla16_fa151_or0;
  wire [0:0] h_u_wallace_cla16_ha8_xor0;
  wire [0:0] h_u_wallace_cla16_ha8_and0;
  wire [0:0] h_u_wallace_cla16_fa152_xor1;
  wire [0:0] h_u_wallace_cla16_fa152_or0;
  wire [0:0] h_u_wallace_cla16_fa153_xor1;
  wire [0:0] h_u_wallace_cla16_fa153_or0;
  wire [0:0] h_u_wallace_cla16_fa154_xor1;
  wire [0:0] h_u_wallace_cla16_fa154_or0;
  wire [0:0] h_u_wallace_cla16_fa155_xor1;
  wire [0:0] h_u_wallace_cla16_fa155_or0;
  wire [0:0] h_u_wallace_cla16_fa156_xor1;
  wire [0:0] h_u_wallace_cla16_fa156_or0;
  wire [0:0] h_u_wallace_cla16_fa157_xor1;
  wire [0:0] h_u_wallace_cla16_fa157_or0;
  wire [0:0] h_u_wallace_cla16_fa158_xor1;
  wire [0:0] h_u_wallace_cla16_fa158_or0;
  wire [0:0] h_u_wallace_cla16_fa159_xor1;
  wire [0:0] h_u_wallace_cla16_fa159_or0;
  wire [0:0] h_u_wallace_cla16_fa160_xor1;
  wire [0:0] h_u_wallace_cla16_fa160_or0;
  wire [0:0] h_u_wallace_cla16_fa161_xor1;
  wire [0:0] h_u_wallace_cla16_fa161_or0;
  wire [0:0] h_u_wallace_cla16_ha9_xor0;
  wire [0:0] h_u_wallace_cla16_ha9_and0;
  wire [0:0] h_u_wallace_cla16_fa162_xor1;
  wire [0:0] h_u_wallace_cla16_fa162_or0;
  wire [0:0] h_u_wallace_cla16_fa163_xor1;
  wire [0:0] h_u_wallace_cla16_fa163_or0;
  wire [0:0] h_u_wallace_cla16_fa164_xor1;
  wire [0:0] h_u_wallace_cla16_fa164_or0;
  wire [0:0] h_u_wallace_cla16_fa165_xor1;
  wire [0:0] h_u_wallace_cla16_fa165_or0;
  wire [0:0] h_u_wallace_cla16_fa166_xor1;
  wire [0:0] h_u_wallace_cla16_fa166_or0;
  wire [0:0] h_u_wallace_cla16_fa167_xor1;
  wire [0:0] h_u_wallace_cla16_fa167_or0;
  wire [0:0] h_u_wallace_cla16_fa168_xor1;
  wire [0:0] h_u_wallace_cla16_fa168_or0;
  wire [0:0] h_u_wallace_cla16_fa169_xor1;
  wire [0:0] h_u_wallace_cla16_fa169_or0;
  wire [0:0] h_u_wallace_cla16_ha10_xor0;
  wire [0:0] h_u_wallace_cla16_ha10_and0;
  wire [0:0] h_u_wallace_cla16_fa170_xor1;
  wire [0:0] h_u_wallace_cla16_fa170_or0;
  wire [0:0] h_u_wallace_cla16_fa171_xor1;
  wire [0:0] h_u_wallace_cla16_fa171_or0;
  wire [0:0] h_u_wallace_cla16_fa172_xor1;
  wire [0:0] h_u_wallace_cla16_fa172_or0;
  wire [0:0] h_u_wallace_cla16_fa173_xor1;
  wire [0:0] h_u_wallace_cla16_fa173_or0;
  wire [0:0] h_u_wallace_cla16_fa174_xor1;
  wire [0:0] h_u_wallace_cla16_fa174_or0;
  wire [0:0] h_u_wallace_cla16_fa175_xor1;
  wire [0:0] h_u_wallace_cla16_fa175_or0;
  wire [0:0] h_u_wallace_cla16_ha11_xor0;
  wire [0:0] h_u_wallace_cla16_ha11_and0;
  wire [0:0] h_u_wallace_cla16_fa176_xor1;
  wire [0:0] h_u_wallace_cla16_fa176_or0;
  wire [0:0] h_u_wallace_cla16_fa177_xor1;
  wire [0:0] h_u_wallace_cla16_fa177_or0;
  wire [0:0] h_u_wallace_cla16_fa178_xor1;
  wire [0:0] h_u_wallace_cla16_fa178_or0;
  wire [0:0] h_u_wallace_cla16_fa179_xor1;
  wire [0:0] h_u_wallace_cla16_fa179_or0;
  wire [0:0] h_u_wallace_cla16_ha12_xor0;
  wire [0:0] h_u_wallace_cla16_ha12_and0;
  wire [0:0] h_u_wallace_cla16_fa180_xor1;
  wire [0:0] h_u_wallace_cla16_fa180_or0;
  wire [0:0] h_u_wallace_cla16_fa181_xor1;
  wire [0:0] h_u_wallace_cla16_fa181_or0;
  wire [0:0] h_u_wallace_cla16_ha13_xor0;
  wire [0:0] h_u_wallace_cla16_ha13_and0;
  wire [0:0] h_u_wallace_cla16_ha14_xor0;
  wire [0:0] h_u_wallace_cla16_ha14_and0;
  wire [0:0] h_u_wallace_cla16_fa182_xor1;
  wire [0:0] h_u_wallace_cla16_fa182_or0;
  wire [0:0] h_u_wallace_cla16_fa183_xor1;
  wire [0:0] h_u_wallace_cla16_fa183_or0;
  wire [0:0] h_u_wallace_cla16_fa184_xor1;
  wire [0:0] h_u_wallace_cla16_fa184_or0;
  wire [0:0] h_u_wallace_cla16_fa185_xor1;
  wire [0:0] h_u_wallace_cla16_fa185_or0;
  wire [0:0] h_u_wallace_cla16_fa186_xor1;
  wire [0:0] h_u_wallace_cla16_fa186_or0;
  wire [0:0] h_u_wallace_cla16_fa187_xor1;
  wire [0:0] h_u_wallace_cla16_fa187_or0;
  wire [0:0] h_u_wallace_cla16_fa188_xor1;
  wire [0:0] h_u_wallace_cla16_fa188_or0;
  wire [0:0] h_u_wallace_cla16_fa189_xor1;
  wire [0:0] h_u_wallace_cla16_fa189_or0;
  wire [0:0] h_u_wallace_cla16_fa190_xor1;
  wire [0:0] h_u_wallace_cla16_fa190_or0;
  wire [0:0] h_u_wallace_cla16_fa191_xor1;
  wire [0:0] h_u_wallace_cla16_fa191_or0;
  wire [0:0] h_u_wallace_cla16_fa192_xor1;
  wire [0:0] h_u_wallace_cla16_fa192_or0;
  wire [0:0] h_u_wallace_cla16_and_13_15;
  wire [0:0] h_u_wallace_cla16_fa193_xor1;
  wire [0:0] h_u_wallace_cla16_fa193_or0;
  wire [0:0] h_u_wallace_cla16_and_15_14;
  wire [0:0] h_u_wallace_cla16_fa194_xor1;
  wire [0:0] h_u_wallace_cla16_fa194_or0;
  wire [0:0] h_u_wallace_cla16_and_0_0;
  wire [0:0] h_u_wallace_cla16_and_1_0;
  wire [0:0] h_u_wallace_cla16_and_0_2;
  wire [0:0] h_u_wallace_cla16_and_14_15;
  wire [0:0] h_u_wallace_cla16_and_0_1;
  wire [0:0] h_u_wallace_cla16_and_15_15;
  wire [29:0] h_u_wallace_cla16_u_cla30_a;
  wire [29:0] h_u_wallace_cla16_u_cla30_b;
  wire [30:0] h_u_wallace_cla16_u_cla30_out;

  and_gate and_gate_h_u_wallace_cla16_and_2_0(.a(a[2]), .b(b[0]), .out(h_u_wallace_cla16_and_2_0));
  and_gate and_gate_h_u_wallace_cla16_and_1_1(.a(a[1]), .b(b[1]), .out(h_u_wallace_cla16_and_1_1));
  ha ha_h_u_wallace_cla16_ha0_out(.a(h_u_wallace_cla16_and_2_0[0]), .b(h_u_wallace_cla16_and_1_1[0]), .ha_xor0(h_u_wallace_cla16_ha0_xor0), .ha_and0(h_u_wallace_cla16_ha0_and0));
  and_gate and_gate_h_u_wallace_cla16_and_3_0(.a(a[3]), .b(b[0]), .out(h_u_wallace_cla16_and_3_0));
  and_gate and_gate_h_u_wallace_cla16_and_2_1(.a(a[2]), .b(b[1]), .out(h_u_wallace_cla16_and_2_1));
  fa fa_h_u_wallace_cla16_fa0_out(.a(h_u_wallace_cla16_ha0_and0[0]), .b(h_u_wallace_cla16_and_3_0[0]), .cin(h_u_wallace_cla16_and_2_1[0]), .fa_xor1(h_u_wallace_cla16_fa0_xor1), .fa_or0(h_u_wallace_cla16_fa0_or0));
  and_gate and_gate_h_u_wallace_cla16_and_4_0(.a(a[4]), .b(b[0]), .out(h_u_wallace_cla16_and_4_0));
  and_gate and_gate_h_u_wallace_cla16_and_3_1(.a(a[3]), .b(b[1]), .out(h_u_wallace_cla16_and_3_1));
  fa fa_h_u_wallace_cla16_fa1_out(.a(h_u_wallace_cla16_fa0_or0[0]), .b(h_u_wallace_cla16_and_4_0[0]), .cin(h_u_wallace_cla16_and_3_1[0]), .fa_xor1(h_u_wallace_cla16_fa1_xor1), .fa_or0(h_u_wallace_cla16_fa1_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_0(.a(a[5]), .b(b[0]), .out(h_u_wallace_cla16_and_5_0));
  and_gate and_gate_h_u_wallace_cla16_and_4_1(.a(a[4]), .b(b[1]), .out(h_u_wallace_cla16_and_4_1));
  fa fa_h_u_wallace_cla16_fa2_out(.a(h_u_wallace_cla16_fa1_or0[0]), .b(h_u_wallace_cla16_and_5_0[0]), .cin(h_u_wallace_cla16_and_4_1[0]), .fa_xor1(h_u_wallace_cla16_fa2_xor1), .fa_or0(h_u_wallace_cla16_fa2_or0));
  and_gate and_gate_h_u_wallace_cla16_and_6_0(.a(a[6]), .b(b[0]), .out(h_u_wallace_cla16_and_6_0));
  and_gate and_gate_h_u_wallace_cla16_and_5_1(.a(a[5]), .b(b[1]), .out(h_u_wallace_cla16_and_5_1));
  fa fa_h_u_wallace_cla16_fa3_out(.a(h_u_wallace_cla16_fa2_or0[0]), .b(h_u_wallace_cla16_and_6_0[0]), .cin(h_u_wallace_cla16_and_5_1[0]), .fa_xor1(h_u_wallace_cla16_fa3_xor1), .fa_or0(h_u_wallace_cla16_fa3_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_0(.a(a[7]), .b(b[0]), .out(h_u_wallace_cla16_and_7_0));
  and_gate and_gate_h_u_wallace_cla16_and_6_1(.a(a[6]), .b(b[1]), .out(h_u_wallace_cla16_and_6_1));
  fa fa_h_u_wallace_cla16_fa4_out(.a(h_u_wallace_cla16_fa3_or0[0]), .b(h_u_wallace_cla16_and_7_0[0]), .cin(h_u_wallace_cla16_and_6_1[0]), .fa_xor1(h_u_wallace_cla16_fa4_xor1), .fa_or0(h_u_wallace_cla16_fa4_or0));
  and_gate and_gate_h_u_wallace_cla16_and_8_0(.a(a[8]), .b(b[0]), .out(h_u_wallace_cla16_and_8_0));
  and_gate and_gate_h_u_wallace_cla16_and_7_1(.a(a[7]), .b(b[1]), .out(h_u_wallace_cla16_and_7_1));
  fa fa_h_u_wallace_cla16_fa5_out(.a(h_u_wallace_cla16_fa4_or0[0]), .b(h_u_wallace_cla16_and_8_0[0]), .cin(h_u_wallace_cla16_and_7_1[0]), .fa_xor1(h_u_wallace_cla16_fa5_xor1), .fa_or0(h_u_wallace_cla16_fa5_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_0(.a(a[9]), .b(b[0]), .out(h_u_wallace_cla16_and_9_0));
  and_gate and_gate_h_u_wallace_cla16_and_8_1(.a(a[8]), .b(b[1]), .out(h_u_wallace_cla16_and_8_1));
  fa fa_h_u_wallace_cla16_fa6_out(.a(h_u_wallace_cla16_fa5_or0[0]), .b(h_u_wallace_cla16_and_9_0[0]), .cin(h_u_wallace_cla16_and_8_1[0]), .fa_xor1(h_u_wallace_cla16_fa6_xor1), .fa_or0(h_u_wallace_cla16_fa6_or0));
  and_gate and_gate_h_u_wallace_cla16_and_10_0(.a(a[10]), .b(b[0]), .out(h_u_wallace_cla16_and_10_0));
  and_gate and_gate_h_u_wallace_cla16_and_9_1(.a(a[9]), .b(b[1]), .out(h_u_wallace_cla16_and_9_1));
  fa fa_h_u_wallace_cla16_fa7_out(.a(h_u_wallace_cla16_fa6_or0[0]), .b(h_u_wallace_cla16_and_10_0[0]), .cin(h_u_wallace_cla16_and_9_1[0]), .fa_xor1(h_u_wallace_cla16_fa7_xor1), .fa_or0(h_u_wallace_cla16_fa7_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_0(.a(a[11]), .b(b[0]), .out(h_u_wallace_cla16_and_11_0));
  and_gate and_gate_h_u_wallace_cla16_and_10_1(.a(a[10]), .b(b[1]), .out(h_u_wallace_cla16_and_10_1));
  fa fa_h_u_wallace_cla16_fa8_out(.a(h_u_wallace_cla16_fa7_or0[0]), .b(h_u_wallace_cla16_and_11_0[0]), .cin(h_u_wallace_cla16_and_10_1[0]), .fa_xor1(h_u_wallace_cla16_fa8_xor1), .fa_or0(h_u_wallace_cla16_fa8_or0));
  and_gate and_gate_h_u_wallace_cla16_and_12_0(.a(a[12]), .b(b[0]), .out(h_u_wallace_cla16_and_12_0));
  and_gate and_gate_h_u_wallace_cla16_and_11_1(.a(a[11]), .b(b[1]), .out(h_u_wallace_cla16_and_11_1));
  fa fa_h_u_wallace_cla16_fa9_out(.a(h_u_wallace_cla16_fa8_or0[0]), .b(h_u_wallace_cla16_and_12_0[0]), .cin(h_u_wallace_cla16_and_11_1[0]), .fa_xor1(h_u_wallace_cla16_fa9_xor1), .fa_or0(h_u_wallace_cla16_fa9_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_0(.a(a[13]), .b(b[0]), .out(h_u_wallace_cla16_and_13_0));
  and_gate and_gate_h_u_wallace_cla16_and_12_1(.a(a[12]), .b(b[1]), .out(h_u_wallace_cla16_and_12_1));
  fa fa_h_u_wallace_cla16_fa10_out(.a(h_u_wallace_cla16_fa9_or0[0]), .b(h_u_wallace_cla16_and_13_0[0]), .cin(h_u_wallace_cla16_and_12_1[0]), .fa_xor1(h_u_wallace_cla16_fa10_xor1), .fa_or0(h_u_wallace_cla16_fa10_or0));
  and_gate and_gate_h_u_wallace_cla16_and_14_0(.a(a[14]), .b(b[0]), .out(h_u_wallace_cla16_and_14_0));
  and_gate and_gate_h_u_wallace_cla16_and_13_1(.a(a[13]), .b(b[1]), .out(h_u_wallace_cla16_and_13_1));
  fa fa_h_u_wallace_cla16_fa11_out(.a(h_u_wallace_cla16_fa10_or0[0]), .b(h_u_wallace_cla16_and_14_0[0]), .cin(h_u_wallace_cla16_and_13_1[0]), .fa_xor1(h_u_wallace_cla16_fa11_xor1), .fa_or0(h_u_wallace_cla16_fa11_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_0(.a(a[15]), .b(b[0]), .out(h_u_wallace_cla16_and_15_0));
  and_gate and_gate_h_u_wallace_cla16_and_14_1(.a(a[14]), .b(b[1]), .out(h_u_wallace_cla16_and_14_1));
  fa fa_h_u_wallace_cla16_fa12_out(.a(h_u_wallace_cla16_fa11_or0[0]), .b(h_u_wallace_cla16_and_15_0[0]), .cin(h_u_wallace_cla16_and_14_1[0]), .fa_xor1(h_u_wallace_cla16_fa12_xor1), .fa_or0(h_u_wallace_cla16_fa12_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_1(.a(a[15]), .b(b[1]), .out(h_u_wallace_cla16_and_15_1));
  and_gate and_gate_h_u_wallace_cla16_and_14_2(.a(a[14]), .b(b[2]), .out(h_u_wallace_cla16_and_14_2));
  fa fa_h_u_wallace_cla16_fa13_out(.a(h_u_wallace_cla16_fa12_or0[0]), .b(h_u_wallace_cla16_and_15_1[0]), .cin(h_u_wallace_cla16_and_14_2[0]), .fa_xor1(h_u_wallace_cla16_fa13_xor1), .fa_or0(h_u_wallace_cla16_fa13_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_2(.a(a[15]), .b(b[2]), .out(h_u_wallace_cla16_and_15_2));
  and_gate and_gate_h_u_wallace_cla16_and_14_3(.a(a[14]), .b(b[3]), .out(h_u_wallace_cla16_and_14_3));
  fa fa_h_u_wallace_cla16_fa14_out(.a(h_u_wallace_cla16_fa13_or0[0]), .b(h_u_wallace_cla16_and_15_2[0]), .cin(h_u_wallace_cla16_and_14_3[0]), .fa_xor1(h_u_wallace_cla16_fa14_xor1), .fa_or0(h_u_wallace_cla16_fa14_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_3(.a(a[15]), .b(b[3]), .out(h_u_wallace_cla16_and_15_3));
  and_gate and_gate_h_u_wallace_cla16_and_14_4(.a(a[14]), .b(b[4]), .out(h_u_wallace_cla16_and_14_4));
  fa fa_h_u_wallace_cla16_fa15_out(.a(h_u_wallace_cla16_fa14_or0[0]), .b(h_u_wallace_cla16_and_15_3[0]), .cin(h_u_wallace_cla16_and_14_4[0]), .fa_xor1(h_u_wallace_cla16_fa15_xor1), .fa_or0(h_u_wallace_cla16_fa15_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_4(.a(a[15]), .b(b[4]), .out(h_u_wallace_cla16_and_15_4));
  and_gate and_gate_h_u_wallace_cla16_and_14_5(.a(a[14]), .b(b[5]), .out(h_u_wallace_cla16_and_14_5));
  fa fa_h_u_wallace_cla16_fa16_out(.a(h_u_wallace_cla16_fa15_or0[0]), .b(h_u_wallace_cla16_and_15_4[0]), .cin(h_u_wallace_cla16_and_14_5[0]), .fa_xor1(h_u_wallace_cla16_fa16_xor1), .fa_or0(h_u_wallace_cla16_fa16_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_5(.a(a[15]), .b(b[5]), .out(h_u_wallace_cla16_and_15_5));
  and_gate and_gate_h_u_wallace_cla16_and_14_6(.a(a[14]), .b(b[6]), .out(h_u_wallace_cla16_and_14_6));
  fa fa_h_u_wallace_cla16_fa17_out(.a(h_u_wallace_cla16_fa16_or0[0]), .b(h_u_wallace_cla16_and_15_5[0]), .cin(h_u_wallace_cla16_and_14_6[0]), .fa_xor1(h_u_wallace_cla16_fa17_xor1), .fa_or0(h_u_wallace_cla16_fa17_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_6(.a(a[15]), .b(b[6]), .out(h_u_wallace_cla16_and_15_6));
  and_gate and_gate_h_u_wallace_cla16_and_14_7(.a(a[14]), .b(b[7]), .out(h_u_wallace_cla16_and_14_7));
  fa fa_h_u_wallace_cla16_fa18_out(.a(h_u_wallace_cla16_fa17_or0[0]), .b(h_u_wallace_cla16_and_15_6[0]), .cin(h_u_wallace_cla16_and_14_7[0]), .fa_xor1(h_u_wallace_cla16_fa18_xor1), .fa_or0(h_u_wallace_cla16_fa18_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_7(.a(a[15]), .b(b[7]), .out(h_u_wallace_cla16_and_15_7));
  and_gate and_gate_h_u_wallace_cla16_and_14_8(.a(a[14]), .b(b[8]), .out(h_u_wallace_cla16_and_14_8));
  fa fa_h_u_wallace_cla16_fa19_out(.a(h_u_wallace_cla16_fa18_or0[0]), .b(h_u_wallace_cla16_and_15_7[0]), .cin(h_u_wallace_cla16_and_14_8[0]), .fa_xor1(h_u_wallace_cla16_fa19_xor1), .fa_or0(h_u_wallace_cla16_fa19_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_8(.a(a[15]), .b(b[8]), .out(h_u_wallace_cla16_and_15_8));
  and_gate and_gate_h_u_wallace_cla16_and_14_9(.a(a[14]), .b(b[9]), .out(h_u_wallace_cla16_and_14_9));
  fa fa_h_u_wallace_cla16_fa20_out(.a(h_u_wallace_cla16_fa19_or0[0]), .b(h_u_wallace_cla16_and_15_8[0]), .cin(h_u_wallace_cla16_and_14_9[0]), .fa_xor1(h_u_wallace_cla16_fa20_xor1), .fa_or0(h_u_wallace_cla16_fa20_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_9(.a(a[15]), .b(b[9]), .out(h_u_wallace_cla16_and_15_9));
  and_gate and_gate_h_u_wallace_cla16_and_14_10(.a(a[14]), .b(b[10]), .out(h_u_wallace_cla16_and_14_10));
  fa fa_h_u_wallace_cla16_fa21_out(.a(h_u_wallace_cla16_fa20_or0[0]), .b(h_u_wallace_cla16_and_15_9[0]), .cin(h_u_wallace_cla16_and_14_10[0]), .fa_xor1(h_u_wallace_cla16_fa21_xor1), .fa_or0(h_u_wallace_cla16_fa21_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_10(.a(a[15]), .b(b[10]), .out(h_u_wallace_cla16_and_15_10));
  and_gate and_gate_h_u_wallace_cla16_and_14_11(.a(a[14]), .b(b[11]), .out(h_u_wallace_cla16_and_14_11));
  fa fa_h_u_wallace_cla16_fa22_out(.a(h_u_wallace_cla16_fa21_or0[0]), .b(h_u_wallace_cla16_and_15_10[0]), .cin(h_u_wallace_cla16_and_14_11[0]), .fa_xor1(h_u_wallace_cla16_fa22_xor1), .fa_or0(h_u_wallace_cla16_fa22_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_11(.a(a[15]), .b(b[11]), .out(h_u_wallace_cla16_and_15_11));
  and_gate and_gate_h_u_wallace_cla16_and_14_12(.a(a[14]), .b(b[12]), .out(h_u_wallace_cla16_and_14_12));
  fa fa_h_u_wallace_cla16_fa23_out(.a(h_u_wallace_cla16_fa22_or0[0]), .b(h_u_wallace_cla16_and_15_11[0]), .cin(h_u_wallace_cla16_and_14_12[0]), .fa_xor1(h_u_wallace_cla16_fa23_xor1), .fa_or0(h_u_wallace_cla16_fa23_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_12(.a(a[15]), .b(b[12]), .out(h_u_wallace_cla16_and_15_12));
  and_gate and_gate_h_u_wallace_cla16_and_14_13(.a(a[14]), .b(b[13]), .out(h_u_wallace_cla16_and_14_13));
  fa fa_h_u_wallace_cla16_fa24_out(.a(h_u_wallace_cla16_fa23_or0[0]), .b(h_u_wallace_cla16_and_15_12[0]), .cin(h_u_wallace_cla16_and_14_13[0]), .fa_xor1(h_u_wallace_cla16_fa24_xor1), .fa_or0(h_u_wallace_cla16_fa24_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_13(.a(a[15]), .b(b[13]), .out(h_u_wallace_cla16_and_15_13));
  and_gate and_gate_h_u_wallace_cla16_and_14_14(.a(a[14]), .b(b[14]), .out(h_u_wallace_cla16_and_14_14));
  fa fa_h_u_wallace_cla16_fa25_out(.a(h_u_wallace_cla16_fa24_or0[0]), .b(h_u_wallace_cla16_and_15_13[0]), .cin(h_u_wallace_cla16_and_14_14[0]), .fa_xor1(h_u_wallace_cla16_fa25_xor1), .fa_or0(h_u_wallace_cla16_fa25_or0));
  and_gate and_gate_h_u_wallace_cla16_and_1_2(.a(a[1]), .b(b[2]), .out(h_u_wallace_cla16_and_1_2));
  and_gate and_gate_h_u_wallace_cla16_and_0_3(.a(a[0]), .b(b[3]), .out(h_u_wallace_cla16_and_0_3));
  ha ha_h_u_wallace_cla16_ha1_out(.a(h_u_wallace_cla16_and_1_2[0]), .b(h_u_wallace_cla16_and_0_3[0]), .ha_xor0(h_u_wallace_cla16_ha1_xor0), .ha_and0(h_u_wallace_cla16_ha1_and0));
  and_gate and_gate_h_u_wallace_cla16_and_2_2(.a(a[2]), .b(b[2]), .out(h_u_wallace_cla16_and_2_2));
  and_gate and_gate_h_u_wallace_cla16_and_1_3(.a(a[1]), .b(b[3]), .out(h_u_wallace_cla16_and_1_3));
  fa fa_h_u_wallace_cla16_fa26_out(.a(h_u_wallace_cla16_ha1_and0[0]), .b(h_u_wallace_cla16_and_2_2[0]), .cin(h_u_wallace_cla16_and_1_3[0]), .fa_xor1(h_u_wallace_cla16_fa26_xor1), .fa_or0(h_u_wallace_cla16_fa26_or0));
  and_gate and_gate_h_u_wallace_cla16_and_3_2(.a(a[3]), .b(b[2]), .out(h_u_wallace_cla16_and_3_2));
  and_gate and_gate_h_u_wallace_cla16_and_2_3(.a(a[2]), .b(b[3]), .out(h_u_wallace_cla16_and_2_3));
  fa fa_h_u_wallace_cla16_fa27_out(.a(h_u_wallace_cla16_fa26_or0[0]), .b(h_u_wallace_cla16_and_3_2[0]), .cin(h_u_wallace_cla16_and_2_3[0]), .fa_xor1(h_u_wallace_cla16_fa27_xor1), .fa_or0(h_u_wallace_cla16_fa27_or0));
  and_gate and_gate_h_u_wallace_cla16_and_4_2(.a(a[4]), .b(b[2]), .out(h_u_wallace_cla16_and_4_2));
  and_gate and_gate_h_u_wallace_cla16_and_3_3(.a(a[3]), .b(b[3]), .out(h_u_wallace_cla16_and_3_3));
  fa fa_h_u_wallace_cla16_fa28_out(.a(h_u_wallace_cla16_fa27_or0[0]), .b(h_u_wallace_cla16_and_4_2[0]), .cin(h_u_wallace_cla16_and_3_3[0]), .fa_xor1(h_u_wallace_cla16_fa28_xor1), .fa_or0(h_u_wallace_cla16_fa28_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_2(.a(a[5]), .b(b[2]), .out(h_u_wallace_cla16_and_5_2));
  and_gate and_gate_h_u_wallace_cla16_and_4_3(.a(a[4]), .b(b[3]), .out(h_u_wallace_cla16_and_4_3));
  fa fa_h_u_wallace_cla16_fa29_out(.a(h_u_wallace_cla16_fa28_or0[0]), .b(h_u_wallace_cla16_and_5_2[0]), .cin(h_u_wallace_cla16_and_4_3[0]), .fa_xor1(h_u_wallace_cla16_fa29_xor1), .fa_or0(h_u_wallace_cla16_fa29_or0));
  and_gate and_gate_h_u_wallace_cla16_and_6_2(.a(a[6]), .b(b[2]), .out(h_u_wallace_cla16_and_6_2));
  and_gate and_gate_h_u_wallace_cla16_and_5_3(.a(a[5]), .b(b[3]), .out(h_u_wallace_cla16_and_5_3));
  fa fa_h_u_wallace_cla16_fa30_out(.a(h_u_wallace_cla16_fa29_or0[0]), .b(h_u_wallace_cla16_and_6_2[0]), .cin(h_u_wallace_cla16_and_5_3[0]), .fa_xor1(h_u_wallace_cla16_fa30_xor1), .fa_or0(h_u_wallace_cla16_fa30_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_2(.a(a[7]), .b(b[2]), .out(h_u_wallace_cla16_and_7_2));
  and_gate and_gate_h_u_wallace_cla16_and_6_3(.a(a[6]), .b(b[3]), .out(h_u_wallace_cla16_and_6_3));
  fa fa_h_u_wallace_cla16_fa31_out(.a(h_u_wallace_cla16_fa30_or0[0]), .b(h_u_wallace_cla16_and_7_2[0]), .cin(h_u_wallace_cla16_and_6_3[0]), .fa_xor1(h_u_wallace_cla16_fa31_xor1), .fa_or0(h_u_wallace_cla16_fa31_or0));
  and_gate and_gate_h_u_wallace_cla16_and_8_2(.a(a[8]), .b(b[2]), .out(h_u_wallace_cla16_and_8_2));
  and_gate and_gate_h_u_wallace_cla16_and_7_3(.a(a[7]), .b(b[3]), .out(h_u_wallace_cla16_and_7_3));
  fa fa_h_u_wallace_cla16_fa32_out(.a(h_u_wallace_cla16_fa31_or0[0]), .b(h_u_wallace_cla16_and_8_2[0]), .cin(h_u_wallace_cla16_and_7_3[0]), .fa_xor1(h_u_wallace_cla16_fa32_xor1), .fa_or0(h_u_wallace_cla16_fa32_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_2(.a(a[9]), .b(b[2]), .out(h_u_wallace_cla16_and_9_2));
  and_gate and_gate_h_u_wallace_cla16_and_8_3(.a(a[8]), .b(b[3]), .out(h_u_wallace_cla16_and_8_3));
  fa fa_h_u_wallace_cla16_fa33_out(.a(h_u_wallace_cla16_fa32_or0[0]), .b(h_u_wallace_cla16_and_9_2[0]), .cin(h_u_wallace_cla16_and_8_3[0]), .fa_xor1(h_u_wallace_cla16_fa33_xor1), .fa_or0(h_u_wallace_cla16_fa33_or0));
  and_gate and_gate_h_u_wallace_cla16_and_10_2(.a(a[10]), .b(b[2]), .out(h_u_wallace_cla16_and_10_2));
  and_gate and_gate_h_u_wallace_cla16_and_9_3(.a(a[9]), .b(b[3]), .out(h_u_wallace_cla16_and_9_3));
  fa fa_h_u_wallace_cla16_fa34_out(.a(h_u_wallace_cla16_fa33_or0[0]), .b(h_u_wallace_cla16_and_10_2[0]), .cin(h_u_wallace_cla16_and_9_3[0]), .fa_xor1(h_u_wallace_cla16_fa34_xor1), .fa_or0(h_u_wallace_cla16_fa34_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_2(.a(a[11]), .b(b[2]), .out(h_u_wallace_cla16_and_11_2));
  and_gate and_gate_h_u_wallace_cla16_and_10_3(.a(a[10]), .b(b[3]), .out(h_u_wallace_cla16_and_10_3));
  fa fa_h_u_wallace_cla16_fa35_out(.a(h_u_wallace_cla16_fa34_or0[0]), .b(h_u_wallace_cla16_and_11_2[0]), .cin(h_u_wallace_cla16_and_10_3[0]), .fa_xor1(h_u_wallace_cla16_fa35_xor1), .fa_or0(h_u_wallace_cla16_fa35_or0));
  and_gate and_gate_h_u_wallace_cla16_and_12_2(.a(a[12]), .b(b[2]), .out(h_u_wallace_cla16_and_12_2));
  and_gate and_gate_h_u_wallace_cla16_and_11_3(.a(a[11]), .b(b[3]), .out(h_u_wallace_cla16_and_11_3));
  fa fa_h_u_wallace_cla16_fa36_out(.a(h_u_wallace_cla16_fa35_or0[0]), .b(h_u_wallace_cla16_and_12_2[0]), .cin(h_u_wallace_cla16_and_11_3[0]), .fa_xor1(h_u_wallace_cla16_fa36_xor1), .fa_or0(h_u_wallace_cla16_fa36_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_2(.a(a[13]), .b(b[2]), .out(h_u_wallace_cla16_and_13_2));
  and_gate and_gate_h_u_wallace_cla16_and_12_3(.a(a[12]), .b(b[3]), .out(h_u_wallace_cla16_and_12_3));
  fa fa_h_u_wallace_cla16_fa37_out(.a(h_u_wallace_cla16_fa36_or0[0]), .b(h_u_wallace_cla16_and_13_2[0]), .cin(h_u_wallace_cla16_and_12_3[0]), .fa_xor1(h_u_wallace_cla16_fa37_xor1), .fa_or0(h_u_wallace_cla16_fa37_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_3(.a(a[13]), .b(b[3]), .out(h_u_wallace_cla16_and_13_3));
  and_gate and_gate_h_u_wallace_cla16_and_12_4(.a(a[12]), .b(b[4]), .out(h_u_wallace_cla16_and_12_4));
  fa fa_h_u_wallace_cla16_fa38_out(.a(h_u_wallace_cla16_fa37_or0[0]), .b(h_u_wallace_cla16_and_13_3[0]), .cin(h_u_wallace_cla16_and_12_4[0]), .fa_xor1(h_u_wallace_cla16_fa38_xor1), .fa_or0(h_u_wallace_cla16_fa38_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_4(.a(a[13]), .b(b[4]), .out(h_u_wallace_cla16_and_13_4));
  and_gate and_gate_h_u_wallace_cla16_and_12_5(.a(a[12]), .b(b[5]), .out(h_u_wallace_cla16_and_12_5));
  fa fa_h_u_wallace_cla16_fa39_out(.a(h_u_wallace_cla16_fa38_or0[0]), .b(h_u_wallace_cla16_and_13_4[0]), .cin(h_u_wallace_cla16_and_12_5[0]), .fa_xor1(h_u_wallace_cla16_fa39_xor1), .fa_or0(h_u_wallace_cla16_fa39_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_5(.a(a[13]), .b(b[5]), .out(h_u_wallace_cla16_and_13_5));
  and_gate and_gate_h_u_wallace_cla16_and_12_6(.a(a[12]), .b(b[6]), .out(h_u_wallace_cla16_and_12_6));
  fa fa_h_u_wallace_cla16_fa40_out(.a(h_u_wallace_cla16_fa39_or0[0]), .b(h_u_wallace_cla16_and_13_5[0]), .cin(h_u_wallace_cla16_and_12_6[0]), .fa_xor1(h_u_wallace_cla16_fa40_xor1), .fa_or0(h_u_wallace_cla16_fa40_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_6(.a(a[13]), .b(b[6]), .out(h_u_wallace_cla16_and_13_6));
  and_gate and_gate_h_u_wallace_cla16_and_12_7(.a(a[12]), .b(b[7]), .out(h_u_wallace_cla16_and_12_7));
  fa fa_h_u_wallace_cla16_fa41_out(.a(h_u_wallace_cla16_fa40_or0[0]), .b(h_u_wallace_cla16_and_13_6[0]), .cin(h_u_wallace_cla16_and_12_7[0]), .fa_xor1(h_u_wallace_cla16_fa41_xor1), .fa_or0(h_u_wallace_cla16_fa41_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_7(.a(a[13]), .b(b[7]), .out(h_u_wallace_cla16_and_13_7));
  and_gate and_gate_h_u_wallace_cla16_and_12_8(.a(a[12]), .b(b[8]), .out(h_u_wallace_cla16_and_12_8));
  fa fa_h_u_wallace_cla16_fa42_out(.a(h_u_wallace_cla16_fa41_or0[0]), .b(h_u_wallace_cla16_and_13_7[0]), .cin(h_u_wallace_cla16_and_12_8[0]), .fa_xor1(h_u_wallace_cla16_fa42_xor1), .fa_or0(h_u_wallace_cla16_fa42_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_8(.a(a[13]), .b(b[8]), .out(h_u_wallace_cla16_and_13_8));
  and_gate and_gate_h_u_wallace_cla16_and_12_9(.a(a[12]), .b(b[9]), .out(h_u_wallace_cla16_and_12_9));
  fa fa_h_u_wallace_cla16_fa43_out(.a(h_u_wallace_cla16_fa42_or0[0]), .b(h_u_wallace_cla16_and_13_8[0]), .cin(h_u_wallace_cla16_and_12_9[0]), .fa_xor1(h_u_wallace_cla16_fa43_xor1), .fa_or0(h_u_wallace_cla16_fa43_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_9(.a(a[13]), .b(b[9]), .out(h_u_wallace_cla16_and_13_9));
  and_gate and_gate_h_u_wallace_cla16_and_12_10(.a(a[12]), .b(b[10]), .out(h_u_wallace_cla16_and_12_10));
  fa fa_h_u_wallace_cla16_fa44_out(.a(h_u_wallace_cla16_fa43_or0[0]), .b(h_u_wallace_cla16_and_13_9[0]), .cin(h_u_wallace_cla16_and_12_10[0]), .fa_xor1(h_u_wallace_cla16_fa44_xor1), .fa_or0(h_u_wallace_cla16_fa44_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_10(.a(a[13]), .b(b[10]), .out(h_u_wallace_cla16_and_13_10));
  and_gate and_gate_h_u_wallace_cla16_and_12_11(.a(a[12]), .b(b[11]), .out(h_u_wallace_cla16_and_12_11));
  fa fa_h_u_wallace_cla16_fa45_out(.a(h_u_wallace_cla16_fa44_or0[0]), .b(h_u_wallace_cla16_and_13_10[0]), .cin(h_u_wallace_cla16_and_12_11[0]), .fa_xor1(h_u_wallace_cla16_fa45_xor1), .fa_or0(h_u_wallace_cla16_fa45_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_11(.a(a[13]), .b(b[11]), .out(h_u_wallace_cla16_and_13_11));
  and_gate and_gate_h_u_wallace_cla16_and_12_12(.a(a[12]), .b(b[12]), .out(h_u_wallace_cla16_and_12_12));
  fa fa_h_u_wallace_cla16_fa46_out(.a(h_u_wallace_cla16_fa45_or0[0]), .b(h_u_wallace_cla16_and_13_11[0]), .cin(h_u_wallace_cla16_and_12_12[0]), .fa_xor1(h_u_wallace_cla16_fa46_xor1), .fa_or0(h_u_wallace_cla16_fa46_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_12(.a(a[13]), .b(b[12]), .out(h_u_wallace_cla16_and_13_12));
  and_gate and_gate_h_u_wallace_cla16_and_12_13(.a(a[12]), .b(b[13]), .out(h_u_wallace_cla16_and_12_13));
  fa fa_h_u_wallace_cla16_fa47_out(.a(h_u_wallace_cla16_fa46_or0[0]), .b(h_u_wallace_cla16_and_13_12[0]), .cin(h_u_wallace_cla16_and_12_13[0]), .fa_xor1(h_u_wallace_cla16_fa47_xor1), .fa_or0(h_u_wallace_cla16_fa47_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_13(.a(a[13]), .b(b[13]), .out(h_u_wallace_cla16_and_13_13));
  and_gate and_gate_h_u_wallace_cla16_and_12_14(.a(a[12]), .b(b[14]), .out(h_u_wallace_cla16_and_12_14));
  fa fa_h_u_wallace_cla16_fa48_out(.a(h_u_wallace_cla16_fa47_or0[0]), .b(h_u_wallace_cla16_and_13_13[0]), .cin(h_u_wallace_cla16_and_12_14[0]), .fa_xor1(h_u_wallace_cla16_fa48_xor1), .fa_or0(h_u_wallace_cla16_fa48_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_14(.a(a[13]), .b(b[14]), .out(h_u_wallace_cla16_and_13_14));
  and_gate and_gate_h_u_wallace_cla16_and_12_15(.a(a[12]), .b(b[15]), .out(h_u_wallace_cla16_and_12_15));
  fa fa_h_u_wallace_cla16_fa49_out(.a(h_u_wallace_cla16_fa48_or0[0]), .b(h_u_wallace_cla16_and_13_14[0]), .cin(h_u_wallace_cla16_and_12_15[0]), .fa_xor1(h_u_wallace_cla16_fa49_xor1), .fa_or0(h_u_wallace_cla16_fa49_or0));
  and_gate and_gate_h_u_wallace_cla16_and_0_4(.a(a[0]), .b(b[4]), .out(h_u_wallace_cla16_and_0_4));
  ha ha_h_u_wallace_cla16_ha2_out(.a(h_u_wallace_cla16_and_0_4[0]), .b(h_u_wallace_cla16_fa1_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha2_xor0), .ha_and0(h_u_wallace_cla16_ha2_and0));
  and_gate and_gate_h_u_wallace_cla16_and_1_4(.a(a[1]), .b(b[4]), .out(h_u_wallace_cla16_and_1_4));
  and_gate and_gate_h_u_wallace_cla16_and_0_5(.a(a[0]), .b(b[5]), .out(h_u_wallace_cla16_and_0_5));
  fa fa_h_u_wallace_cla16_fa50_out(.a(h_u_wallace_cla16_ha2_and0[0]), .b(h_u_wallace_cla16_and_1_4[0]), .cin(h_u_wallace_cla16_and_0_5[0]), .fa_xor1(h_u_wallace_cla16_fa50_xor1), .fa_or0(h_u_wallace_cla16_fa50_or0));
  and_gate and_gate_h_u_wallace_cla16_and_2_4(.a(a[2]), .b(b[4]), .out(h_u_wallace_cla16_and_2_4));
  and_gate and_gate_h_u_wallace_cla16_and_1_5(.a(a[1]), .b(b[5]), .out(h_u_wallace_cla16_and_1_5));
  fa fa_h_u_wallace_cla16_fa51_out(.a(h_u_wallace_cla16_fa50_or0[0]), .b(h_u_wallace_cla16_and_2_4[0]), .cin(h_u_wallace_cla16_and_1_5[0]), .fa_xor1(h_u_wallace_cla16_fa51_xor1), .fa_or0(h_u_wallace_cla16_fa51_or0));
  and_gate and_gate_h_u_wallace_cla16_and_3_4(.a(a[3]), .b(b[4]), .out(h_u_wallace_cla16_and_3_4));
  and_gate and_gate_h_u_wallace_cla16_and_2_5(.a(a[2]), .b(b[5]), .out(h_u_wallace_cla16_and_2_5));
  fa fa_h_u_wallace_cla16_fa52_out(.a(h_u_wallace_cla16_fa51_or0[0]), .b(h_u_wallace_cla16_and_3_4[0]), .cin(h_u_wallace_cla16_and_2_5[0]), .fa_xor1(h_u_wallace_cla16_fa52_xor1), .fa_or0(h_u_wallace_cla16_fa52_or0));
  and_gate and_gate_h_u_wallace_cla16_and_4_4(.a(a[4]), .b(b[4]), .out(h_u_wallace_cla16_and_4_4));
  and_gate and_gate_h_u_wallace_cla16_and_3_5(.a(a[3]), .b(b[5]), .out(h_u_wallace_cla16_and_3_5));
  fa fa_h_u_wallace_cla16_fa53_out(.a(h_u_wallace_cla16_fa52_or0[0]), .b(h_u_wallace_cla16_and_4_4[0]), .cin(h_u_wallace_cla16_and_3_5[0]), .fa_xor1(h_u_wallace_cla16_fa53_xor1), .fa_or0(h_u_wallace_cla16_fa53_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_4(.a(a[5]), .b(b[4]), .out(h_u_wallace_cla16_and_5_4));
  and_gate and_gate_h_u_wallace_cla16_and_4_5(.a(a[4]), .b(b[5]), .out(h_u_wallace_cla16_and_4_5));
  fa fa_h_u_wallace_cla16_fa54_out(.a(h_u_wallace_cla16_fa53_or0[0]), .b(h_u_wallace_cla16_and_5_4[0]), .cin(h_u_wallace_cla16_and_4_5[0]), .fa_xor1(h_u_wallace_cla16_fa54_xor1), .fa_or0(h_u_wallace_cla16_fa54_or0));
  and_gate and_gate_h_u_wallace_cla16_and_6_4(.a(a[6]), .b(b[4]), .out(h_u_wallace_cla16_and_6_4));
  and_gate and_gate_h_u_wallace_cla16_and_5_5(.a(a[5]), .b(b[5]), .out(h_u_wallace_cla16_and_5_5));
  fa fa_h_u_wallace_cla16_fa55_out(.a(h_u_wallace_cla16_fa54_or0[0]), .b(h_u_wallace_cla16_and_6_4[0]), .cin(h_u_wallace_cla16_and_5_5[0]), .fa_xor1(h_u_wallace_cla16_fa55_xor1), .fa_or0(h_u_wallace_cla16_fa55_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_4(.a(a[7]), .b(b[4]), .out(h_u_wallace_cla16_and_7_4));
  and_gate and_gate_h_u_wallace_cla16_and_6_5(.a(a[6]), .b(b[5]), .out(h_u_wallace_cla16_and_6_5));
  fa fa_h_u_wallace_cla16_fa56_out(.a(h_u_wallace_cla16_fa55_or0[0]), .b(h_u_wallace_cla16_and_7_4[0]), .cin(h_u_wallace_cla16_and_6_5[0]), .fa_xor1(h_u_wallace_cla16_fa56_xor1), .fa_or0(h_u_wallace_cla16_fa56_or0));
  and_gate and_gate_h_u_wallace_cla16_and_8_4(.a(a[8]), .b(b[4]), .out(h_u_wallace_cla16_and_8_4));
  and_gate and_gate_h_u_wallace_cla16_and_7_5(.a(a[7]), .b(b[5]), .out(h_u_wallace_cla16_and_7_5));
  fa fa_h_u_wallace_cla16_fa57_out(.a(h_u_wallace_cla16_fa56_or0[0]), .b(h_u_wallace_cla16_and_8_4[0]), .cin(h_u_wallace_cla16_and_7_5[0]), .fa_xor1(h_u_wallace_cla16_fa57_xor1), .fa_or0(h_u_wallace_cla16_fa57_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_4(.a(a[9]), .b(b[4]), .out(h_u_wallace_cla16_and_9_4));
  and_gate and_gate_h_u_wallace_cla16_and_8_5(.a(a[8]), .b(b[5]), .out(h_u_wallace_cla16_and_8_5));
  fa fa_h_u_wallace_cla16_fa58_out(.a(h_u_wallace_cla16_fa57_or0[0]), .b(h_u_wallace_cla16_and_9_4[0]), .cin(h_u_wallace_cla16_and_8_5[0]), .fa_xor1(h_u_wallace_cla16_fa58_xor1), .fa_or0(h_u_wallace_cla16_fa58_or0));
  and_gate and_gate_h_u_wallace_cla16_and_10_4(.a(a[10]), .b(b[4]), .out(h_u_wallace_cla16_and_10_4));
  and_gate and_gate_h_u_wallace_cla16_and_9_5(.a(a[9]), .b(b[5]), .out(h_u_wallace_cla16_and_9_5));
  fa fa_h_u_wallace_cla16_fa59_out(.a(h_u_wallace_cla16_fa58_or0[0]), .b(h_u_wallace_cla16_and_10_4[0]), .cin(h_u_wallace_cla16_and_9_5[0]), .fa_xor1(h_u_wallace_cla16_fa59_xor1), .fa_or0(h_u_wallace_cla16_fa59_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_4(.a(a[11]), .b(b[4]), .out(h_u_wallace_cla16_and_11_4));
  and_gate and_gate_h_u_wallace_cla16_and_10_5(.a(a[10]), .b(b[5]), .out(h_u_wallace_cla16_and_10_5));
  fa fa_h_u_wallace_cla16_fa60_out(.a(h_u_wallace_cla16_fa59_or0[0]), .b(h_u_wallace_cla16_and_11_4[0]), .cin(h_u_wallace_cla16_and_10_5[0]), .fa_xor1(h_u_wallace_cla16_fa60_xor1), .fa_or0(h_u_wallace_cla16_fa60_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_5(.a(a[11]), .b(b[5]), .out(h_u_wallace_cla16_and_11_5));
  and_gate and_gate_h_u_wallace_cla16_and_10_6(.a(a[10]), .b(b[6]), .out(h_u_wallace_cla16_and_10_6));
  fa fa_h_u_wallace_cla16_fa61_out(.a(h_u_wallace_cla16_fa60_or0[0]), .b(h_u_wallace_cla16_and_11_5[0]), .cin(h_u_wallace_cla16_and_10_6[0]), .fa_xor1(h_u_wallace_cla16_fa61_xor1), .fa_or0(h_u_wallace_cla16_fa61_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_6(.a(a[11]), .b(b[6]), .out(h_u_wallace_cla16_and_11_6));
  and_gate and_gate_h_u_wallace_cla16_and_10_7(.a(a[10]), .b(b[7]), .out(h_u_wallace_cla16_and_10_7));
  fa fa_h_u_wallace_cla16_fa62_out(.a(h_u_wallace_cla16_fa61_or0[0]), .b(h_u_wallace_cla16_and_11_6[0]), .cin(h_u_wallace_cla16_and_10_7[0]), .fa_xor1(h_u_wallace_cla16_fa62_xor1), .fa_or0(h_u_wallace_cla16_fa62_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_7(.a(a[11]), .b(b[7]), .out(h_u_wallace_cla16_and_11_7));
  and_gate and_gate_h_u_wallace_cla16_and_10_8(.a(a[10]), .b(b[8]), .out(h_u_wallace_cla16_and_10_8));
  fa fa_h_u_wallace_cla16_fa63_out(.a(h_u_wallace_cla16_fa62_or0[0]), .b(h_u_wallace_cla16_and_11_7[0]), .cin(h_u_wallace_cla16_and_10_8[0]), .fa_xor1(h_u_wallace_cla16_fa63_xor1), .fa_or0(h_u_wallace_cla16_fa63_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_8(.a(a[11]), .b(b[8]), .out(h_u_wallace_cla16_and_11_8));
  and_gate and_gate_h_u_wallace_cla16_and_10_9(.a(a[10]), .b(b[9]), .out(h_u_wallace_cla16_and_10_9));
  fa fa_h_u_wallace_cla16_fa64_out(.a(h_u_wallace_cla16_fa63_or0[0]), .b(h_u_wallace_cla16_and_11_8[0]), .cin(h_u_wallace_cla16_and_10_9[0]), .fa_xor1(h_u_wallace_cla16_fa64_xor1), .fa_or0(h_u_wallace_cla16_fa64_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_9(.a(a[11]), .b(b[9]), .out(h_u_wallace_cla16_and_11_9));
  and_gate and_gate_h_u_wallace_cla16_and_10_10(.a(a[10]), .b(b[10]), .out(h_u_wallace_cla16_and_10_10));
  fa fa_h_u_wallace_cla16_fa65_out(.a(h_u_wallace_cla16_fa64_or0[0]), .b(h_u_wallace_cla16_and_11_9[0]), .cin(h_u_wallace_cla16_and_10_10[0]), .fa_xor1(h_u_wallace_cla16_fa65_xor1), .fa_or0(h_u_wallace_cla16_fa65_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_10(.a(a[11]), .b(b[10]), .out(h_u_wallace_cla16_and_11_10));
  and_gate and_gate_h_u_wallace_cla16_and_10_11(.a(a[10]), .b(b[11]), .out(h_u_wallace_cla16_and_10_11));
  fa fa_h_u_wallace_cla16_fa66_out(.a(h_u_wallace_cla16_fa65_or0[0]), .b(h_u_wallace_cla16_and_11_10[0]), .cin(h_u_wallace_cla16_and_10_11[0]), .fa_xor1(h_u_wallace_cla16_fa66_xor1), .fa_or0(h_u_wallace_cla16_fa66_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_11(.a(a[11]), .b(b[11]), .out(h_u_wallace_cla16_and_11_11));
  and_gate and_gate_h_u_wallace_cla16_and_10_12(.a(a[10]), .b(b[12]), .out(h_u_wallace_cla16_and_10_12));
  fa fa_h_u_wallace_cla16_fa67_out(.a(h_u_wallace_cla16_fa66_or0[0]), .b(h_u_wallace_cla16_and_11_11[0]), .cin(h_u_wallace_cla16_and_10_12[0]), .fa_xor1(h_u_wallace_cla16_fa67_xor1), .fa_or0(h_u_wallace_cla16_fa67_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_12(.a(a[11]), .b(b[12]), .out(h_u_wallace_cla16_and_11_12));
  and_gate and_gate_h_u_wallace_cla16_and_10_13(.a(a[10]), .b(b[13]), .out(h_u_wallace_cla16_and_10_13));
  fa fa_h_u_wallace_cla16_fa68_out(.a(h_u_wallace_cla16_fa67_or0[0]), .b(h_u_wallace_cla16_and_11_12[0]), .cin(h_u_wallace_cla16_and_10_13[0]), .fa_xor1(h_u_wallace_cla16_fa68_xor1), .fa_or0(h_u_wallace_cla16_fa68_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_13(.a(a[11]), .b(b[13]), .out(h_u_wallace_cla16_and_11_13));
  and_gate and_gate_h_u_wallace_cla16_and_10_14(.a(a[10]), .b(b[14]), .out(h_u_wallace_cla16_and_10_14));
  fa fa_h_u_wallace_cla16_fa69_out(.a(h_u_wallace_cla16_fa68_or0[0]), .b(h_u_wallace_cla16_and_11_13[0]), .cin(h_u_wallace_cla16_and_10_14[0]), .fa_xor1(h_u_wallace_cla16_fa69_xor1), .fa_or0(h_u_wallace_cla16_fa69_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_14(.a(a[11]), .b(b[14]), .out(h_u_wallace_cla16_and_11_14));
  and_gate and_gate_h_u_wallace_cla16_and_10_15(.a(a[10]), .b(b[15]), .out(h_u_wallace_cla16_and_10_15));
  fa fa_h_u_wallace_cla16_fa70_out(.a(h_u_wallace_cla16_fa69_or0[0]), .b(h_u_wallace_cla16_and_11_14[0]), .cin(h_u_wallace_cla16_and_10_15[0]), .fa_xor1(h_u_wallace_cla16_fa70_xor1), .fa_or0(h_u_wallace_cla16_fa70_or0));
  and_gate and_gate_h_u_wallace_cla16_and_11_15(.a(a[11]), .b(b[15]), .out(h_u_wallace_cla16_and_11_15));
  fa fa_h_u_wallace_cla16_fa71_out(.a(h_u_wallace_cla16_fa70_or0[0]), .b(h_u_wallace_cla16_and_11_15[0]), .cin(h_u_wallace_cla16_fa23_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa71_xor1), .fa_or0(h_u_wallace_cla16_fa71_or0));
  ha ha_h_u_wallace_cla16_ha3_out(.a(h_u_wallace_cla16_fa2_xor1[0]), .b(h_u_wallace_cla16_fa27_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha3_xor0), .ha_and0(h_u_wallace_cla16_ha3_and0));
  and_gate and_gate_h_u_wallace_cla16_and_0_6(.a(a[0]), .b(b[6]), .out(h_u_wallace_cla16_and_0_6));
  fa fa_h_u_wallace_cla16_fa72_out(.a(h_u_wallace_cla16_ha3_and0[0]), .b(h_u_wallace_cla16_and_0_6[0]), .cin(h_u_wallace_cla16_fa3_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa72_xor1), .fa_or0(h_u_wallace_cla16_fa72_or0));
  and_gate and_gate_h_u_wallace_cla16_and_1_6(.a(a[1]), .b(b[6]), .out(h_u_wallace_cla16_and_1_6));
  and_gate and_gate_h_u_wallace_cla16_and_0_7(.a(a[0]), .b(b[7]), .out(h_u_wallace_cla16_and_0_7));
  fa fa_h_u_wallace_cla16_fa73_out(.a(h_u_wallace_cla16_fa72_or0[0]), .b(h_u_wallace_cla16_and_1_6[0]), .cin(h_u_wallace_cla16_and_0_7[0]), .fa_xor1(h_u_wallace_cla16_fa73_xor1), .fa_or0(h_u_wallace_cla16_fa73_or0));
  and_gate and_gate_h_u_wallace_cla16_and_2_6(.a(a[2]), .b(b[6]), .out(h_u_wallace_cla16_and_2_6));
  and_gate and_gate_h_u_wallace_cla16_and_1_7(.a(a[1]), .b(b[7]), .out(h_u_wallace_cla16_and_1_7));
  fa fa_h_u_wallace_cla16_fa74_out(.a(h_u_wallace_cla16_fa73_or0[0]), .b(h_u_wallace_cla16_and_2_6[0]), .cin(h_u_wallace_cla16_and_1_7[0]), .fa_xor1(h_u_wallace_cla16_fa74_xor1), .fa_or0(h_u_wallace_cla16_fa74_or0));
  and_gate and_gate_h_u_wallace_cla16_and_3_6(.a(a[3]), .b(b[6]), .out(h_u_wallace_cla16_and_3_6));
  and_gate and_gate_h_u_wallace_cla16_and_2_7(.a(a[2]), .b(b[7]), .out(h_u_wallace_cla16_and_2_7));
  fa fa_h_u_wallace_cla16_fa75_out(.a(h_u_wallace_cla16_fa74_or0[0]), .b(h_u_wallace_cla16_and_3_6[0]), .cin(h_u_wallace_cla16_and_2_7[0]), .fa_xor1(h_u_wallace_cla16_fa75_xor1), .fa_or0(h_u_wallace_cla16_fa75_or0));
  and_gate and_gate_h_u_wallace_cla16_and_4_6(.a(a[4]), .b(b[6]), .out(h_u_wallace_cla16_and_4_6));
  and_gate and_gate_h_u_wallace_cla16_and_3_7(.a(a[3]), .b(b[7]), .out(h_u_wallace_cla16_and_3_7));
  fa fa_h_u_wallace_cla16_fa76_out(.a(h_u_wallace_cla16_fa75_or0[0]), .b(h_u_wallace_cla16_and_4_6[0]), .cin(h_u_wallace_cla16_and_3_7[0]), .fa_xor1(h_u_wallace_cla16_fa76_xor1), .fa_or0(h_u_wallace_cla16_fa76_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_6(.a(a[5]), .b(b[6]), .out(h_u_wallace_cla16_and_5_6));
  and_gate and_gate_h_u_wallace_cla16_and_4_7(.a(a[4]), .b(b[7]), .out(h_u_wallace_cla16_and_4_7));
  fa fa_h_u_wallace_cla16_fa77_out(.a(h_u_wallace_cla16_fa76_or0[0]), .b(h_u_wallace_cla16_and_5_6[0]), .cin(h_u_wallace_cla16_and_4_7[0]), .fa_xor1(h_u_wallace_cla16_fa77_xor1), .fa_or0(h_u_wallace_cla16_fa77_or0));
  and_gate and_gate_h_u_wallace_cla16_and_6_6(.a(a[6]), .b(b[6]), .out(h_u_wallace_cla16_and_6_6));
  and_gate and_gate_h_u_wallace_cla16_and_5_7(.a(a[5]), .b(b[7]), .out(h_u_wallace_cla16_and_5_7));
  fa fa_h_u_wallace_cla16_fa78_out(.a(h_u_wallace_cla16_fa77_or0[0]), .b(h_u_wallace_cla16_and_6_6[0]), .cin(h_u_wallace_cla16_and_5_7[0]), .fa_xor1(h_u_wallace_cla16_fa78_xor1), .fa_or0(h_u_wallace_cla16_fa78_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_6(.a(a[7]), .b(b[6]), .out(h_u_wallace_cla16_and_7_6));
  and_gate and_gate_h_u_wallace_cla16_and_6_7(.a(a[6]), .b(b[7]), .out(h_u_wallace_cla16_and_6_7));
  fa fa_h_u_wallace_cla16_fa79_out(.a(h_u_wallace_cla16_fa78_or0[0]), .b(h_u_wallace_cla16_and_7_6[0]), .cin(h_u_wallace_cla16_and_6_7[0]), .fa_xor1(h_u_wallace_cla16_fa79_xor1), .fa_or0(h_u_wallace_cla16_fa79_or0));
  and_gate and_gate_h_u_wallace_cla16_and_8_6(.a(a[8]), .b(b[6]), .out(h_u_wallace_cla16_and_8_6));
  and_gate and_gate_h_u_wallace_cla16_and_7_7(.a(a[7]), .b(b[7]), .out(h_u_wallace_cla16_and_7_7));
  fa fa_h_u_wallace_cla16_fa80_out(.a(h_u_wallace_cla16_fa79_or0[0]), .b(h_u_wallace_cla16_and_8_6[0]), .cin(h_u_wallace_cla16_and_7_7[0]), .fa_xor1(h_u_wallace_cla16_fa80_xor1), .fa_or0(h_u_wallace_cla16_fa80_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_6(.a(a[9]), .b(b[6]), .out(h_u_wallace_cla16_and_9_6));
  and_gate and_gate_h_u_wallace_cla16_and_8_7(.a(a[8]), .b(b[7]), .out(h_u_wallace_cla16_and_8_7));
  fa fa_h_u_wallace_cla16_fa81_out(.a(h_u_wallace_cla16_fa80_or0[0]), .b(h_u_wallace_cla16_and_9_6[0]), .cin(h_u_wallace_cla16_and_8_7[0]), .fa_xor1(h_u_wallace_cla16_fa81_xor1), .fa_or0(h_u_wallace_cla16_fa81_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_7(.a(a[9]), .b(b[7]), .out(h_u_wallace_cla16_and_9_7));
  and_gate and_gate_h_u_wallace_cla16_and_8_8(.a(a[8]), .b(b[8]), .out(h_u_wallace_cla16_and_8_8));
  fa fa_h_u_wallace_cla16_fa82_out(.a(h_u_wallace_cla16_fa81_or0[0]), .b(h_u_wallace_cla16_and_9_7[0]), .cin(h_u_wallace_cla16_and_8_8[0]), .fa_xor1(h_u_wallace_cla16_fa82_xor1), .fa_or0(h_u_wallace_cla16_fa82_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_8(.a(a[9]), .b(b[8]), .out(h_u_wallace_cla16_and_9_8));
  and_gate and_gate_h_u_wallace_cla16_and_8_9(.a(a[8]), .b(b[9]), .out(h_u_wallace_cla16_and_8_9));
  fa fa_h_u_wallace_cla16_fa83_out(.a(h_u_wallace_cla16_fa82_or0[0]), .b(h_u_wallace_cla16_and_9_8[0]), .cin(h_u_wallace_cla16_and_8_9[0]), .fa_xor1(h_u_wallace_cla16_fa83_xor1), .fa_or0(h_u_wallace_cla16_fa83_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_9(.a(a[9]), .b(b[9]), .out(h_u_wallace_cla16_and_9_9));
  and_gate and_gate_h_u_wallace_cla16_and_8_10(.a(a[8]), .b(b[10]), .out(h_u_wallace_cla16_and_8_10));
  fa fa_h_u_wallace_cla16_fa84_out(.a(h_u_wallace_cla16_fa83_or0[0]), .b(h_u_wallace_cla16_and_9_9[0]), .cin(h_u_wallace_cla16_and_8_10[0]), .fa_xor1(h_u_wallace_cla16_fa84_xor1), .fa_or0(h_u_wallace_cla16_fa84_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_10(.a(a[9]), .b(b[10]), .out(h_u_wallace_cla16_and_9_10));
  and_gate and_gate_h_u_wallace_cla16_and_8_11(.a(a[8]), .b(b[11]), .out(h_u_wallace_cla16_and_8_11));
  fa fa_h_u_wallace_cla16_fa85_out(.a(h_u_wallace_cla16_fa84_or0[0]), .b(h_u_wallace_cla16_and_9_10[0]), .cin(h_u_wallace_cla16_and_8_11[0]), .fa_xor1(h_u_wallace_cla16_fa85_xor1), .fa_or0(h_u_wallace_cla16_fa85_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_11(.a(a[9]), .b(b[11]), .out(h_u_wallace_cla16_and_9_11));
  and_gate and_gate_h_u_wallace_cla16_and_8_12(.a(a[8]), .b(b[12]), .out(h_u_wallace_cla16_and_8_12));
  fa fa_h_u_wallace_cla16_fa86_out(.a(h_u_wallace_cla16_fa85_or0[0]), .b(h_u_wallace_cla16_and_9_11[0]), .cin(h_u_wallace_cla16_and_8_12[0]), .fa_xor1(h_u_wallace_cla16_fa86_xor1), .fa_or0(h_u_wallace_cla16_fa86_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_12(.a(a[9]), .b(b[12]), .out(h_u_wallace_cla16_and_9_12));
  and_gate and_gate_h_u_wallace_cla16_and_8_13(.a(a[8]), .b(b[13]), .out(h_u_wallace_cla16_and_8_13));
  fa fa_h_u_wallace_cla16_fa87_out(.a(h_u_wallace_cla16_fa86_or0[0]), .b(h_u_wallace_cla16_and_9_12[0]), .cin(h_u_wallace_cla16_and_8_13[0]), .fa_xor1(h_u_wallace_cla16_fa87_xor1), .fa_or0(h_u_wallace_cla16_fa87_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_13(.a(a[9]), .b(b[13]), .out(h_u_wallace_cla16_and_9_13));
  and_gate and_gate_h_u_wallace_cla16_and_8_14(.a(a[8]), .b(b[14]), .out(h_u_wallace_cla16_and_8_14));
  fa fa_h_u_wallace_cla16_fa88_out(.a(h_u_wallace_cla16_fa87_or0[0]), .b(h_u_wallace_cla16_and_9_13[0]), .cin(h_u_wallace_cla16_and_8_14[0]), .fa_xor1(h_u_wallace_cla16_fa88_xor1), .fa_or0(h_u_wallace_cla16_fa88_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_14(.a(a[9]), .b(b[14]), .out(h_u_wallace_cla16_and_9_14));
  and_gate and_gate_h_u_wallace_cla16_and_8_15(.a(a[8]), .b(b[15]), .out(h_u_wallace_cla16_and_8_15));
  fa fa_h_u_wallace_cla16_fa89_out(.a(h_u_wallace_cla16_fa88_or0[0]), .b(h_u_wallace_cla16_and_9_14[0]), .cin(h_u_wallace_cla16_and_8_15[0]), .fa_xor1(h_u_wallace_cla16_fa89_xor1), .fa_or0(h_u_wallace_cla16_fa89_or0));
  and_gate and_gate_h_u_wallace_cla16_and_9_15(.a(a[9]), .b(b[15]), .out(h_u_wallace_cla16_and_9_15));
  fa fa_h_u_wallace_cla16_fa90_out(.a(h_u_wallace_cla16_fa89_or0[0]), .b(h_u_wallace_cla16_and_9_15[0]), .cin(h_u_wallace_cla16_fa21_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa90_xor1), .fa_or0(h_u_wallace_cla16_fa90_or0));
  fa fa_h_u_wallace_cla16_fa91_out(.a(h_u_wallace_cla16_fa90_or0[0]), .b(h_u_wallace_cla16_fa22_xor1[0]), .cin(h_u_wallace_cla16_fa47_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa91_xor1), .fa_or0(h_u_wallace_cla16_fa91_or0));
  ha ha_h_u_wallace_cla16_ha4_out(.a(h_u_wallace_cla16_fa28_xor1[0]), .b(h_u_wallace_cla16_fa51_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha4_xor0), .ha_and0(h_u_wallace_cla16_ha4_and0));
  fa fa_h_u_wallace_cla16_fa92_out(.a(h_u_wallace_cla16_ha4_and0[0]), .b(h_u_wallace_cla16_fa4_xor1[0]), .cin(h_u_wallace_cla16_fa29_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa92_xor1), .fa_or0(h_u_wallace_cla16_fa92_or0));
  and_gate and_gate_h_u_wallace_cla16_and_0_8(.a(a[0]), .b(b[8]), .out(h_u_wallace_cla16_and_0_8));
  fa fa_h_u_wallace_cla16_fa93_out(.a(h_u_wallace_cla16_fa92_or0[0]), .b(h_u_wallace_cla16_and_0_8[0]), .cin(h_u_wallace_cla16_fa5_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa93_xor1), .fa_or0(h_u_wallace_cla16_fa93_or0));
  and_gate and_gate_h_u_wallace_cla16_and_1_8(.a(a[1]), .b(b[8]), .out(h_u_wallace_cla16_and_1_8));
  and_gate and_gate_h_u_wallace_cla16_and_0_9(.a(a[0]), .b(b[9]), .out(h_u_wallace_cla16_and_0_9));
  fa fa_h_u_wallace_cla16_fa94_out(.a(h_u_wallace_cla16_fa93_or0[0]), .b(h_u_wallace_cla16_and_1_8[0]), .cin(h_u_wallace_cla16_and_0_9[0]), .fa_xor1(h_u_wallace_cla16_fa94_xor1), .fa_or0(h_u_wallace_cla16_fa94_or0));
  and_gate and_gate_h_u_wallace_cla16_and_2_8(.a(a[2]), .b(b[8]), .out(h_u_wallace_cla16_and_2_8));
  and_gate and_gate_h_u_wallace_cla16_and_1_9(.a(a[1]), .b(b[9]), .out(h_u_wallace_cla16_and_1_9));
  fa fa_h_u_wallace_cla16_fa95_out(.a(h_u_wallace_cla16_fa94_or0[0]), .b(h_u_wallace_cla16_and_2_8[0]), .cin(h_u_wallace_cla16_and_1_9[0]), .fa_xor1(h_u_wallace_cla16_fa95_xor1), .fa_or0(h_u_wallace_cla16_fa95_or0));
  and_gate and_gate_h_u_wallace_cla16_and_3_8(.a(a[3]), .b(b[8]), .out(h_u_wallace_cla16_and_3_8));
  and_gate and_gate_h_u_wallace_cla16_and_2_9(.a(a[2]), .b(b[9]), .out(h_u_wallace_cla16_and_2_9));
  fa fa_h_u_wallace_cla16_fa96_out(.a(h_u_wallace_cla16_fa95_or0[0]), .b(h_u_wallace_cla16_and_3_8[0]), .cin(h_u_wallace_cla16_and_2_9[0]), .fa_xor1(h_u_wallace_cla16_fa96_xor1), .fa_or0(h_u_wallace_cla16_fa96_or0));
  and_gate and_gate_h_u_wallace_cla16_and_4_8(.a(a[4]), .b(b[8]), .out(h_u_wallace_cla16_and_4_8));
  and_gate and_gate_h_u_wallace_cla16_and_3_9(.a(a[3]), .b(b[9]), .out(h_u_wallace_cla16_and_3_9));
  fa fa_h_u_wallace_cla16_fa97_out(.a(h_u_wallace_cla16_fa96_or0[0]), .b(h_u_wallace_cla16_and_4_8[0]), .cin(h_u_wallace_cla16_and_3_9[0]), .fa_xor1(h_u_wallace_cla16_fa97_xor1), .fa_or0(h_u_wallace_cla16_fa97_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_8(.a(a[5]), .b(b[8]), .out(h_u_wallace_cla16_and_5_8));
  and_gate and_gate_h_u_wallace_cla16_and_4_9(.a(a[4]), .b(b[9]), .out(h_u_wallace_cla16_and_4_9));
  fa fa_h_u_wallace_cla16_fa98_out(.a(h_u_wallace_cla16_fa97_or0[0]), .b(h_u_wallace_cla16_and_5_8[0]), .cin(h_u_wallace_cla16_and_4_9[0]), .fa_xor1(h_u_wallace_cla16_fa98_xor1), .fa_or0(h_u_wallace_cla16_fa98_or0));
  and_gate and_gate_h_u_wallace_cla16_and_6_8(.a(a[6]), .b(b[8]), .out(h_u_wallace_cla16_and_6_8));
  and_gate and_gate_h_u_wallace_cla16_and_5_9(.a(a[5]), .b(b[9]), .out(h_u_wallace_cla16_and_5_9));
  fa fa_h_u_wallace_cla16_fa99_out(.a(h_u_wallace_cla16_fa98_or0[0]), .b(h_u_wallace_cla16_and_6_8[0]), .cin(h_u_wallace_cla16_and_5_9[0]), .fa_xor1(h_u_wallace_cla16_fa99_xor1), .fa_or0(h_u_wallace_cla16_fa99_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_8(.a(a[7]), .b(b[8]), .out(h_u_wallace_cla16_and_7_8));
  and_gate and_gate_h_u_wallace_cla16_and_6_9(.a(a[6]), .b(b[9]), .out(h_u_wallace_cla16_and_6_9));
  fa fa_h_u_wallace_cla16_fa100_out(.a(h_u_wallace_cla16_fa99_or0[0]), .b(h_u_wallace_cla16_and_7_8[0]), .cin(h_u_wallace_cla16_and_6_9[0]), .fa_xor1(h_u_wallace_cla16_fa100_xor1), .fa_or0(h_u_wallace_cla16_fa100_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_9(.a(a[7]), .b(b[9]), .out(h_u_wallace_cla16_and_7_9));
  and_gate and_gate_h_u_wallace_cla16_and_6_10(.a(a[6]), .b(b[10]), .out(h_u_wallace_cla16_and_6_10));
  fa fa_h_u_wallace_cla16_fa101_out(.a(h_u_wallace_cla16_fa100_or0[0]), .b(h_u_wallace_cla16_and_7_9[0]), .cin(h_u_wallace_cla16_and_6_10[0]), .fa_xor1(h_u_wallace_cla16_fa101_xor1), .fa_or0(h_u_wallace_cla16_fa101_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_10(.a(a[7]), .b(b[10]), .out(h_u_wallace_cla16_and_7_10));
  and_gate and_gate_h_u_wallace_cla16_and_6_11(.a(a[6]), .b(b[11]), .out(h_u_wallace_cla16_and_6_11));
  fa fa_h_u_wallace_cla16_fa102_out(.a(h_u_wallace_cla16_fa101_or0[0]), .b(h_u_wallace_cla16_and_7_10[0]), .cin(h_u_wallace_cla16_and_6_11[0]), .fa_xor1(h_u_wallace_cla16_fa102_xor1), .fa_or0(h_u_wallace_cla16_fa102_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_11(.a(a[7]), .b(b[11]), .out(h_u_wallace_cla16_and_7_11));
  and_gate and_gate_h_u_wallace_cla16_and_6_12(.a(a[6]), .b(b[12]), .out(h_u_wallace_cla16_and_6_12));
  fa fa_h_u_wallace_cla16_fa103_out(.a(h_u_wallace_cla16_fa102_or0[0]), .b(h_u_wallace_cla16_and_7_11[0]), .cin(h_u_wallace_cla16_and_6_12[0]), .fa_xor1(h_u_wallace_cla16_fa103_xor1), .fa_or0(h_u_wallace_cla16_fa103_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_12(.a(a[7]), .b(b[12]), .out(h_u_wallace_cla16_and_7_12));
  and_gate and_gate_h_u_wallace_cla16_and_6_13(.a(a[6]), .b(b[13]), .out(h_u_wallace_cla16_and_6_13));
  fa fa_h_u_wallace_cla16_fa104_out(.a(h_u_wallace_cla16_fa103_or0[0]), .b(h_u_wallace_cla16_and_7_12[0]), .cin(h_u_wallace_cla16_and_6_13[0]), .fa_xor1(h_u_wallace_cla16_fa104_xor1), .fa_or0(h_u_wallace_cla16_fa104_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_13(.a(a[7]), .b(b[13]), .out(h_u_wallace_cla16_and_7_13));
  and_gate and_gate_h_u_wallace_cla16_and_6_14(.a(a[6]), .b(b[14]), .out(h_u_wallace_cla16_and_6_14));
  fa fa_h_u_wallace_cla16_fa105_out(.a(h_u_wallace_cla16_fa104_or0[0]), .b(h_u_wallace_cla16_and_7_13[0]), .cin(h_u_wallace_cla16_and_6_14[0]), .fa_xor1(h_u_wallace_cla16_fa105_xor1), .fa_or0(h_u_wallace_cla16_fa105_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_14(.a(a[7]), .b(b[14]), .out(h_u_wallace_cla16_and_7_14));
  and_gate and_gate_h_u_wallace_cla16_and_6_15(.a(a[6]), .b(b[15]), .out(h_u_wallace_cla16_and_6_15));
  fa fa_h_u_wallace_cla16_fa106_out(.a(h_u_wallace_cla16_fa105_or0[0]), .b(h_u_wallace_cla16_and_7_14[0]), .cin(h_u_wallace_cla16_and_6_15[0]), .fa_xor1(h_u_wallace_cla16_fa106_xor1), .fa_or0(h_u_wallace_cla16_fa106_or0));
  and_gate and_gate_h_u_wallace_cla16_and_7_15(.a(a[7]), .b(b[15]), .out(h_u_wallace_cla16_and_7_15));
  fa fa_h_u_wallace_cla16_fa107_out(.a(h_u_wallace_cla16_fa106_or0[0]), .b(h_u_wallace_cla16_and_7_15[0]), .cin(h_u_wallace_cla16_fa19_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa107_xor1), .fa_or0(h_u_wallace_cla16_fa107_or0));
  fa fa_h_u_wallace_cla16_fa108_out(.a(h_u_wallace_cla16_fa107_or0[0]), .b(h_u_wallace_cla16_fa20_xor1[0]), .cin(h_u_wallace_cla16_fa45_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa108_xor1), .fa_or0(h_u_wallace_cla16_fa108_or0));
  fa fa_h_u_wallace_cla16_fa109_out(.a(h_u_wallace_cla16_fa108_or0[0]), .b(h_u_wallace_cla16_fa46_xor1[0]), .cin(h_u_wallace_cla16_fa69_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa109_xor1), .fa_or0(h_u_wallace_cla16_fa109_or0));
  ha ha_h_u_wallace_cla16_ha5_out(.a(h_u_wallace_cla16_fa52_xor1[0]), .b(h_u_wallace_cla16_fa73_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha5_xor0), .ha_and0(h_u_wallace_cla16_ha5_and0));
  fa fa_h_u_wallace_cla16_fa110_out(.a(h_u_wallace_cla16_ha5_and0[0]), .b(h_u_wallace_cla16_fa30_xor1[0]), .cin(h_u_wallace_cla16_fa53_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa110_xor1), .fa_or0(h_u_wallace_cla16_fa110_or0));
  fa fa_h_u_wallace_cla16_fa111_out(.a(h_u_wallace_cla16_fa110_or0[0]), .b(h_u_wallace_cla16_fa6_xor1[0]), .cin(h_u_wallace_cla16_fa31_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa111_xor1), .fa_or0(h_u_wallace_cla16_fa111_or0));
  and_gate and_gate_h_u_wallace_cla16_and_0_10(.a(a[0]), .b(b[10]), .out(h_u_wallace_cla16_and_0_10));
  fa fa_h_u_wallace_cla16_fa112_out(.a(h_u_wallace_cla16_fa111_or0[0]), .b(h_u_wallace_cla16_and_0_10[0]), .cin(h_u_wallace_cla16_fa7_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa112_xor1), .fa_or0(h_u_wallace_cla16_fa112_or0));
  and_gate and_gate_h_u_wallace_cla16_and_1_10(.a(a[1]), .b(b[10]), .out(h_u_wallace_cla16_and_1_10));
  and_gate and_gate_h_u_wallace_cla16_and_0_11(.a(a[0]), .b(b[11]), .out(h_u_wallace_cla16_and_0_11));
  fa fa_h_u_wallace_cla16_fa113_out(.a(h_u_wallace_cla16_fa112_or0[0]), .b(h_u_wallace_cla16_and_1_10[0]), .cin(h_u_wallace_cla16_and_0_11[0]), .fa_xor1(h_u_wallace_cla16_fa113_xor1), .fa_or0(h_u_wallace_cla16_fa113_or0));
  and_gate and_gate_h_u_wallace_cla16_and_2_10(.a(a[2]), .b(b[10]), .out(h_u_wallace_cla16_and_2_10));
  and_gate and_gate_h_u_wallace_cla16_and_1_11(.a(a[1]), .b(b[11]), .out(h_u_wallace_cla16_and_1_11));
  fa fa_h_u_wallace_cla16_fa114_out(.a(h_u_wallace_cla16_fa113_or0[0]), .b(h_u_wallace_cla16_and_2_10[0]), .cin(h_u_wallace_cla16_and_1_11[0]), .fa_xor1(h_u_wallace_cla16_fa114_xor1), .fa_or0(h_u_wallace_cla16_fa114_or0));
  and_gate and_gate_h_u_wallace_cla16_and_3_10(.a(a[3]), .b(b[10]), .out(h_u_wallace_cla16_and_3_10));
  and_gate and_gate_h_u_wallace_cla16_and_2_11(.a(a[2]), .b(b[11]), .out(h_u_wallace_cla16_and_2_11));
  fa fa_h_u_wallace_cla16_fa115_out(.a(h_u_wallace_cla16_fa114_or0[0]), .b(h_u_wallace_cla16_and_3_10[0]), .cin(h_u_wallace_cla16_and_2_11[0]), .fa_xor1(h_u_wallace_cla16_fa115_xor1), .fa_or0(h_u_wallace_cla16_fa115_or0));
  and_gate and_gate_h_u_wallace_cla16_and_4_10(.a(a[4]), .b(b[10]), .out(h_u_wallace_cla16_and_4_10));
  and_gate and_gate_h_u_wallace_cla16_and_3_11(.a(a[3]), .b(b[11]), .out(h_u_wallace_cla16_and_3_11));
  fa fa_h_u_wallace_cla16_fa116_out(.a(h_u_wallace_cla16_fa115_or0[0]), .b(h_u_wallace_cla16_and_4_10[0]), .cin(h_u_wallace_cla16_and_3_11[0]), .fa_xor1(h_u_wallace_cla16_fa116_xor1), .fa_or0(h_u_wallace_cla16_fa116_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_10(.a(a[5]), .b(b[10]), .out(h_u_wallace_cla16_and_5_10));
  and_gate and_gate_h_u_wallace_cla16_and_4_11(.a(a[4]), .b(b[11]), .out(h_u_wallace_cla16_and_4_11));
  fa fa_h_u_wallace_cla16_fa117_out(.a(h_u_wallace_cla16_fa116_or0[0]), .b(h_u_wallace_cla16_and_5_10[0]), .cin(h_u_wallace_cla16_and_4_11[0]), .fa_xor1(h_u_wallace_cla16_fa117_xor1), .fa_or0(h_u_wallace_cla16_fa117_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_11(.a(a[5]), .b(b[11]), .out(h_u_wallace_cla16_and_5_11));
  and_gate and_gate_h_u_wallace_cla16_and_4_12(.a(a[4]), .b(b[12]), .out(h_u_wallace_cla16_and_4_12));
  fa fa_h_u_wallace_cla16_fa118_out(.a(h_u_wallace_cla16_fa117_or0[0]), .b(h_u_wallace_cla16_and_5_11[0]), .cin(h_u_wallace_cla16_and_4_12[0]), .fa_xor1(h_u_wallace_cla16_fa118_xor1), .fa_or0(h_u_wallace_cla16_fa118_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_12(.a(a[5]), .b(b[12]), .out(h_u_wallace_cla16_and_5_12));
  and_gate and_gate_h_u_wallace_cla16_and_4_13(.a(a[4]), .b(b[13]), .out(h_u_wallace_cla16_and_4_13));
  fa fa_h_u_wallace_cla16_fa119_out(.a(h_u_wallace_cla16_fa118_or0[0]), .b(h_u_wallace_cla16_and_5_12[0]), .cin(h_u_wallace_cla16_and_4_13[0]), .fa_xor1(h_u_wallace_cla16_fa119_xor1), .fa_or0(h_u_wallace_cla16_fa119_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_13(.a(a[5]), .b(b[13]), .out(h_u_wallace_cla16_and_5_13));
  and_gate and_gate_h_u_wallace_cla16_and_4_14(.a(a[4]), .b(b[14]), .out(h_u_wallace_cla16_and_4_14));
  fa fa_h_u_wallace_cla16_fa120_out(.a(h_u_wallace_cla16_fa119_or0[0]), .b(h_u_wallace_cla16_and_5_13[0]), .cin(h_u_wallace_cla16_and_4_14[0]), .fa_xor1(h_u_wallace_cla16_fa120_xor1), .fa_or0(h_u_wallace_cla16_fa120_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_14(.a(a[5]), .b(b[14]), .out(h_u_wallace_cla16_and_5_14));
  and_gate and_gate_h_u_wallace_cla16_and_4_15(.a(a[4]), .b(b[15]), .out(h_u_wallace_cla16_and_4_15));
  fa fa_h_u_wallace_cla16_fa121_out(.a(h_u_wallace_cla16_fa120_or0[0]), .b(h_u_wallace_cla16_and_5_14[0]), .cin(h_u_wallace_cla16_and_4_15[0]), .fa_xor1(h_u_wallace_cla16_fa121_xor1), .fa_or0(h_u_wallace_cla16_fa121_or0));
  and_gate and_gate_h_u_wallace_cla16_and_5_15(.a(a[5]), .b(b[15]), .out(h_u_wallace_cla16_and_5_15));
  fa fa_h_u_wallace_cla16_fa122_out(.a(h_u_wallace_cla16_fa121_or0[0]), .b(h_u_wallace_cla16_and_5_15[0]), .cin(h_u_wallace_cla16_fa17_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa122_xor1), .fa_or0(h_u_wallace_cla16_fa122_or0));
  fa fa_h_u_wallace_cla16_fa123_out(.a(h_u_wallace_cla16_fa122_or0[0]), .b(h_u_wallace_cla16_fa18_xor1[0]), .cin(h_u_wallace_cla16_fa43_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa123_xor1), .fa_or0(h_u_wallace_cla16_fa123_or0));
  fa fa_h_u_wallace_cla16_fa124_out(.a(h_u_wallace_cla16_fa123_or0[0]), .b(h_u_wallace_cla16_fa44_xor1[0]), .cin(h_u_wallace_cla16_fa67_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa124_xor1), .fa_or0(h_u_wallace_cla16_fa124_or0));
  fa fa_h_u_wallace_cla16_fa125_out(.a(h_u_wallace_cla16_fa124_or0[0]), .b(h_u_wallace_cla16_fa68_xor1[0]), .cin(h_u_wallace_cla16_fa89_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa125_xor1), .fa_or0(h_u_wallace_cla16_fa125_or0));
  ha ha_h_u_wallace_cla16_ha6_out(.a(h_u_wallace_cla16_fa74_xor1[0]), .b(h_u_wallace_cla16_fa93_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha6_xor0), .ha_and0(h_u_wallace_cla16_ha6_and0));
  fa fa_h_u_wallace_cla16_fa126_out(.a(h_u_wallace_cla16_ha6_and0[0]), .b(h_u_wallace_cla16_fa54_xor1[0]), .cin(h_u_wallace_cla16_fa75_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa126_xor1), .fa_or0(h_u_wallace_cla16_fa126_or0));
  fa fa_h_u_wallace_cla16_fa127_out(.a(h_u_wallace_cla16_fa126_or0[0]), .b(h_u_wallace_cla16_fa32_xor1[0]), .cin(h_u_wallace_cla16_fa55_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa127_xor1), .fa_or0(h_u_wallace_cla16_fa127_or0));
  fa fa_h_u_wallace_cla16_fa128_out(.a(h_u_wallace_cla16_fa127_or0[0]), .b(h_u_wallace_cla16_fa8_xor1[0]), .cin(h_u_wallace_cla16_fa33_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa128_xor1), .fa_or0(h_u_wallace_cla16_fa128_or0));
  and_gate and_gate_h_u_wallace_cla16_and_0_12(.a(a[0]), .b(b[12]), .out(h_u_wallace_cla16_and_0_12));
  fa fa_h_u_wallace_cla16_fa129_out(.a(h_u_wallace_cla16_fa128_or0[0]), .b(h_u_wallace_cla16_and_0_12[0]), .cin(h_u_wallace_cla16_fa9_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa129_xor1), .fa_or0(h_u_wallace_cla16_fa129_or0));
  and_gate and_gate_h_u_wallace_cla16_and_1_12(.a(a[1]), .b(b[12]), .out(h_u_wallace_cla16_and_1_12));
  and_gate and_gate_h_u_wallace_cla16_and_0_13(.a(a[0]), .b(b[13]), .out(h_u_wallace_cla16_and_0_13));
  fa fa_h_u_wallace_cla16_fa130_out(.a(h_u_wallace_cla16_fa129_or0[0]), .b(h_u_wallace_cla16_and_1_12[0]), .cin(h_u_wallace_cla16_and_0_13[0]), .fa_xor1(h_u_wallace_cla16_fa130_xor1), .fa_or0(h_u_wallace_cla16_fa130_or0));
  and_gate and_gate_h_u_wallace_cla16_and_2_12(.a(a[2]), .b(b[12]), .out(h_u_wallace_cla16_and_2_12));
  and_gate and_gate_h_u_wallace_cla16_and_1_13(.a(a[1]), .b(b[13]), .out(h_u_wallace_cla16_and_1_13));
  fa fa_h_u_wallace_cla16_fa131_out(.a(h_u_wallace_cla16_fa130_or0[0]), .b(h_u_wallace_cla16_and_2_12[0]), .cin(h_u_wallace_cla16_and_1_13[0]), .fa_xor1(h_u_wallace_cla16_fa131_xor1), .fa_or0(h_u_wallace_cla16_fa131_or0));
  and_gate and_gate_h_u_wallace_cla16_and_3_12(.a(a[3]), .b(b[12]), .out(h_u_wallace_cla16_and_3_12));
  and_gate and_gate_h_u_wallace_cla16_and_2_13(.a(a[2]), .b(b[13]), .out(h_u_wallace_cla16_and_2_13));
  fa fa_h_u_wallace_cla16_fa132_out(.a(h_u_wallace_cla16_fa131_or0[0]), .b(h_u_wallace_cla16_and_3_12[0]), .cin(h_u_wallace_cla16_and_2_13[0]), .fa_xor1(h_u_wallace_cla16_fa132_xor1), .fa_or0(h_u_wallace_cla16_fa132_or0));
  and_gate and_gate_h_u_wallace_cla16_and_3_13(.a(a[3]), .b(b[13]), .out(h_u_wallace_cla16_and_3_13));
  and_gate and_gate_h_u_wallace_cla16_and_2_14(.a(a[2]), .b(b[14]), .out(h_u_wallace_cla16_and_2_14));
  fa fa_h_u_wallace_cla16_fa133_out(.a(h_u_wallace_cla16_fa132_or0[0]), .b(h_u_wallace_cla16_and_3_13[0]), .cin(h_u_wallace_cla16_and_2_14[0]), .fa_xor1(h_u_wallace_cla16_fa133_xor1), .fa_or0(h_u_wallace_cla16_fa133_or0));
  and_gate and_gate_h_u_wallace_cla16_and_3_14(.a(a[3]), .b(b[14]), .out(h_u_wallace_cla16_and_3_14));
  and_gate and_gate_h_u_wallace_cla16_and_2_15(.a(a[2]), .b(b[15]), .out(h_u_wallace_cla16_and_2_15));
  fa fa_h_u_wallace_cla16_fa134_out(.a(h_u_wallace_cla16_fa133_or0[0]), .b(h_u_wallace_cla16_and_3_14[0]), .cin(h_u_wallace_cla16_and_2_15[0]), .fa_xor1(h_u_wallace_cla16_fa134_xor1), .fa_or0(h_u_wallace_cla16_fa134_or0));
  and_gate and_gate_h_u_wallace_cla16_and_3_15(.a(a[3]), .b(b[15]), .out(h_u_wallace_cla16_and_3_15));
  fa fa_h_u_wallace_cla16_fa135_out(.a(h_u_wallace_cla16_fa134_or0[0]), .b(h_u_wallace_cla16_and_3_15[0]), .cin(h_u_wallace_cla16_fa15_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa135_xor1), .fa_or0(h_u_wallace_cla16_fa135_or0));
  fa fa_h_u_wallace_cla16_fa136_out(.a(h_u_wallace_cla16_fa135_or0[0]), .b(h_u_wallace_cla16_fa16_xor1[0]), .cin(h_u_wallace_cla16_fa41_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa136_xor1), .fa_or0(h_u_wallace_cla16_fa136_or0));
  fa fa_h_u_wallace_cla16_fa137_out(.a(h_u_wallace_cla16_fa136_or0[0]), .b(h_u_wallace_cla16_fa42_xor1[0]), .cin(h_u_wallace_cla16_fa65_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa137_xor1), .fa_or0(h_u_wallace_cla16_fa137_or0));
  fa fa_h_u_wallace_cla16_fa138_out(.a(h_u_wallace_cla16_fa137_or0[0]), .b(h_u_wallace_cla16_fa66_xor1[0]), .cin(h_u_wallace_cla16_fa87_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa138_xor1), .fa_or0(h_u_wallace_cla16_fa138_or0));
  fa fa_h_u_wallace_cla16_fa139_out(.a(h_u_wallace_cla16_fa138_or0[0]), .b(h_u_wallace_cla16_fa88_xor1[0]), .cin(h_u_wallace_cla16_fa107_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa139_xor1), .fa_or0(h_u_wallace_cla16_fa139_or0));
  ha ha_h_u_wallace_cla16_ha7_out(.a(h_u_wallace_cla16_fa94_xor1[0]), .b(h_u_wallace_cla16_fa111_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha7_xor0), .ha_and0(h_u_wallace_cla16_ha7_and0));
  fa fa_h_u_wallace_cla16_fa140_out(.a(h_u_wallace_cla16_ha7_and0[0]), .b(h_u_wallace_cla16_fa76_xor1[0]), .cin(h_u_wallace_cla16_fa95_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa140_xor1), .fa_or0(h_u_wallace_cla16_fa140_or0));
  fa fa_h_u_wallace_cla16_fa141_out(.a(h_u_wallace_cla16_fa140_or0[0]), .b(h_u_wallace_cla16_fa56_xor1[0]), .cin(h_u_wallace_cla16_fa77_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa141_xor1), .fa_or0(h_u_wallace_cla16_fa141_or0));
  fa fa_h_u_wallace_cla16_fa142_out(.a(h_u_wallace_cla16_fa141_or0[0]), .b(h_u_wallace_cla16_fa34_xor1[0]), .cin(h_u_wallace_cla16_fa57_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa142_xor1), .fa_or0(h_u_wallace_cla16_fa142_or0));
  fa fa_h_u_wallace_cla16_fa143_out(.a(h_u_wallace_cla16_fa142_or0[0]), .b(h_u_wallace_cla16_fa10_xor1[0]), .cin(h_u_wallace_cla16_fa35_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa143_xor1), .fa_or0(h_u_wallace_cla16_fa143_or0));
  and_gate and_gate_h_u_wallace_cla16_and_0_14(.a(a[0]), .b(b[14]), .out(h_u_wallace_cla16_and_0_14));
  fa fa_h_u_wallace_cla16_fa144_out(.a(h_u_wallace_cla16_fa143_or0[0]), .b(h_u_wallace_cla16_and_0_14[0]), .cin(h_u_wallace_cla16_fa11_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa144_xor1), .fa_or0(h_u_wallace_cla16_fa144_or0));
  and_gate and_gate_h_u_wallace_cla16_and_1_14(.a(a[1]), .b(b[14]), .out(h_u_wallace_cla16_and_1_14));
  and_gate and_gate_h_u_wallace_cla16_and_0_15(.a(a[0]), .b(b[15]), .out(h_u_wallace_cla16_and_0_15));
  fa fa_h_u_wallace_cla16_fa145_out(.a(h_u_wallace_cla16_fa144_or0[0]), .b(h_u_wallace_cla16_and_1_14[0]), .cin(h_u_wallace_cla16_and_0_15[0]), .fa_xor1(h_u_wallace_cla16_fa145_xor1), .fa_or0(h_u_wallace_cla16_fa145_or0));
  and_gate and_gate_h_u_wallace_cla16_and_1_15(.a(a[1]), .b(b[15]), .out(h_u_wallace_cla16_and_1_15));
  fa fa_h_u_wallace_cla16_fa146_out(.a(h_u_wallace_cla16_fa145_or0[0]), .b(h_u_wallace_cla16_and_1_15[0]), .cin(h_u_wallace_cla16_fa13_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa146_xor1), .fa_or0(h_u_wallace_cla16_fa146_or0));
  fa fa_h_u_wallace_cla16_fa147_out(.a(h_u_wallace_cla16_fa146_or0[0]), .b(h_u_wallace_cla16_fa14_xor1[0]), .cin(h_u_wallace_cla16_fa39_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa147_xor1), .fa_or0(h_u_wallace_cla16_fa147_or0));
  fa fa_h_u_wallace_cla16_fa148_out(.a(h_u_wallace_cla16_fa147_or0[0]), .b(h_u_wallace_cla16_fa40_xor1[0]), .cin(h_u_wallace_cla16_fa63_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa148_xor1), .fa_or0(h_u_wallace_cla16_fa148_or0));
  fa fa_h_u_wallace_cla16_fa149_out(.a(h_u_wallace_cla16_fa148_or0[0]), .b(h_u_wallace_cla16_fa64_xor1[0]), .cin(h_u_wallace_cla16_fa85_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa149_xor1), .fa_or0(h_u_wallace_cla16_fa149_or0));
  fa fa_h_u_wallace_cla16_fa150_out(.a(h_u_wallace_cla16_fa149_or0[0]), .b(h_u_wallace_cla16_fa86_xor1[0]), .cin(h_u_wallace_cla16_fa105_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa150_xor1), .fa_or0(h_u_wallace_cla16_fa150_or0));
  fa fa_h_u_wallace_cla16_fa151_out(.a(h_u_wallace_cla16_fa150_or0[0]), .b(h_u_wallace_cla16_fa106_xor1[0]), .cin(h_u_wallace_cla16_fa123_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa151_xor1), .fa_or0(h_u_wallace_cla16_fa151_or0));
  ha ha_h_u_wallace_cla16_ha8_out(.a(h_u_wallace_cla16_fa112_xor1[0]), .b(h_u_wallace_cla16_fa127_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha8_xor0), .ha_and0(h_u_wallace_cla16_ha8_and0));
  fa fa_h_u_wallace_cla16_fa152_out(.a(h_u_wallace_cla16_ha8_and0[0]), .b(h_u_wallace_cla16_fa96_xor1[0]), .cin(h_u_wallace_cla16_fa113_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa152_xor1), .fa_or0(h_u_wallace_cla16_fa152_or0));
  fa fa_h_u_wallace_cla16_fa153_out(.a(h_u_wallace_cla16_fa152_or0[0]), .b(h_u_wallace_cla16_fa78_xor1[0]), .cin(h_u_wallace_cla16_fa97_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa153_xor1), .fa_or0(h_u_wallace_cla16_fa153_or0));
  fa fa_h_u_wallace_cla16_fa154_out(.a(h_u_wallace_cla16_fa153_or0[0]), .b(h_u_wallace_cla16_fa58_xor1[0]), .cin(h_u_wallace_cla16_fa79_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa154_xor1), .fa_or0(h_u_wallace_cla16_fa154_or0));
  fa fa_h_u_wallace_cla16_fa155_out(.a(h_u_wallace_cla16_fa154_or0[0]), .b(h_u_wallace_cla16_fa36_xor1[0]), .cin(h_u_wallace_cla16_fa59_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa155_xor1), .fa_or0(h_u_wallace_cla16_fa155_or0));
  fa fa_h_u_wallace_cla16_fa156_out(.a(h_u_wallace_cla16_fa155_or0[0]), .b(h_u_wallace_cla16_fa12_xor1[0]), .cin(h_u_wallace_cla16_fa37_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa156_xor1), .fa_or0(h_u_wallace_cla16_fa156_or0));
  fa fa_h_u_wallace_cla16_fa157_out(.a(h_u_wallace_cla16_fa156_or0[0]), .b(h_u_wallace_cla16_fa38_xor1[0]), .cin(h_u_wallace_cla16_fa61_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa157_xor1), .fa_or0(h_u_wallace_cla16_fa157_or0));
  fa fa_h_u_wallace_cla16_fa158_out(.a(h_u_wallace_cla16_fa157_or0[0]), .b(h_u_wallace_cla16_fa62_xor1[0]), .cin(h_u_wallace_cla16_fa83_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa158_xor1), .fa_or0(h_u_wallace_cla16_fa158_or0));
  fa fa_h_u_wallace_cla16_fa159_out(.a(h_u_wallace_cla16_fa158_or0[0]), .b(h_u_wallace_cla16_fa84_xor1[0]), .cin(h_u_wallace_cla16_fa103_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa159_xor1), .fa_or0(h_u_wallace_cla16_fa159_or0));
  fa fa_h_u_wallace_cla16_fa160_out(.a(h_u_wallace_cla16_fa159_or0[0]), .b(h_u_wallace_cla16_fa104_xor1[0]), .cin(h_u_wallace_cla16_fa121_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa160_xor1), .fa_or0(h_u_wallace_cla16_fa160_or0));
  fa fa_h_u_wallace_cla16_fa161_out(.a(h_u_wallace_cla16_fa160_or0[0]), .b(h_u_wallace_cla16_fa122_xor1[0]), .cin(h_u_wallace_cla16_fa137_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa161_xor1), .fa_or0(h_u_wallace_cla16_fa161_or0));
  ha ha_h_u_wallace_cla16_ha9_out(.a(h_u_wallace_cla16_fa128_xor1[0]), .b(h_u_wallace_cla16_fa141_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha9_xor0), .ha_and0(h_u_wallace_cla16_ha9_and0));
  fa fa_h_u_wallace_cla16_fa162_out(.a(h_u_wallace_cla16_ha9_and0[0]), .b(h_u_wallace_cla16_fa114_xor1[0]), .cin(h_u_wallace_cla16_fa129_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa162_xor1), .fa_or0(h_u_wallace_cla16_fa162_or0));
  fa fa_h_u_wallace_cla16_fa163_out(.a(h_u_wallace_cla16_fa162_or0[0]), .b(h_u_wallace_cla16_fa98_xor1[0]), .cin(h_u_wallace_cla16_fa115_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa163_xor1), .fa_or0(h_u_wallace_cla16_fa163_or0));
  fa fa_h_u_wallace_cla16_fa164_out(.a(h_u_wallace_cla16_fa163_or0[0]), .b(h_u_wallace_cla16_fa80_xor1[0]), .cin(h_u_wallace_cla16_fa99_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa164_xor1), .fa_or0(h_u_wallace_cla16_fa164_or0));
  fa fa_h_u_wallace_cla16_fa165_out(.a(h_u_wallace_cla16_fa164_or0[0]), .b(h_u_wallace_cla16_fa60_xor1[0]), .cin(h_u_wallace_cla16_fa81_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa165_xor1), .fa_or0(h_u_wallace_cla16_fa165_or0));
  fa fa_h_u_wallace_cla16_fa166_out(.a(h_u_wallace_cla16_fa165_or0[0]), .b(h_u_wallace_cla16_fa82_xor1[0]), .cin(h_u_wallace_cla16_fa101_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa166_xor1), .fa_or0(h_u_wallace_cla16_fa166_or0));
  fa fa_h_u_wallace_cla16_fa167_out(.a(h_u_wallace_cla16_fa166_or0[0]), .b(h_u_wallace_cla16_fa102_xor1[0]), .cin(h_u_wallace_cla16_fa119_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa167_xor1), .fa_or0(h_u_wallace_cla16_fa167_or0));
  fa fa_h_u_wallace_cla16_fa168_out(.a(h_u_wallace_cla16_fa167_or0[0]), .b(h_u_wallace_cla16_fa120_xor1[0]), .cin(h_u_wallace_cla16_fa135_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa168_xor1), .fa_or0(h_u_wallace_cla16_fa168_or0));
  fa fa_h_u_wallace_cla16_fa169_out(.a(h_u_wallace_cla16_fa168_or0[0]), .b(h_u_wallace_cla16_fa136_xor1[0]), .cin(h_u_wallace_cla16_fa149_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa169_xor1), .fa_or0(h_u_wallace_cla16_fa169_or0));
  ha ha_h_u_wallace_cla16_ha10_out(.a(h_u_wallace_cla16_fa142_xor1[0]), .b(h_u_wallace_cla16_fa153_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha10_xor0), .ha_and0(h_u_wallace_cla16_ha10_and0));
  fa fa_h_u_wallace_cla16_fa170_out(.a(h_u_wallace_cla16_ha10_and0[0]), .b(h_u_wallace_cla16_fa130_xor1[0]), .cin(h_u_wallace_cla16_fa143_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa170_xor1), .fa_or0(h_u_wallace_cla16_fa170_or0));
  fa fa_h_u_wallace_cla16_fa171_out(.a(h_u_wallace_cla16_fa170_or0[0]), .b(h_u_wallace_cla16_fa116_xor1[0]), .cin(h_u_wallace_cla16_fa131_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa171_xor1), .fa_or0(h_u_wallace_cla16_fa171_or0));
  fa fa_h_u_wallace_cla16_fa172_out(.a(h_u_wallace_cla16_fa171_or0[0]), .b(h_u_wallace_cla16_fa100_xor1[0]), .cin(h_u_wallace_cla16_fa117_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa172_xor1), .fa_or0(h_u_wallace_cla16_fa172_or0));
  fa fa_h_u_wallace_cla16_fa173_out(.a(h_u_wallace_cla16_fa172_or0[0]), .b(h_u_wallace_cla16_fa118_xor1[0]), .cin(h_u_wallace_cla16_fa133_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa173_xor1), .fa_or0(h_u_wallace_cla16_fa173_or0));
  fa fa_h_u_wallace_cla16_fa174_out(.a(h_u_wallace_cla16_fa173_or0[0]), .b(h_u_wallace_cla16_fa134_xor1[0]), .cin(h_u_wallace_cla16_fa147_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa174_xor1), .fa_or0(h_u_wallace_cla16_fa174_or0));
  fa fa_h_u_wallace_cla16_fa175_out(.a(h_u_wallace_cla16_fa174_or0[0]), .b(h_u_wallace_cla16_fa148_xor1[0]), .cin(h_u_wallace_cla16_fa159_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa175_xor1), .fa_or0(h_u_wallace_cla16_fa175_or0));
  ha ha_h_u_wallace_cla16_ha11_out(.a(h_u_wallace_cla16_fa154_xor1[0]), .b(h_u_wallace_cla16_fa163_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha11_xor0), .ha_and0(h_u_wallace_cla16_ha11_and0));
  fa fa_h_u_wallace_cla16_fa176_out(.a(h_u_wallace_cla16_ha11_and0[0]), .b(h_u_wallace_cla16_fa144_xor1[0]), .cin(h_u_wallace_cla16_fa155_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa176_xor1), .fa_or0(h_u_wallace_cla16_fa176_or0));
  fa fa_h_u_wallace_cla16_fa177_out(.a(h_u_wallace_cla16_fa176_or0[0]), .b(h_u_wallace_cla16_fa132_xor1[0]), .cin(h_u_wallace_cla16_fa145_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa177_xor1), .fa_or0(h_u_wallace_cla16_fa177_or0));
  fa fa_h_u_wallace_cla16_fa178_out(.a(h_u_wallace_cla16_fa177_or0[0]), .b(h_u_wallace_cla16_fa146_xor1[0]), .cin(h_u_wallace_cla16_fa157_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa178_xor1), .fa_or0(h_u_wallace_cla16_fa178_or0));
  fa fa_h_u_wallace_cla16_fa179_out(.a(h_u_wallace_cla16_fa178_or0[0]), .b(h_u_wallace_cla16_fa158_xor1[0]), .cin(h_u_wallace_cla16_fa167_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa179_xor1), .fa_or0(h_u_wallace_cla16_fa179_or0));
  ha ha_h_u_wallace_cla16_ha12_out(.a(h_u_wallace_cla16_fa164_xor1[0]), .b(h_u_wallace_cla16_fa171_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha12_xor0), .ha_and0(h_u_wallace_cla16_ha12_and0));
  fa fa_h_u_wallace_cla16_fa180_out(.a(h_u_wallace_cla16_ha12_and0[0]), .b(h_u_wallace_cla16_fa156_xor1[0]), .cin(h_u_wallace_cla16_fa165_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa180_xor1), .fa_or0(h_u_wallace_cla16_fa180_or0));
  fa fa_h_u_wallace_cla16_fa181_out(.a(h_u_wallace_cla16_fa180_or0[0]), .b(h_u_wallace_cla16_fa166_xor1[0]), .cin(h_u_wallace_cla16_fa173_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa181_xor1), .fa_or0(h_u_wallace_cla16_fa181_or0));
  ha ha_h_u_wallace_cla16_ha13_out(.a(h_u_wallace_cla16_fa172_xor1[0]), .b(h_u_wallace_cla16_fa177_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha13_xor0), .ha_and0(h_u_wallace_cla16_ha13_and0));
  ha ha_h_u_wallace_cla16_ha14_out(.a(h_u_wallace_cla16_ha13_and0[0]), .b(h_u_wallace_cla16_fa178_xor1[0]), .ha_xor0(h_u_wallace_cla16_ha14_xor0), .ha_and0(h_u_wallace_cla16_ha14_and0));
  fa fa_h_u_wallace_cla16_fa182_out(.a(h_u_wallace_cla16_ha14_and0[0]), .b(h_u_wallace_cla16_fa181_or0[0]), .cin(h_u_wallace_cla16_fa174_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa182_xor1), .fa_or0(h_u_wallace_cla16_fa182_or0));
  fa fa_h_u_wallace_cla16_fa183_out(.a(h_u_wallace_cla16_fa182_or0[0]), .b(h_u_wallace_cla16_fa179_or0[0]), .cin(h_u_wallace_cla16_fa168_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa183_xor1), .fa_or0(h_u_wallace_cla16_fa183_or0));
  fa fa_h_u_wallace_cla16_fa184_out(.a(h_u_wallace_cla16_fa183_or0[0]), .b(h_u_wallace_cla16_fa175_or0[0]), .cin(h_u_wallace_cla16_fa160_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa184_xor1), .fa_or0(h_u_wallace_cla16_fa184_or0));
  fa fa_h_u_wallace_cla16_fa185_out(.a(h_u_wallace_cla16_fa184_or0[0]), .b(h_u_wallace_cla16_fa169_or0[0]), .cin(h_u_wallace_cla16_fa150_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa185_xor1), .fa_or0(h_u_wallace_cla16_fa185_or0));
  fa fa_h_u_wallace_cla16_fa186_out(.a(h_u_wallace_cla16_fa185_or0[0]), .b(h_u_wallace_cla16_fa161_or0[0]), .cin(h_u_wallace_cla16_fa138_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa186_xor1), .fa_or0(h_u_wallace_cla16_fa186_or0));
  fa fa_h_u_wallace_cla16_fa187_out(.a(h_u_wallace_cla16_fa186_or0[0]), .b(h_u_wallace_cla16_fa151_or0[0]), .cin(h_u_wallace_cla16_fa124_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa187_xor1), .fa_or0(h_u_wallace_cla16_fa187_or0));
  fa fa_h_u_wallace_cla16_fa188_out(.a(h_u_wallace_cla16_fa187_or0[0]), .b(h_u_wallace_cla16_fa139_or0[0]), .cin(h_u_wallace_cla16_fa108_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa188_xor1), .fa_or0(h_u_wallace_cla16_fa188_or0));
  fa fa_h_u_wallace_cla16_fa189_out(.a(h_u_wallace_cla16_fa188_or0[0]), .b(h_u_wallace_cla16_fa125_or0[0]), .cin(h_u_wallace_cla16_fa90_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa189_xor1), .fa_or0(h_u_wallace_cla16_fa189_or0));
  fa fa_h_u_wallace_cla16_fa190_out(.a(h_u_wallace_cla16_fa189_or0[0]), .b(h_u_wallace_cla16_fa109_or0[0]), .cin(h_u_wallace_cla16_fa70_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa190_xor1), .fa_or0(h_u_wallace_cla16_fa190_or0));
  fa fa_h_u_wallace_cla16_fa191_out(.a(h_u_wallace_cla16_fa190_or0[0]), .b(h_u_wallace_cla16_fa91_or0[0]), .cin(h_u_wallace_cla16_fa48_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa191_xor1), .fa_or0(h_u_wallace_cla16_fa191_or0));
  fa fa_h_u_wallace_cla16_fa192_out(.a(h_u_wallace_cla16_fa191_or0[0]), .b(h_u_wallace_cla16_fa71_or0[0]), .cin(h_u_wallace_cla16_fa24_xor1[0]), .fa_xor1(h_u_wallace_cla16_fa192_xor1), .fa_or0(h_u_wallace_cla16_fa192_or0));
  and_gate and_gate_h_u_wallace_cla16_and_13_15(.a(a[13]), .b(b[15]), .out(h_u_wallace_cla16_and_13_15));
  fa fa_h_u_wallace_cla16_fa193_out(.a(h_u_wallace_cla16_fa192_or0[0]), .b(h_u_wallace_cla16_fa49_or0[0]), .cin(h_u_wallace_cla16_and_13_15[0]), .fa_xor1(h_u_wallace_cla16_fa193_xor1), .fa_or0(h_u_wallace_cla16_fa193_or0));
  and_gate and_gate_h_u_wallace_cla16_and_15_14(.a(a[15]), .b(b[14]), .out(h_u_wallace_cla16_and_15_14));
  fa fa_h_u_wallace_cla16_fa194_out(.a(h_u_wallace_cla16_fa193_or0[0]), .b(h_u_wallace_cla16_fa25_or0[0]), .cin(h_u_wallace_cla16_and_15_14[0]), .fa_xor1(h_u_wallace_cla16_fa194_xor1), .fa_or0(h_u_wallace_cla16_fa194_or0));
  and_gate and_gate_h_u_wallace_cla16_and_0_0(.a(a[0]), .b(b[0]), .out(h_u_wallace_cla16_and_0_0));
  and_gate and_gate_h_u_wallace_cla16_and_1_0(.a(a[1]), .b(b[0]), .out(h_u_wallace_cla16_and_1_0));
  and_gate and_gate_h_u_wallace_cla16_and_0_2(.a(a[0]), .b(b[2]), .out(h_u_wallace_cla16_and_0_2));
  and_gate and_gate_h_u_wallace_cla16_and_14_15(.a(a[14]), .b(b[15]), .out(h_u_wallace_cla16_and_14_15));
  and_gate and_gate_h_u_wallace_cla16_and_0_1(.a(a[0]), .b(b[1]), .out(h_u_wallace_cla16_and_0_1));
  and_gate and_gate_h_u_wallace_cla16_and_15_15(.a(a[15]), .b(b[15]), .out(h_u_wallace_cla16_and_15_15));
  assign h_u_wallace_cla16_u_cla30_a[0] = h_u_wallace_cla16_and_1_0[0];
  assign h_u_wallace_cla16_u_cla30_a[1] = h_u_wallace_cla16_and_0_2[0];
  assign h_u_wallace_cla16_u_cla30_a[2] = h_u_wallace_cla16_fa0_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[3] = h_u_wallace_cla16_fa26_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[4] = h_u_wallace_cla16_fa50_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[5] = h_u_wallace_cla16_fa72_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[6] = h_u_wallace_cla16_fa92_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[7] = h_u_wallace_cla16_fa110_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[8] = h_u_wallace_cla16_fa126_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[9] = h_u_wallace_cla16_fa140_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[10] = h_u_wallace_cla16_fa152_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[11] = h_u_wallace_cla16_fa162_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[12] = h_u_wallace_cla16_fa170_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[13] = h_u_wallace_cla16_fa176_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[14] = h_u_wallace_cla16_fa180_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[15] = h_u_wallace_cla16_fa181_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[16] = h_u_wallace_cla16_fa179_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[17] = h_u_wallace_cla16_fa175_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[18] = h_u_wallace_cla16_fa169_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[19] = h_u_wallace_cla16_fa161_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[20] = h_u_wallace_cla16_fa151_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[21] = h_u_wallace_cla16_fa139_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[22] = h_u_wallace_cla16_fa125_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[23] = h_u_wallace_cla16_fa109_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[24] = h_u_wallace_cla16_fa91_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[25] = h_u_wallace_cla16_fa71_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[26] = h_u_wallace_cla16_fa49_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[27] = h_u_wallace_cla16_fa25_xor1[0];
  assign h_u_wallace_cla16_u_cla30_a[28] = h_u_wallace_cla16_and_14_15[0];
  assign h_u_wallace_cla16_u_cla30_a[29] = h_u_wallace_cla16_fa194_or0[0];
  assign h_u_wallace_cla16_u_cla30_b[0] = h_u_wallace_cla16_and_0_1[0];
  assign h_u_wallace_cla16_u_cla30_b[1] = h_u_wallace_cla16_ha0_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[2] = h_u_wallace_cla16_ha1_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[3] = h_u_wallace_cla16_ha2_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[4] = h_u_wallace_cla16_ha3_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[5] = h_u_wallace_cla16_ha4_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[6] = h_u_wallace_cla16_ha5_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[7] = h_u_wallace_cla16_ha6_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[8] = h_u_wallace_cla16_ha7_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[9] = h_u_wallace_cla16_ha8_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[10] = h_u_wallace_cla16_ha9_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[11] = h_u_wallace_cla16_ha10_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[12] = h_u_wallace_cla16_ha11_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[13] = h_u_wallace_cla16_ha12_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[14] = h_u_wallace_cla16_ha13_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[15] = h_u_wallace_cla16_ha14_xor0[0];
  assign h_u_wallace_cla16_u_cla30_b[16] = h_u_wallace_cla16_fa182_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[17] = h_u_wallace_cla16_fa183_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[18] = h_u_wallace_cla16_fa184_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[19] = h_u_wallace_cla16_fa185_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[20] = h_u_wallace_cla16_fa186_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[21] = h_u_wallace_cla16_fa187_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[22] = h_u_wallace_cla16_fa188_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[23] = h_u_wallace_cla16_fa189_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[24] = h_u_wallace_cla16_fa190_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[25] = h_u_wallace_cla16_fa191_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[26] = h_u_wallace_cla16_fa192_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[27] = h_u_wallace_cla16_fa193_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[28] = h_u_wallace_cla16_fa194_xor1[0];
  assign h_u_wallace_cla16_u_cla30_b[29] = h_u_wallace_cla16_and_15_15[0];
  u_cla30 u_cla30_h_u_wallace_cla16_u_cla30_out(.a(h_u_wallace_cla16_u_cla30_a), .b(h_u_wallace_cla16_u_cla30_b), .u_cla30_out(h_u_wallace_cla16_u_cla30_out));

  assign h_u_wallace_cla16_out[0] = h_u_wallace_cla16_and_0_0[0];
  assign h_u_wallace_cla16_out[1] = h_u_wallace_cla16_u_cla30_out[0];
  assign h_u_wallace_cla16_out[2] = h_u_wallace_cla16_u_cla30_out[1];
  assign h_u_wallace_cla16_out[3] = h_u_wallace_cla16_u_cla30_out[2];
  assign h_u_wallace_cla16_out[4] = h_u_wallace_cla16_u_cla30_out[3];
  assign h_u_wallace_cla16_out[5] = h_u_wallace_cla16_u_cla30_out[4];
  assign h_u_wallace_cla16_out[6] = h_u_wallace_cla16_u_cla30_out[5];
  assign h_u_wallace_cla16_out[7] = h_u_wallace_cla16_u_cla30_out[6];
  assign h_u_wallace_cla16_out[8] = h_u_wallace_cla16_u_cla30_out[7];
  assign h_u_wallace_cla16_out[9] = h_u_wallace_cla16_u_cla30_out[8];
  assign h_u_wallace_cla16_out[10] = h_u_wallace_cla16_u_cla30_out[9];
  assign h_u_wallace_cla16_out[11] = h_u_wallace_cla16_u_cla30_out[10];
  assign h_u_wallace_cla16_out[12] = h_u_wallace_cla16_u_cla30_out[11];
  assign h_u_wallace_cla16_out[13] = h_u_wallace_cla16_u_cla30_out[12];
  assign h_u_wallace_cla16_out[14] = h_u_wallace_cla16_u_cla30_out[13];
  assign h_u_wallace_cla16_out[15] = h_u_wallace_cla16_u_cla30_out[14];
  assign h_u_wallace_cla16_out[16] = h_u_wallace_cla16_u_cla30_out[15];
  assign h_u_wallace_cla16_out[17] = h_u_wallace_cla16_u_cla30_out[16];
  assign h_u_wallace_cla16_out[18] = h_u_wallace_cla16_u_cla30_out[17];
  assign h_u_wallace_cla16_out[19] = h_u_wallace_cla16_u_cla30_out[18];
  assign h_u_wallace_cla16_out[20] = h_u_wallace_cla16_u_cla30_out[19];
  assign h_u_wallace_cla16_out[21] = h_u_wallace_cla16_u_cla30_out[20];
  assign h_u_wallace_cla16_out[22] = h_u_wallace_cla16_u_cla30_out[21];
  assign h_u_wallace_cla16_out[23] = h_u_wallace_cla16_u_cla30_out[22];
  assign h_u_wallace_cla16_out[24] = h_u_wallace_cla16_u_cla30_out[23];
  assign h_u_wallace_cla16_out[25] = h_u_wallace_cla16_u_cla30_out[24];
  assign h_u_wallace_cla16_out[26] = h_u_wallace_cla16_u_cla30_out[25];
  assign h_u_wallace_cla16_out[27] = h_u_wallace_cla16_u_cla30_out[26];
  assign h_u_wallace_cla16_out[28] = h_u_wallace_cla16_u_cla30_out[27];
  assign h_u_wallace_cla16_out[29] = h_u_wallace_cla16_u_cla30_out[28];
  assign h_u_wallace_cla16_out[30] = h_u_wallace_cla16_u_cla30_out[29];
  assign h_u_wallace_cla16_out[31] = h_u_wallace_cla16_u_cla30_out[30];
endmodule