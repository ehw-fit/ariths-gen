module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module nor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a | _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module constant_wire_value_0(input a, input b, output constant_wire_0);
  wire constant_wire_value_0_a;
  wire constant_wire_value_0_b;

  assign constant_wire_value_0_a = a;
  assign constant_wire_value_0_b = b;

  xor_gate xor_gate_constant_wire_value_0_y0(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y0);
  xnor_gate xnor_gate_constant_wire_value_0_y1(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y1);
  nor_gate nor_gate_constant_wire_0(constant_wire_value_0_y0, constant_wire_value_0_y1, constant_wire_0);
endmodule

module pg_logic(input a, input b, output pg_logic_y0, output pg_logic_y1, output pg_logic_y2);
  wire pg_logic_a;
  wire pg_logic_b;

  assign pg_logic_a = a;
  assign pg_logic_b = b;

  or_gate or_gate_pg_logic_y0(pg_logic_a, pg_logic_b, pg_logic_y0);
  and_gate and_gate_pg_logic_y1(pg_logic_a, pg_logic_b, pg_logic_y1);
  xor_gate xor_gate_pg_logic_y2(pg_logic_a, pg_logic_b, pg_logic_y2);
endmodule

module h_u_cla24(input [23:0] a, input [23:0] b, output [24:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire constant_wire_0;
  wire h_u_cla24_pg_logic0_y0;
  wire h_u_cla24_pg_logic0_y1;
  wire h_u_cla24_pg_logic0_y2;
  wire h_u_cla24_xor0_y0;
  wire h_u_cla24_and0_y0;
  wire h_u_cla24_or0_y0;
  wire h_u_cla24_pg_logic1_y0;
  wire h_u_cla24_pg_logic1_y1;
  wire h_u_cla24_pg_logic1_y2;
  wire h_u_cla24_xor1_y0;
  wire h_u_cla24_and1_y0;
  wire h_u_cla24_and2_y0;
  wire h_u_cla24_and3_y0;
  wire h_u_cla24_and4_y0;
  wire h_u_cla24_or1_y0;
  wire h_u_cla24_or2_y0;
  wire h_u_cla24_pg_logic2_y0;
  wire h_u_cla24_pg_logic2_y1;
  wire h_u_cla24_pg_logic2_y2;
  wire h_u_cla24_xor2_y0;
  wire h_u_cla24_and5_y0;
  wire h_u_cla24_and6_y0;
  wire h_u_cla24_and7_y0;
  wire h_u_cla24_and8_y0;
  wire h_u_cla24_and9_y0;
  wire h_u_cla24_and10_y0;
  wire h_u_cla24_and11_y0;
  wire h_u_cla24_and12_y0;
  wire h_u_cla24_and13_y0;
  wire h_u_cla24_or3_y0;
  wire h_u_cla24_or4_y0;
  wire h_u_cla24_or5_y0;
  wire h_u_cla24_pg_logic3_y0;
  wire h_u_cla24_pg_logic3_y1;
  wire h_u_cla24_pg_logic3_y2;
  wire h_u_cla24_xor3_y0;
  wire h_u_cla24_and14_y0;
  wire h_u_cla24_and15_y0;
  wire h_u_cla24_and16_y0;
  wire h_u_cla24_and17_y0;
  wire h_u_cla24_and18_y0;
  wire h_u_cla24_and19_y0;
  wire h_u_cla24_and20_y0;
  wire h_u_cla24_and21_y0;
  wire h_u_cla24_and22_y0;
  wire h_u_cla24_and23_y0;
  wire h_u_cla24_and24_y0;
  wire h_u_cla24_and25_y0;
  wire h_u_cla24_and26_y0;
  wire h_u_cla24_and27_y0;
  wire h_u_cla24_and28_y0;
  wire h_u_cla24_and29_y0;
  wire h_u_cla24_or6_y0;
  wire h_u_cla24_or7_y0;
  wire h_u_cla24_or8_y0;
  wire h_u_cla24_or9_y0;
  wire h_u_cla24_pg_logic4_y0;
  wire h_u_cla24_pg_logic4_y1;
  wire h_u_cla24_pg_logic4_y2;
  wire h_u_cla24_xor4_y0;
  wire h_u_cla24_and30_y0;
  wire h_u_cla24_and31_y0;
  wire h_u_cla24_and32_y0;
  wire h_u_cla24_and33_y0;
  wire h_u_cla24_and34_y0;
  wire h_u_cla24_and35_y0;
  wire h_u_cla24_and36_y0;
  wire h_u_cla24_and37_y0;
  wire h_u_cla24_and38_y0;
  wire h_u_cla24_and39_y0;
  wire h_u_cla24_and40_y0;
  wire h_u_cla24_and41_y0;
  wire h_u_cla24_and42_y0;
  wire h_u_cla24_and43_y0;
  wire h_u_cla24_and44_y0;
  wire h_u_cla24_and45_y0;
  wire h_u_cla24_and46_y0;
  wire h_u_cla24_and47_y0;
  wire h_u_cla24_and48_y0;
  wire h_u_cla24_and49_y0;
  wire h_u_cla24_and50_y0;
  wire h_u_cla24_and51_y0;
  wire h_u_cla24_and52_y0;
  wire h_u_cla24_and53_y0;
  wire h_u_cla24_and54_y0;
  wire h_u_cla24_or10_y0;
  wire h_u_cla24_or11_y0;
  wire h_u_cla24_or12_y0;
  wire h_u_cla24_or13_y0;
  wire h_u_cla24_or14_y0;
  wire h_u_cla24_pg_logic5_y0;
  wire h_u_cla24_pg_logic5_y1;
  wire h_u_cla24_pg_logic5_y2;
  wire h_u_cla24_xor5_y0;
  wire h_u_cla24_and55_y0;
  wire h_u_cla24_and56_y0;
  wire h_u_cla24_and57_y0;
  wire h_u_cla24_and58_y0;
  wire h_u_cla24_and59_y0;
  wire h_u_cla24_and60_y0;
  wire h_u_cla24_and61_y0;
  wire h_u_cla24_and62_y0;
  wire h_u_cla24_and63_y0;
  wire h_u_cla24_and64_y0;
  wire h_u_cla24_and65_y0;
  wire h_u_cla24_and66_y0;
  wire h_u_cla24_and67_y0;
  wire h_u_cla24_and68_y0;
  wire h_u_cla24_and69_y0;
  wire h_u_cla24_and70_y0;
  wire h_u_cla24_and71_y0;
  wire h_u_cla24_and72_y0;
  wire h_u_cla24_and73_y0;
  wire h_u_cla24_and74_y0;
  wire h_u_cla24_and75_y0;
  wire h_u_cla24_and76_y0;
  wire h_u_cla24_and77_y0;
  wire h_u_cla24_and78_y0;
  wire h_u_cla24_and79_y0;
  wire h_u_cla24_and80_y0;
  wire h_u_cla24_and81_y0;
  wire h_u_cla24_and82_y0;
  wire h_u_cla24_and83_y0;
  wire h_u_cla24_and84_y0;
  wire h_u_cla24_and85_y0;
  wire h_u_cla24_and86_y0;
  wire h_u_cla24_and87_y0;
  wire h_u_cla24_and88_y0;
  wire h_u_cla24_and89_y0;
  wire h_u_cla24_and90_y0;
  wire h_u_cla24_or15_y0;
  wire h_u_cla24_or16_y0;
  wire h_u_cla24_or17_y0;
  wire h_u_cla24_or18_y0;
  wire h_u_cla24_or19_y0;
  wire h_u_cla24_or20_y0;
  wire h_u_cla24_pg_logic6_y0;
  wire h_u_cla24_pg_logic6_y1;
  wire h_u_cla24_pg_logic6_y2;
  wire h_u_cla24_xor6_y0;
  wire h_u_cla24_and91_y0;
  wire h_u_cla24_and92_y0;
  wire h_u_cla24_and93_y0;
  wire h_u_cla24_and94_y0;
  wire h_u_cla24_and95_y0;
  wire h_u_cla24_and96_y0;
  wire h_u_cla24_and97_y0;
  wire h_u_cla24_and98_y0;
  wire h_u_cla24_and99_y0;
  wire h_u_cla24_and100_y0;
  wire h_u_cla24_and101_y0;
  wire h_u_cla24_and102_y0;
  wire h_u_cla24_and103_y0;
  wire h_u_cla24_and104_y0;
  wire h_u_cla24_and105_y0;
  wire h_u_cla24_and106_y0;
  wire h_u_cla24_and107_y0;
  wire h_u_cla24_and108_y0;
  wire h_u_cla24_and109_y0;
  wire h_u_cla24_and110_y0;
  wire h_u_cla24_and111_y0;
  wire h_u_cla24_and112_y0;
  wire h_u_cla24_and113_y0;
  wire h_u_cla24_and114_y0;
  wire h_u_cla24_and115_y0;
  wire h_u_cla24_and116_y0;
  wire h_u_cla24_and117_y0;
  wire h_u_cla24_and118_y0;
  wire h_u_cla24_and119_y0;
  wire h_u_cla24_and120_y0;
  wire h_u_cla24_and121_y0;
  wire h_u_cla24_and122_y0;
  wire h_u_cla24_and123_y0;
  wire h_u_cla24_and124_y0;
  wire h_u_cla24_and125_y0;
  wire h_u_cla24_and126_y0;
  wire h_u_cla24_and127_y0;
  wire h_u_cla24_and128_y0;
  wire h_u_cla24_and129_y0;
  wire h_u_cla24_and130_y0;
  wire h_u_cla24_and131_y0;
  wire h_u_cla24_and132_y0;
  wire h_u_cla24_and133_y0;
  wire h_u_cla24_and134_y0;
  wire h_u_cla24_and135_y0;
  wire h_u_cla24_and136_y0;
  wire h_u_cla24_and137_y0;
  wire h_u_cla24_and138_y0;
  wire h_u_cla24_and139_y0;
  wire h_u_cla24_or21_y0;
  wire h_u_cla24_or22_y0;
  wire h_u_cla24_or23_y0;
  wire h_u_cla24_or24_y0;
  wire h_u_cla24_or25_y0;
  wire h_u_cla24_or26_y0;
  wire h_u_cla24_or27_y0;
  wire h_u_cla24_pg_logic7_y0;
  wire h_u_cla24_pg_logic7_y1;
  wire h_u_cla24_pg_logic7_y2;
  wire h_u_cla24_xor7_y0;
  wire h_u_cla24_and140_y0;
  wire h_u_cla24_and141_y0;
  wire h_u_cla24_and142_y0;
  wire h_u_cla24_and143_y0;
  wire h_u_cla24_and144_y0;
  wire h_u_cla24_and145_y0;
  wire h_u_cla24_and146_y0;
  wire h_u_cla24_and147_y0;
  wire h_u_cla24_and148_y0;
  wire h_u_cla24_and149_y0;
  wire h_u_cla24_and150_y0;
  wire h_u_cla24_and151_y0;
  wire h_u_cla24_and152_y0;
  wire h_u_cla24_and153_y0;
  wire h_u_cla24_and154_y0;
  wire h_u_cla24_and155_y0;
  wire h_u_cla24_and156_y0;
  wire h_u_cla24_and157_y0;
  wire h_u_cla24_and158_y0;
  wire h_u_cla24_and159_y0;
  wire h_u_cla24_and160_y0;
  wire h_u_cla24_and161_y0;
  wire h_u_cla24_and162_y0;
  wire h_u_cla24_and163_y0;
  wire h_u_cla24_and164_y0;
  wire h_u_cla24_and165_y0;
  wire h_u_cla24_and166_y0;
  wire h_u_cla24_and167_y0;
  wire h_u_cla24_and168_y0;
  wire h_u_cla24_and169_y0;
  wire h_u_cla24_and170_y0;
  wire h_u_cla24_and171_y0;
  wire h_u_cla24_and172_y0;
  wire h_u_cla24_and173_y0;
  wire h_u_cla24_and174_y0;
  wire h_u_cla24_and175_y0;
  wire h_u_cla24_and176_y0;
  wire h_u_cla24_and177_y0;
  wire h_u_cla24_and178_y0;
  wire h_u_cla24_and179_y0;
  wire h_u_cla24_and180_y0;
  wire h_u_cla24_and181_y0;
  wire h_u_cla24_and182_y0;
  wire h_u_cla24_and183_y0;
  wire h_u_cla24_and184_y0;
  wire h_u_cla24_and185_y0;
  wire h_u_cla24_and186_y0;
  wire h_u_cla24_and187_y0;
  wire h_u_cla24_and188_y0;
  wire h_u_cla24_and189_y0;
  wire h_u_cla24_and190_y0;
  wire h_u_cla24_and191_y0;
  wire h_u_cla24_and192_y0;
  wire h_u_cla24_and193_y0;
  wire h_u_cla24_and194_y0;
  wire h_u_cla24_and195_y0;
  wire h_u_cla24_and196_y0;
  wire h_u_cla24_and197_y0;
  wire h_u_cla24_and198_y0;
  wire h_u_cla24_and199_y0;
  wire h_u_cla24_and200_y0;
  wire h_u_cla24_and201_y0;
  wire h_u_cla24_and202_y0;
  wire h_u_cla24_and203_y0;
  wire h_u_cla24_or28_y0;
  wire h_u_cla24_or29_y0;
  wire h_u_cla24_or30_y0;
  wire h_u_cla24_or31_y0;
  wire h_u_cla24_or32_y0;
  wire h_u_cla24_or33_y0;
  wire h_u_cla24_or34_y0;
  wire h_u_cla24_or35_y0;
  wire h_u_cla24_pg_logic8_y0;
  wire h_u_cla24_pg_logic8_y1;
  wire h_u_cla24_pg_logic8_y2;
  wire h_u_cla24_xor8_y0;
  wire h_u_cla24_and204_y0;
  wire h_u_cla24_and205_y0;
  wire h_u_cla24_and206_y0;
  wire h_u_cla24_and207_y0;
  wire h_u_cla24_and208_y0;
  wire h_u_cla24_and209_y0;
  wire h_u_cla24_and210_y0;
  wire h_u_cla24_and211_y0;
  wire h_u_cla24_and212_y0;
  wire h_u_cla24_and213_y0;
  wire h_u_cla24_and214_y0;
  wire h_u_cla24_and215_y0;
  wire h_u_cla24_and216_y0;
  wire h_u_cla24_and217_y0;
  wire h_u_cla24_and218_y0;
  wire h_u_cla24_and219_y0;
  wire h_u_cla24_and220_y0;
  wire h_u_cla24_and221_y0;
  wire h_u_cla24_and222_y0;
  wire h_u_cla24_and223_y0;
  wire h_u_cla24_and224_y0;
  wire h_u_cla24_and225_y0;
  wire h_u_cla24_and226_y0;
  wire h_u_cla24_and227_y0;
  wire h_u_cla24_and228_y0;
  wire h_u_cla24_and229_y0;
  wire h_u_cla24_and230_y0;
  wire h_u_cla24_and231_y0;
  wire h_u_cla24_and232_y0;
  wire h_u_cla24_and233_y0;
  wire h_u_cla24_and234_y0;
  wire h_u_cla24_and235_y0;
  wire h_u_cla24_and236_y0;
  wire h_u_cla24_and237_y0;
  wire h_u_cla24_and238_y0;
  wire h_u_cla24_and239_y0;
  wire h_u_cla24_and240_y0;
  wire h_u_cla24_and241_y0;
  wire h_u_cla24_and242_y0;
  wire h_u_cla24_and243_y0;
  wire h_u_cla24_and244_y0;
  wire h_u_cla24_and245_y0;
  wire h_u_cla24_and246_y0;
  wire h_u_cla24_and247_y0;
  wire h_u_cla24_and248_y0;
  wire h_u_cla24_and249_y0;
  wire h_u_cla24_and250_y0;
  wire h_u_cla24_and251_y0;
  wire h_u_cla24_and252_y0;
  wire h_u_cla24_and253_y0;
  wire h_u_cla24_and254_y0;
  wire h_u_cla24_and255_y0;
  wire h_u_cla24_and256_y0;
  wire h_u_cla24_and257_y0;
  wire h_u_cla24_and258_y0;
  wire h_u_cla24_and259_y0;
  wire h_u_cla24_and260_y0;
  wire h_u_cla24_and261_y0;
  wire h_u_cla24_and262_y0;
  wire h_u_cla24_and263_y0;
  wire h_u_cla24_and264_y0;
  wire h_u_cla24_and265_y0;
  wire h_u_cla24_and266_y0;
  wire h_u_cla24_and267_y0;
  wire h_u_cla24_and268_y0;
  wire h_u_cla24_and269_y0;
  wire h_u_cla24_and270_y0;
  wire h_u_cla24_and271_y0;
  wire h_u_cla24_and272_y0;
  wire h_u_cla24_and273_y0;
  wire h_u_cla24_and274_y0;
  wire h_u_cla24_and275_y0;
  wire h_u_cla24_and276_y0;
  wire h_u_cla24_and277_y0;
  wire h_u_cla24_and278_y0;
  wire h_u_cla24_and279_y0;
  wire h_u_cla24_and280_y0;
  wire h_u_cla24_and281_y0;
  wire h_u_cla24_and282_y0;
  wire h_u_cla24_and283_y0;
  wire h_u_cla24_and284_y0;
  wire h_u_cla24_or36_y0;
  wire h_u_cla24_or37_y0;
  wire h_u_cla24_or38_y0;
  wire h_u_cla24_or39_y0;
  wire h_u_cla24_or40_y0;
  wire h_u_cla24_or41_y0;
  wire h_u_cla24_or42_y0;
  wire h_u_cla24_or43_y0;
  wire h_u_cla24_or44_y0;
  wire h_u_cla24_pg_logic9_y0;
  wire h_u_cla24_pg_logic9_y1;
  wire h_u_cla24_pg_logic9_y2;
  wire h_u_cla24_xor9_y0;
  wire h_u_cla24_and285_y0;
  wire h_u_cla24_and286_y0;
  wire h_u_cla24_and287_y0;
  wire h_u_cla24_and288_y0;
  wire h_u_cla24_and289_y0;
  wire h_u_cla24_and290_y0;
  wire h_u_cla24_and291_y0;
  wire h_u_cla24_and292_y0;
  wire h_u_cla24_and293_y0;
  wire h_u_cla24_and294_y0;
  wire h_u_cla24_and295_y0;
  wire h_u_cla24_and296_y0;
  wire h_u_cla24_and297_y0;
  wire h_u_cla24_and298_y0;
  wire h_u_cla24_and299_y0;
  wire h_u_cla24_and300_y0;
  wire h_u_cla24_and301_y0;
  wire h_u_cla24_and302_y0;
  wire h_u_cla24_and303_y0;
  wire h_u_cla24_and304_y0;
  wire h_u_cla24_and305_y0;
  wire h_u_cla24_and306_y0;
  wire h_u_cla24_and307_y0;
  wire h_u_cla24_and308_y0;
  wire h_u_cla24_and309_y0;
  wire h_u_cla24_and310_y0;
  wire h_u_cla24_and311_y0;
  wire h_u_cla24_and312_y0;
  wire h_u_cla24_and313_y0;
  wire h_u_cla24_and314_y0;
  wire h_u_cla24_and315_y0;
  wire h_u_cla24_and316_y0;
  wire h_u_cla24_and317_y0;
  wire h_u_cla24_and318_y0;
  wire h_u_cla24_and319_y0;
  wire h_u_cla24_and320_y0;
  wire h_u_cla24_and321_y0;
  wire h_u_cla24_and322_y0;
  wire h_u_cla24_and323_y0;
  wire h_u_cla24_and324_y0;
  wire h_u_cla24_and325_y0;
  wire h_u_cla24_and326_y0;
  wire h_u_cla24_and327_y0;
  wire h_u_cla24_and328_y0;
  wire h_u_cla24_and329_y0;
  wire h_u_cla24_and330_y0;
  wire h_u_cla24_and331_y0;
  wire h_u_cla24_and332_y0;
  wire h_u_cla24_and333_y0;
  wire h_u_cla24_and334_y0;
  wire h_u_cla24_and335_y0;
  wire h_u_cla24_and336_y0;
  wire h_u_cla24_and337_y0;
  wire h_u_cla24_and338_y0;
  wire h_u_cla24_and339_y0;
  wire h_u_cla24_and340_y0;
  wire h_u_cla24_and341_y0;
  wire h_u_cla24_and342_y0;
  wire h_u_cla24_and343_y0;
  wire h_u_cla24_and344_y0;
  wire h_u_cla24_and345_y0;
  wire h_u_cla24_and346_y0;
  wire h_u_cla24_and347_y0;
  wire h_u_cla24_and348_y0;
  wire h_u_cla24_and349_y0;
  wire h_u_cla24_and350_y0;
  wire h_u_cla24_and351_y0;
  wire h_u_cla24_and352_y0;
  wire h_u_cla24_and353_y0;
  wire h_u_cla24_and354_y0;
  wire h_u_cla24_and355_y0;
  wire h_u_cla24_and356_y0;
  wire h_u_cla24_and357_y0;
  wire h_u_cla24_and358_y0;
  wire h_u_cla24_and359_y0;
  wire h_u_cla24_and360_y0;
  wire h_u_cla24_and361_y0;
  wire h_u_cla24_and362_y0;
  wire h_u_cla24_and363_y0;
  wire h_u_cla24_and364_y0;
  wire h_u_cla24_and365_y0;
  wire h_u_cla24_and366_y0;
  wire h_u_cla24_and367_y0;
  wire h_u_cla24_and368_y0;
  wire h_u_cla24_and369_y0;
  wire h_u_cla24_and370_y0;
  wire h_u_cla24_and371_y0;
  wire h_u_cla24_and372_y0;
  wire h_u_cla24_and373_y0;
  wire h_u_cla24_and374_y0;
  wire h_u_cla24_and375_y0;
  wire h_u_cla24_and376_y0;
  wire h_u_cla24_and377_y0;
  wire h_u_cla24_and378_y0;
  wire h_u_cla24_and379_y0;
  wire h_u_cla24_and380_y0;
  wire h_u_cla24_and381_y0;
  wire h_u_cla24_and382_y0;
  wire h_u_cla24_and383_y0;
  wire h_u_cla24_and384_y0;
  wire h_u_cla24_or45_y0;
  wire h_u_cla24_or46_y0;
  wire h_u_cla24_or47_y0;
  wire h_u_cla24_or48_y0;
  wire h_u_cla24_or49_y0;
  wire h_u_cla24_or50_y0;
  wire h_u_cla24_or51_y0;
  wire h_u_cla24_or52_y0;
  wire h_u_cla24_or53_y0;
  wire h_u_cla24_or54_y0;
  wire h_u_cla24_pg_logic10_y0;
  wire h_u_cla24_pg_logic10_y1;
  wire h_u_cla24_pg_logic10_y2;
  wire h_u_cla24_xor10_y0;
  wire h_u_cla24_and385_y0;
  wire h_u_cla24_and386_y0;
  wire h_u_cla24_and387_y0;
  wire h_u_cla24_and388_y0;
  wire h_u_cla24_and389_y0;
  wire h_u_cla24_and390_y0;
  wire h_u_cla24_and391_y0;
  wire h_u_cla24_and392_y0;
  wire h_u_cla24_and393_y0;
  wire h_u_cla24_and394_y0;
  wire h_u_cla24_and395_y0;
  wire h_u_cla24_and396_y0;
  wire h_u_cla24_and397_y0;
  wire h_u_cla24_and398_y0;
  wire h_u_cla24_and399_y0;
  wire h_u_cla24_and400_y0;
  wire h_u_cla24_and401_y0;
  wire h_u_cla24_and402_y0;
  wire h_u_cla24_and403_y0;
  wire h_u_cla24_and404_y0;
  wire h_u_cla24_and405_y0;
  wire h_u_cla24_and406_y0;
  wire h_u_cla24_and407_y0;
  wire h_u_cla24_and408_y0;
  wire h_u_cla24_and409_y0;
  wire h_u_cla24_and410_y0;
  wire h_u_cla24_and411_y0;
  wire h_u_cla24_and412_y0;
  wire h_u_cla24_and413_y0;
  wire h_u_cla24_and414_y0;
  wire h_u_cla24_and415_y0;
  wire h_u_cla24_and416_y0;
  wire h_u_cla24_and417_y0;
  wire h_u_cla24_and418_y0;
  wire h_u_cla24_and419_y0;
  wire h_u_cla24_and420_y0;
  wire h_u_cla24_and421_y0;
  wire h_u_cla24_and422_y0;
  wire h_u_cla24_and423_y0;
  wire h_u_cla24_and424_y0;
  wire h_u_cla24_and425_y0;
  wire h_u_cla24_and426_y0;
  wire h_u_cla24_and427_y0;
  wire h_u_cla24_and428_y0;
  wire h_u_cla24_and429_y0;
  wire h_u_cla24_and430_y0;
  wire h_u_cla24_and431_y0;
  wire h_u_cla24_and432_y0;
  wire h_u_cla24_and433_y0;
  wire h_u_cla24_and434_y0;
  wire h_u_cla24_and435_y0;
  wire h_u_cla24_and436_y0;
  wire h_u_cla24_and437_y0;
  wire h_u_cla24_and438_y0;
  wire h_u_cla24_and439_y0;
  wire h_u_cla24_and440_y0;
  wire h_u_cla24_and441_y0;
  wire h_u_cla24_and442_y0;
  wire h_u_cla24_and443_y0;
  wire h_u_cla24_and444_y0;
  wire h_u_cla24_and445_y0;
  wire h_u_cla24_and446_y0;
  wire h_u_cla24_and447_y0;
  wire h_u_cla24_and448_y0;
  wire h_u_cla24_and449_y0;
  wire h_u_cla24_and450_y0;
  wire h_u_cla24_and451_y0;
  wire h_u_cla24_and452_y0;
  wire h_u_cla24_and453_y0;
  wire h_u_cla24_and454_y0;
  wire h_u_cla24_and455_y0;
  wire h_u_cla24_and456_y0;
  wire h_u_cla24_and457_y0;
  wire h_u_cla24_and458_y0;
  wire h_u_cla24_and459_y0;
  wire h_u_cla24_and460_y0;
  wire h_u_cla24_and461_y0;
  wire h_u_cla24_and462_y0;
  wire h_u_cla24_and463_y0;
  wire h_u_cla24_and464_y0;
  wire h_u_cla24_and465_y0;
  wire h_u_cla24_and466_y0;
  wire h_u_cla24_and467_y0;
  wire h_u_cla24_and468_y0;
  wire h_u_cla24_and469_y0;
  wire h_u_cla24_and470_y0;
  wire h_u_cla24_and471_y0;
  wire h_u_cla24_and472_y0;
  wire h_u_cla24_and473_y0;
  wire h_u_cla24_and474_y0;
  wire h_u_cla24_and475_y0;
  wire h_u_cla24_and476_y0;
  wire h_u_cla24_and477_y0;
  wire h_u_cla24_and478_y0;
  wire h_u_cla24_and479_y0;
  wire h_u_cla24_and480_y0;
  wire h_u_cla24_and481_y0;
  wire h_u_cla24_and482_y0;
  wire h_u_cla24_and483_y0;
  wire h_u_cla24_and484_y0;
  wire h_u_cla24_and485_y0;
  wire h_u_cla24_and486_y0;
  wire h_u_cla24_and487_y0;
  wire h_u_cla24_and488_y0;
  wire h_u_cla24_and489_y0;
  wire h_u_cla24_and490_y0;
  wire h_u_cla24_and491_y0;
  wire h_u_cla24_and492_y0;
  wire h_u_cla24_and493_y0;
  wire h_u_cla24_and494_y0;
  wire h_u_cla24_and495_y0;
  wire h_u_cla24_and496_y0;
  wire h_u_cla24_and497_y0;
  wire h_u_cla24_and498_y0;
  wire h_u_cla24_and499_y0;
  wire h_u_cla24_and500_y0;
  wire h_u_cla24_and501_y0;
  wire h_u_cla24_and502_y0;
  wire h_u_cla24_and503_y0;
  wire h_u_cla24_and504_y0;
  wire h_u_cla24_and505_y0;
  wire h_u_cla24_or55_y0;
  wire h_u_cla24_or56_y0;
  wire h_u_cla24_or57_y0;
  wire h_u_cla24_or58_y0;
  wire h_u_cla24_or59_y0;
  wire h_u_cla24_or60_y0;
  wire h_u_cla24_or61_y0;
  wire h_u_cla24_or62_y0;
  wire h_u_cla24_or63_y0;
  wire h_u_cla24_or64_y0;
  wire h_u_cla24_or65_y0;
  wire h_u_cla24_pg_logic11_y0;
  wire h_u_cla24_pg_logic11_y1;
  wire h_u_cla24_pg_logic11_y2;
  wire h_u_cla24_xor11_y0;
  wire h_u_cla24_and506_y0;
  wire h_u_cla24_and507_y0;
  wire h_u_cla24_and508_y0;
  wire h_u_cla24_and509_y0;
  wire h_u_cla24_and510_y0;
  wire h_u_cla24_and511_y0;
  wire h_u_cla24_and512_y0;
  wire h_u_cla24_and513_y0;
  wire h_u_cla24_and514_y0;
  wire h_u_cla24_and515_y0;
  wire h_u_cla24_and516_y0;
  wire h_u_cla24_and517_y0;
  wire h_u_cla24_and518_y0;
  wire h_u_cla24_and519_y0;
  wire h_u_cla24_and520_y0;
  wire h_u_cla24_and521_y0;
  wire h_u_cla24_and522_y0;
  wire h_u_cla24_and523_y0;
  wire h_u_cla24_and524_y0;
  wire h_u_cla24_and525_y0;
  wire h_u_cla24_and526_y0;
  wire h_u_cla24_and527_y0;
  wire h_u_cla24_and528_y0;
  wire h_u_cla24_and529_y0;
  wire h_u_cla24_and530_y0;
  wire h_u_cla24_and531_y0;
  wire h_u_cla24_and532_y0;
  wire h_u_cla24_and533_y0;
  wire h_u_cla24_and534_y0;
  wire h_u_cla24_and535_y0;
  wire h_u_cla24_and536_y0;
  wire h_u_cla24_and537_y0;
  wire h_u_cla24_and538_y0;
  wire h_u_cla24_and539_y0;
  wire h_u_cla24_and540_y0;
  wire h_u_cla24_and541_y0;
  wire h_u_cla24_and542_y0;
  wire h_u_cla24_and543_y0;
  wire h_u_cla24_and544_y0;
  wire h_u_cla24_and545_y0;
  wire h_u_cla24_and546_y0;
  wire h_u_cla24_and547_y0;
  wire h_u_cla24_and548_y0;
  wire h_u_cla24_and549_y0;
  wire h_u_cla24_and550_y0;
  wire h_u_cla24_and551_y0;
  wire h_u_cla24_and552_y0;
  wire h_u_cla24_and553_y0;
  wire h_u_cla24_and554_y0;
  wire h_u_cla24_and555_y0;
  wire h_u_cla24_and556_y0;
  wire h_u_cla24_and557_y0;
  wire h_u_cla24_and558_y0;
  wire h_u_cla24_and559_y0;
  wire h_u_cla24_and560_y0;
  wire h_u_cla24_and561_y0;
  wire h_u_cla24_and562_y0;
  wire h_u_cla24_and563_y0;
  wire h_u_cla24_and564_y0;
  wire h_u_cla24_and565_y0;
  wire h_u_cla24_and566_y0;
  wire h_u_cla24_and567_y0;
  wire h_u_cla24_and568_y0;
  wire h_u_cla24_and569_y0;
  wire h_u_cla24_and570_y0;
  wire h_u_cla24_and571_y0;
  wire h_u_cla24_and572_y0;
  wire h_u_cla24_and573_y0;
  wire h_u_cla24_and574_y0;
  wire h_u_cla24_and575_y0;
  wire h_u_cla24_and576_y0;
  wire h_u_cla24_and577_y0;
  wire h_u_cla24_and578_y0;
  wire h_u_cla24_and579_y0;
  wire h_u_cla24_and580_y0;
  wire h_u_cla24_and581_y0;
  wire h_u_cla24_and582_y0;
  wire h_u_cla24_and583_y0;
  wire h_u_cla24_and584_y0;
  wire h_u_cla24_and585_y0;
  wire h_u_cla24_and586_y0;
  wire h_u_cla24_and587_y0;
  wire h_u_cla24_and588_y0;
  wire h_u_cla24_and589_y0;
  wire h_u_cla24_and590_y0;
  wire h_u_cla24_and591_y0;
  wire h_u_cla24_and592_y0;
  wire h_u_cla24_and593_y0;
  wire h_u_cla24_and594_y0;
  wire h_u_cla24_and595_y0;
  wire h_u_cla24_and596_y0;
  wire h_u_cla24_and597_y0;
  wire h_u_cla24_and598_y0;
  wire h_u_cla24_and599_y0;
  wire h_u_cla24_and600_y0;
  wire h_u_cla24_and601_y0;
  wire h_u_cla24_and602_y0;
  wire h_u_cla24_and603_y0;
  wire h_u_cla24_and604_y0;
  wire h_u_cla24_and605_y0;
  wire h_u_cla24_and606_y0;
  wire h_u_cla24_and607_y0;
  wire h_u_cla24_and608_y0;
  wire h_u_cla24_and609_y0;
  wire h_u_cla24_and610_y0;
  wire h_u_cla24_and611_y0;
  wire h_u_cla24_and612_y0;
  wire h_u_cla24_and613_y0;
  wire h_u_cla24_and614_y0;
  wire h_u_cla24_and615_y0;
  wire h_u_cla24_and616_y0;
  wire h_u_cla24_and617_y0;
  wire h_u_cla24_and618_y0;
  wire h_u_cla24_and619_y0;
  wire h_u_cla24_and620_y0;
  wire h_u_cla24_and621_y0;
  wire h_u_cla24_and622_y0;
  wire h_u_cla24_and623_y0;
  wire h_u_cla24_and624_y0;
  wire h_u_cla24_and625_y0;
  wire h_u_cla24_and626_y0;
  wire h_u_cla24_and627_y0;
  wire h_u_cla24_and628_y0;
  wire h_u_cla24_and629_y0;
  wire h_u_cla24_and630_y0;
  wire h_u_cla24_and631_y0;
  wire h_u_cla24_and632_y0;
  wire h_u_cla24_and633_y0;
  wire h_u_cla24_and634_y0;
  wire h_u_cla24_and635_y0;
  wire h_u_cla24_and636_y0;
  wire h_u_cla24_and637_y0;
  wire h_u_cla24_and638_y0;
  wire h_u_cla24_and639_y0;
  wire h_u_cla24_and640_y0;
  wire h_u_cla24_and641_y0;
  wire h_u_cla24_and642_y0;
  wire h_u_cla24_and643_y0;
  wire h_u_cla24_and644_y0;
  wire h_u_cla24_and645_y0;
  wire h_u_cla24_and646_y0;
  wire h_u_cla24_and647_y0;
  wire h_u_cla24_and648_y0;
  wire h_u_cla24_and649_y0;
  wire h_u_cla24_or66_y0;
  wire h_u_cla24_or67_y0;
  wire h_u_cla24_or68_y0;
  wire h_u_cla24_or69_y0;
  wire h_u_cla24_or70_y0;
  wire h_u_cla24_or71_y0;
  wire h_u_cla24_or72_y0;
  wire h_u_cla24_or73_y0;
  wire h_u_cla24_or74_y0;
  wire h_u_cla24_or75_y0;
  wire h_u_cla24_or76_y0;
  wire h_u_cla24_or77_y0;
  wire h_u_cla24_pg_logic12_y0;
  wire h_u_cla24_pg_logic12_y1;
  wire h_u_cla24_pg_logic12_y2;
  wire h_u_cla24_xor12_y0;
  wire h_u_cla24_and650_y0;
  wire h_u_cla24_and651_y0;
  wire h_u_cla24_and652_y0;
  wire h_u_cla24_and653_y0;
  wire h_u_cla24_and654_y0;
  wire h_u_cla24_and655_y0;
  wire h_u_cla24_and656_y0;
  wire h_u_cla24_and657_y0;
  wire h_u_cla24_and658_y0;
  wire h_u_cla24_and659_y0;
  wire h_u_cla24_and660_y0;
  wire h_u_cla24_and661_y0;
  wire h_u_cla24_and662_y0;
  wire h_u_cla24_and663_y0;
  wire h_u_cla24_and664_y0;
  wire h_u_cla24_and665_y0;
  wire h_u_cla24_and666_y0;
  wire h_u_cla24_and667_y0;
  wire h_u_cla24_and668_y0;
  wire h_u_cla24_and669_y0;
  wire h_u_cla24_and670_y0;
  wire h_u_cla24_and671_y0;
  wire h_u_cla24_and672_y0;
  wire h_u_cla24_and673_y0;
  wire h_u_cla24_and674_y0;
  wire h_u_cla24_and675_y0;
  wire h_u_cla24_and676_y0;
  wire h_u_cla24_and677_y0;
  wire h_u_cla24_and678_y0;
  wire h_u_cla24_and679_y0;
  wire h_u_cla24_and680_y0;
  wire h_u_cla24_and681_y0;
  wire h_u_cla24_and682_y0;
  wire h_u_cla24_and683_y0;
  wire h_u_cla24_and684_y0;
  wire h_u_cla24_and685_y0;
  wire h_u_cla24_and686_y0;
  wire h_u_cla24_and687_y0;
  wire h_u_cla24_and688_y0;
  wire h_u_cla24_and689_y0;
  wire h_u_cla24_and690_y0;
  wire h_u_cla24_and691_y0;
  wire h_u_cla24_and692_y0;
  wire h_u_cla24_and693_y0;
  wire h_u_cla24_and694_y0;
  wire h_u_cla24_and695_y0;
  wire h_u_cla24_and696_y0;
  wire h_u_cla24_and697_y0;
  wire h_u_cla24_and698_y0;
  wire h_u_cla24_and699_y0;
  wire h_u_cla24_and700_y0;
  wire h_u_cla24_and701_y0;
  wire h_u_cla24_and702_y0;
  wire h_u_cla24_and703_y0;
  wire h_u_cla24_and704_y0;
  wire h_u_cla24_and705_y0;
  wire h_u_cla24_and706_y0;
  wire h_u_cla24_and707_y0;
  wire h_u_cla24_and708_y0;
  wire h_u_cla24_and709_y0;
  wire h_u_cla24_and710_y0;
  wire h_u_cla24_and711_y0;
  wire h_u_cla24_and712_y0;
  wire h_u_cla24_and713_y0;
  wire h_u_cla24_and714_y0;
  wire h_u_cla24_and715_y0;
  wire h_u_cla24_and716_y0;
  wire h_u_cla24_and717_y0;
  wire h_u_cla24_and718_y0;
  wire h_u_cla24_and719_y0;
  wire h_u_cla24_and720_y0;
  wire h_u_cla24_and721_y0;
  wire h_u_cla24_and722_y0;
  wire h_u_cla24_and723_y0;
  wire h_u_cla24_and724_y0;
  wire h_u_cla24_and725_y0;
  wire h_u_cla24_and726_y0;
  wire h_u_cla24_and727_y0;
  wire h_u_cla24_and728_y0;
  wire h_u_cla24_and729_y0;
  wire h_u_cla24_and730_y0;
  wire h_u_cla24_and731_y0;
  wire h_u_cla24_and732_y0;
  wire h_u_cla24_and733_y0;
  wire h_u_cla24_and734_y0;
  wire h_u_cla24_and735_y0;
  wire h_u_cla24_and736_y0;
  wire h_u_cla24_and737_y0;
  wire h_u_cla24_and738_y0;
  wire h_u_cla24_and739_y0;
  wire h_u_cla24_and740_y0;
  wire h_u_cla24_and741_y0;
  wire h_u_cla24_and742_y0;
  wire h_u_cla24_and743_y0;
  wire h_u_cla24_and744_y0;
  wire h_u_cla24_and745_y0;
  wire h_u_cla24_and746_y0;
  wire h_u_cla24_and747_y0;
  wire h_u_cla24_and748_y0;
  wire h_u_cla24_and749_y0;
  wire h_u_cla24_and750_y0;
  wire h_u_cla24_and751_y0;
  wire h_u_cla24_and752_y0;
  wire h_u_cla24_and753_y0;
  wire h_u_cla24_and754_y0;
  wire h_u_cla24_and755_y0;
  wire h_u_cla24_and756_y0;
  wire h_u_cla24_and757_y0;
  wire h_u_cla24_and758_y0;
  wire h_u_cla24_and759_y0;
  wire h_u_cla24_and760_y0;
  wire h_u_cla24_and761_y0;
  wire h_u_cla24_and762_y0;
  wire h_u_cla24_and763_y0;
  wire h_u_cla24_and764_y0;
  wire h_u_cla24_and765_y0;
  wire h_u_cla24_and766_y0;
  wire h_u_cla24_and767_y0;
  wire h_u_cla24_and768_y0;
  wire h_u_cla24_and769_y0;
  wire h_u_cla24_and770_y0;
  wire h_u_cla24_and771_y0;
  wire h_u_cla24_and772_y0;
  wire h_u_cla24_and773_y0;
  wire h_u_cla24_and774_y0;
  wire h_u_cla24_and775_y0;
  wire h_u_cla24_and776_y0;
  wire h_u_cla24_and777_y0;
  wire h_u_cla24_and778_y0;
  wire h_u_cla24_and779_y0;
  wire h_u_cla24_and780_y0;
  wire h_u_cla24_and781_y0;
  wire h_u_cla24_and782_y0;
  wire h_u_cla24_and783_y0;
  wire h_u_cla24_and784_y0;
  wire h_u_cla24_and785_y0;
  wire h_u_cla24_and786_y0;
  wire h_u_cla24_and787_y0;
  wire h_u_cla24_and788_y0;
  wire h_u_cla24_and789_y0;
  wire h_u_cla24_and790_y0;
  wire h_u_cla24_and791_y0;
  wire h_u_cla24_and792_y0;
  wire h_u_cla24_and793_y0;
  wire h_u_cla24_and794_y0;
  wire h_u_cla24_and795_y0;
  wire h_u_cla24_and796_y0;
  wire h_u_cla24_and797_y0;
  wire h_u_cla24_and798_y0;
  wire h_u_cla24_and799_y0;
  wire h_u_cla24_and800_y0;
  wire h_u_cla24_and801_y0;
  wire h_u_cla24_and802_y0;
  wire h_u_cla24_and803_y0;
  wire h_u_cla24_and804_y0;
  wire h_u_cla24_and805_y0;
  wire h_u_cla24_and806_y0;
  wire h_u_cla24_and807_y0;
  wire h_u_cla24_and808_y0;
  wire h_u_cla24_and809_y0;
  wire h_u_cla24_and810_y0;
  wire h_u_cla24_and811_y0;
  wire h_u_cla24_and812_y0;
  wire h_u_cla24_and813_y0;
  wire h_u_cla24_and814_y0;
  wire h_u_cla24_and815_y0;
  wire h_u_cla24_and816_y0;
  wire h_u_cla24_and817_y0;
  wire h_u_cla24_and818_y0;
  wire h_u_cla24_or78_y0;
  wire h_u_cla24_or79_y0;
  wire h_u_cla24_or80_y0;
  wire h_u_cla24_or81_y0;
  wire h_u_cla24_or82_y0;
  wire h_u_cla24_or83_y0;
  wire h_u_cla24_or84_y0;
  wire h_u_cla24_or85_y0;
  wire h_u_cla24_or86_y0;
  wire h_u_cla24_or87_y0;
  wire h_u_cla24_or88_y0;
  wire h_u_cla24_or89_y0;
  wire h_u_cla24_or90_y0;
  wire h_u_cla24_pg_logic13_y0;
  wire h_u_cla24_pg_logic13_y1;
  wire h_u_cla24_pg_logic13_y2;
  wire h_u_cla24_xor13_y0;
  wire h_u_cla24_and819_y0;
  wire h_u_cla24_and820_y0;
  wire h_u_cla24_and821_y0;
  wire h_u_cla24_and822_y0;
  wire h_u_cla24_and823_y0;
  wire h_u_cla24_and824_y0;
  wire h_u_cla24_and825_y0;
  wire h_u_cla24_and826_y0;
  wire h_u_cla24_and827_y0;
  wire h_u_cla24_and828_y0;
  wire h_u_cla24_and829_y0;
  wire h_u_cla24_and830_y0;
  wire h_u_cla24_and831_y0;
  wire h_u_cla24_and832_y0;
  wire h_u_cla24_and833_y0;
  wire h_u_cla24_and834_y0;
  wire h_u_cla24_and835_y0;
  wire h_u_cla24_and836_y0;
  wire h_u_cla24_and837_y0;
  wire h_u_cla24_and838_y0;
  wire h_u_cla24_and839_y0;
  wire h_u_cla24_and840_y0;
  wire h_u_cla24_and841_y0;
  wire h_u_cla24_and842_y0;
  wire h_u_cla24_and843_y0;
  wire h_u_cla24_and844_y0;
  wire h_u_cla24_and845_y0;
  wire h_u_cla24_and846_y0;
  wire h_u_cla24_and847_y0;
  wire h_u_cla24_and848_y0;
  wire h_u_cla24_and849_y0;
  wire h_u_cla24_and850_y0;
  wire h_u_cla24_and851_y0;
  wire h_u_cla24_and852_y0;
  wire h_u_cla24_and853_y0;
  wire h_u_cla24_and854_y0;
  wire h_u_cla24_and855_y0;
  wire h_u_cla24_and856_y0;
  wire h_u_cla24_and857_y0;
  wire h_u_cla24_and858_y0;
  wire h_u_cla24_and859_y0;
  wire h_u_cla24_and860_y0;
  wire h_u_cla24_and861_y0;
  wire h_u_cla24_and862_y0;
  wire h_u_cla24_and863_y0;
  wire h_u_cla24_and864_y0;
  wire h_u_cla24_and865_y0;
  wire h_u_cla24_and866_y0;
  wire h_u_cla24_and867_y0;
  wire h_u_cla24_and868_y0;
  wire h_u_cla24_and869_y0;
  wire h_u_cla24_and870_y0;
  wire h_u_cla24_and871_y0;
  wire h_u_cla24_and872_y0;
  wire h_u_cla24_and873_y0;
  wire h_u_cla24_and874_y0;
  wire h_u_cla24_and875_y0;
  wire h_u_cla24_and876_y0;
  wire h_u_cla24_and877_y0;
  wire h_u_cla24_and878_y0;
  wire h_u_cla24_and879_y0;
  wire h_u_cla24_and880_y0;
  wire h_u_cla24_and881_y0;
  wire h_u_cla24_and882_y0;
  wire h_u_cla24_and883_y0;
  wire h_u_cla24_and884_y0;
  wire h_u_cla24_and885_y0;
  wire h_u_cla24_and886_y0;
  wire h_u_cla24_and887_y0;
  wire h_u_cla24_and888_y0;
  wire h_u_cla24_and889_y0;
  wire h_u_cla24_and890_y0;
  wire h_u_cla24_and891_y0;
  wire h_u_cla24_and892_y0;
  wire h_u_cla24_and893_y0;
  wire h_u_cla24_and894_y0;
  wire h_u_cla24_and895_y0;
  wire h_u_cla24_and896_y0;
  wire h_u_cla24_and897_y0;
  wire h_u_cla24_and898_y0;
  wire h_u_cla24_and899_y0;
  wire h_u_cla24_and900_y0;
  wire h_u_cla24_and901_y0;
  wire h_u_cla24_and902_y0;
  wire h_u_cla24_and903_y0;
  wire h_u_cla24_and904_y0;
  wire h_u_cla24_and905_y0;
  wire h_u_cla24_and906_y0;
  wire h_u_cla24_and907_y0;
  wire h_u_cla24_and908_y0;
  wire h_u_cla24_and909_y0;
  wire h_u_cla24_and910_y0;
  wire h_u_cla24_and911_y0;
  wire h_u_cla24_and912_y0;
  wire h_u_cla24_and913_y0;
  wire h_u_cla24_and914_y0;
  wire h_u_cla24_and915_y0;
  wire h_u_cla24_and916_y0;
  wire h_u_cla24_and917_y0;
  wire h_u_cla24_and918_y0;
  wire h_u_cla24_and919_y0;
  wire h_u_cla24_and920_y0;
  wire h_u_cla24_and921_y0;
  wire h_u_cla24_and922_y0;
  wire h_u_cla24_and923_y0;
  wire h_u_cla24_and924_y0;
  wire h_u_cla24_and925_y0;
  wire h_u_cla24_and926_y0;
  wire h_u_cla24_and927_y0;
  wire h_u_cla24_and928_y0;
  wire h_u_cla24_and929_y0;
  wire h_u_cla24_and930_y0;
  wire h_u_cla24_and931_y0;
  wire h_u_cla24_and932_y0;
  wire h_u_cla24_and933_y0;
  wire h_u_cla24_and934_y0;
  wire h_u_cla24_and935_y0;
  wire h_u_cla24_and936_y0;
  wire h_u_cla24_and937_y0;
  wire h_u_cla24_and938_y0;
  wire h_u_cla24_and939_y0;
  wire h_u_cla24_and940_y0;
  wire h_u_cla24_and941_y0;
  wire h_u_cla24_and942_y0;
  wire h_u_cla24_and943_y0;
  wire h_u_cla24_and944_y0;
  wire h_u_cla24_and945_y0;
  wire h_u_cla24_and946_y0;
  wire h_u_cla24_and947_y0;
  wire h_u_cla24_and948_y0;
  wire h_u_cla24_and949_y0;
  wire h_u_cla24_and950_y0;
  wire h_u_cla24_and951_y0;
  wire h_u_cla24_and952_y0;
  wire h_u_cla24_and953_y0;
  wire h_u_cla24_and954_y0;
  wire h_u_cla24_and955_y0;
  wire h_u_cla24_and956_y0;
  wire h_u_cla24_and957_y0;
  wire h_u_cla24_and958_y0;
  wire h_u_cla24_and959_y0;
  wire h_u_cla24_and960_y0;
  wire h_u_cla24_and961_y0;
  wire h_u_cla24_and962_y0;
  wire h_u_cla24_and963_y0;
  wire h_u_cla24_and964_y0;
  wire h_u_cla24_and965_y0;
  wire h_u_cla24_and966_y0;
  wire h_u_cla24_and967_y0;
  wire h_u_cla24_and968_y0;
  wire h_u_cla24_and969_y0;
  wire h_u_cla24_and970_y0;
  wire h_u_cla24_and971_y0;
  wire h_u_cla24_and972_y0;
  wire h_u_cla24_and973_y0;
  wire h_u_cla24_and974_y0;
  wire h_u_cla24_and975_y0;
  wire h_u_cla24_and976_y0;
  wire h_u_cla24_and977_y0;
  wire h_u_cla24_and978_y0;
  wire h_u_cla24_and979_y0;
  wire h_u_cla24_and980_y0;
  wire h_u_cla24_and981_y0;
  wire h_u_cla24_and982_y0;
  wire h_u_cla24_and983_y0;
  wire h_u_cla24_and984_y0;
  wire h_u_cla24_and985_y0;
  wire h_u_cla24_and986_y0;
  wire h_u_cla24_and987_y0;
  wire h_u_cla24_and988_y0;
  wire h_u_cla24_and989_y0;
  wire h_u_cla24_and990_y0;
  wire h_u_cla24_and991_y0;
  wire h_u_cla24_and992_y0;
  wire h_u_cla24_and993_y0;
  wire h_u_cla24_and994_y0;
  wire h_u_cla24_and995_y0;
  wire h_u_cla24_and996_y0;
  wire h_u_cla24_and997_y0;
  wire h_u_cla24_and998_y0;
  wire h_u_cla24_and999_y0;
  wire h_u_cla24_and1000_y0;
  wire h_u_cla24_and1001_y0;
  wire h_u_cla24_and1002_y0;
  wire h_u_cla24_and1003_y0;
  wire h_u_cla24_and1004_y0;
  wire h_u_cla24_and1005_y0;
  wire h_u_cla24_and1006_y0;
  wire h_u_cla24_and1007_y0;
  wire h_u_cla24_and1008_y0;
  wire h_u_cla24_and1009_y0;
  wire h_u_cla24_and1010_y0;
  wire h_u_cla24_and1011_y0;
  wire h_u_cla24_and1012_y0;
  wire h_u_cla24_and1013_y0;
  wire h_u_cla24_and1014_y0;
  wire h_u_cla24_or91_y0;
  wire h_u_cla24_or92_y0;
  wire h_u_cla24_or93_y0;
  wire h_u_cla24_or94_y0;
  wire h_u_cla24_or95_y0;
  wire h_u_cla24_or96_y0;
  wire h_u_cla24_or97_y0;
  wire h_u_cla24_or98_y0;
  wire h_u_cla24_or99_y0;
  wire h_u_cla24_or100_y0;
  wire h_u_cla24_or101_y0;
  wire h_u_cla24_or102_y0;
  wire h_u_cla24_or103_y0;
  wire h_u_cla24_or104_y0;
  wire h_u_cla24_pg_logic14_y0;
  wire h_u_cla24_pg_logic14_y1;
  wire h_u_cla24_pg_logic14_y2;
  wire h_u_cla24_xor14_y0;
  wire h_u_cla24_and1015_y0;
  wire h_u_cla24_and1016_y0;
  wire h_u_cla24_and1017_y0;
  wire h_u_cla24_and1018_y0;
  wire h_u_cla24_and1019_y0;
  wire h_u_cla24_and1020_y0;
  wire h_u_cla24_and1021_y0;
  wire h_u_cla24_and1022_y0;
  wire h_u_cla24_and1023_y0;
  wire h_u_cla24_and1024_y0;
  wire h_u_cla24_and1025_y0;
  wire h_u_cla24_and1026_y0;
  wire h_u_cla24_and1027_y0;
  wire h_u_cla24_and1028_y0;
  wire h_u_cla24_and1029_y0;
  wire h_u_cla24_and1030_y0;
  wire h_u_cla24_and1031_y0;
  wire h_u_cla24_and1032_y0;
  wire h_u_cla24_and1033_y0;
  wire h_u_cla24_and1034_y0;
  wire h_u_cla24_and1035_y0;
  wire h_u_cla24_and1036_y0;
  wire h_u_cla24_and1037_y0;
  wire h_u_cla24_and1038_y0;
  wire h_u_cla24_and1039_y0;
  wire h_u_cla24_and1040_y0;
  wire h_u_cla24_and1041_y0;
  wire h_u_cla24_and1042_y0;
  wire h_u_cla24_and1043_y0;
  wire h_u_cla24_and1044_y0;
  wire h_u_cla24_and1045_y0;
  wire h_u_cla24_and1046_y0;
  wire h_u_cla24_and1047_y0;
  wire h_u_cla24_and1048_y0;
  wire h_u_cla24_and1049_y0;
  wire h_u_cla24_and1050_y0;
  wire h_u_cla24_and1051_y0;
  wire h_u_cla24_and1052_y0;
  wire h_u_cla24_and1053_y0;
  wire h_u_cla24_and1054_y0;
  wire h_u_cla24_and1055_y0;
  wire h_u_cla24_and1056_y0;
  wire h_u_cla24_and1057_y0;
  wire h_u_cla24_and1058_y0;
  wire h_u_cla24_and1059_y0;
  wire h_u_cla24_and1060_y0;
  wire h_u_cla24_and1061_y0;
  wire h_u_cla24_and1062_y0;
  wire h_u_cla24_and1063_y0;
  wire h_u_cla24_and1064_y0;
  wire h_u_cla24_and1065_y0;
  wire h_u_cla24_and1066_y0;
  wire h_u_cla24_and1067_y0;
  wire h_u_cla24_and1068_y0;
  wire h_u_cla24_and1069_y0;
  wire h_u_cla24_and1070_y0;
  wire h_u_cla24_and1071_y0;
  wire h_u_cla24_and1072_y0;
  wire h_u_cla24_and1073_y0;
  wire h_u_cla24_and1074_y0;
  wire h_u_cla24_and1075_y0;
  wire h_u_cla24_and1076_y0;
  wire h_u_cla24_and1077_y0;
  wire h_u_cla24_and1078_y0;
  wire h_u_cla24_and1079_y0;
  wire h_u_cla24_and1080_y0;
  wire h_u_cla24_and1081_y0;
  wire h_u_cla24_and1082_y0;
  wire h_u_cla24_and1083_y0;
  wire h_u_cla24_and1084_y0;
  wire h_u_cla24_and1085_y0;
  wire h_u_cla24_and1086_y0;
  wire h_u_cla24_and1087_y0;
  wire h_u_cla24_and1088_y0;
  wire h_u_cla24_and1089_y0;
  wire h_u_cla24_and1090_y0;
  wire h_u_cla24_and1091_y0;
  wire h_u_cla24_and1092_y0;
  wire h_u_cla24_and1093_y0;
  wire h_u_cla24_and1094_y0;
  wire h_u_cla24_and1095_y0;
  wire h_u_cla24_and1096_y0;
  wire h_u_cla24_and1097_y0;
  wire h_u_cla24_and1098_y0;
  wire h_u_cla24_and1099_y0;
  wire h_u_cla24_and1100_y0;
  wire h_u_cla24_and1101_y0;
  wire h_u_cla24_and1102_y0;
  wire h_u_cla24_and1103_y0;
  wire h_u_cla24_and1104_y0;
  wire h_u_cla24_and1105_y0;
  wire h_u_cla24_and1106_y0;
  wire h_u_cla24_and1107_y0;
  wire h_u_cla24_and1108_y0;
  wire h_u_cla24_and1109_y0;
  wire h_u_cla24_and1110_y0;
  wire h_u_cla24_and1111_y0;
  wire h_u_cla24_and1112_y0;
  wire h_u_cla24_and1113_y0;
  wire h_u_cla24_and1114_y0;
  wire h_u_cla24_and1115_y0;
  wire h_u_cla24_and1116_y0;
  wire h_u_cla24_and1117_y0;
  wire h_u_cla24_and1118_y0;
  wire h_u_cla24_and1119_y0;
  wire h_u_cla24_and1120_y0;
  wire h_u_cla24_and1121_y0;
  wire h_u_cla24_and1122_y0;
  wire h_u_cla24_and1123_y0;
  wire h_u_cla24_and1124_y0;
  wire h_u_cla24_and1125_y0;
  wire h_u_cla24_and1126_y0;
  wire h_u_cla24_and1127_y0;
  wire h_u_cla24_and1128_y0;
  wire h_u_cla24_and1129_y0;
  wire h_u_cla24_and1130_y0;
  wire h_u_cla24_and1131_y0;
  wire h_u_cla24_and1132_y0;
  wire h_u_cla24_and1133_y0;
  wire h_u_cla24_and1134_y0;
  wire h_u_cla24_and1135_y0;
  wire h_u_cla24_and1136_y0;
  wire h_u_cla24_and1137_y0;
  wire h_u_cla24_and1138_y0;
  wire h_u_cla24_and1139_y0;
  wire h_u_cla24_and1140_y0;
  wire h_u_cla24_and1141_y0;
  wire h_u_cla24_and1142_y0;
  wire h_u_cla24_and1143_y0;
  wire h_u_cla24_and1144_y0;
  wire h_u_cla24_and1145_y0;
  wire h_u_cla24_and1146_y0;
  wire h_u_cla24_and1147_y0;
  wire h_u_cla24_and1148_y0;
  wire h_u_cla24_and1149_y0;
  wire h_u_cla24_and1150_y0;
  wire h_u_cla24_and1151_y0;
  wire h_u_cla24_and1152_y0;
  wire h_u_cla24_and1153_y0;
  wire h_u_cla24_and1154_y0;
  wire h_u_cla24_and1155_y0;
  wire h_u_cla24_and1156_y0;
  wire h_u_cla24_and1157_y0;
  wire h_u_cla24_and1158_y0;
  wire h_u_cla24_and1159_y0;
  wire h_u_cla24_and1160_y0;
  wire h_u_cla24_and1161_y0;
  wire h_u_cla24_and1162_y0;
  wire h_u_cla24_and1163_y0;
  wire h_u_cla24_and1164_y0;
  wire h_u_cla24_and1165_y0;
  wire h_u_cla24_and1166_y0;
  wire h_u_cla24_and1167_y0;
  wire h_u_cla24_and1168_y0;
  wire h_u_cla24_and1169_y0;
  wire h_u_cla24_and1170_y0;
  wire h_u_cla24_and1171_y0;
  wire h_u_cla24_and1172_y0;
  wire h_u_cla24_and1173_y0;
  wire h_u_cla24_and1174_y0;
  wire h_u_cla24_and1175_y0;
  wire h_u_cla24_and1176_y0;
  wire h_u_cla24_and1177_y0;
  wire h_u_cla24_and1178_y0;
  wire h_u_cla24_and1179_y0;
  wire h_u_cla24_and1180_y0;
  wire h_u_cla24_and1181_y0;
  wire h_u_cla24_and1182_y0;
  wire h_u_cla24_and1183_y0;
  wire h_u_cla24_and1184_y0;
  wire h_u_cla24_and1185_y0;
  wire h_u_cla24_and1186_y0;
  wire h_u_cla24_and1187_y0;
  wire h_u_cla24_and1188_y0;
  wire h_u_cla24_and1189_y0;
  wire h_u_cla24_and1190_y0;
  wire h_u_cla24_and1191_y0;
  wire h_u_cla24_and1192_y0;
  wire h_u_cla24_and1193_y0;
  wire h_u_cla24_and1194_y0;
  wire h_u_cla24_and1195_y0;
  wire h_u_cla24_and1196_y0;
  wire h_u_cla24_and1197_y0;
  wire h_u_cla24_and1198_y0;
  wire h_u_cla24_and1199_y0;
  wire h_u_cla24_and1200_y0;
  wire h_u_cla24_and1201_y0;
  wire h_u_cla24_and1202_y0;
  wire h_u_cla24_and1203_y0;
  wire h_u_cla24_and1204_y0;
  wire h_u_cla24_and1205_y0;
  wire h_u_cla24_and1206_y0;
  wire h_u_cla24_and1207_y0;
  wire h_u_cla24_and1208_y0;
  wire h_u_cla24_and1209_y0;
  wire h_u_cla24_and1210_y0;
  wire h_u_cla24_and1211_y0;
  wire h_u_cla24_and1212_y0;
  wire h_u_cla24_and1213_y0;
  wire h_u_cla24_and1214_y0;
  wire h_u_cla24_and1215_y0;
  wire h_u_cla24_and1216_y0;
  wire h_u_cla24_and1217_y0;
  wire h_u_cla24_and1218_y0;
  wire h_u_cla24_and1219_y0;
  wire h_u_cla24_and1220_y0;
  wire h_u_cla24_and1221_y0;
  wire h_u_cla24_and1222_y0;
  wire h_u_cla24_and1223_y0;
  wire h_u_cla24_and1224_y0;
  wire h_u_cla24_and1225_y0;
  wire h_u_cla24_and1226_y0;
  wire h_u_cla24_and1227_y0;
  wire h_u_cla24_and1228_y0;
  wire h_u_cla24_and1229_y0;
  wire h_u_cla24_and1230_y0;
  wire h_u_cla24_and1231_y0;
  wire h_u_cla24_and1232_y0;
  wire h_u_cla24_and1233_y0;
  wire h_u_cla24_and1234_y0;
  wire h_u_cla24_and1235_y0;
  wire h_u_cla24_and1236_y0;
  wire h_u_cla24_and1237_y0;
  wire h_u_cla24_and1238_y0;
  wire h_u_cla24_and1239_y0;
  wire h_u_cla24_or105_y0;
  wire h_u_cla24_or106_y0;
  wire h_u_cla24_or107_y0;
  wire h_u_cla24_or108_y0;
  wire h_u_cla24_or109_y0;
  wire h_u_cla24_or110_y0;
  wire h_u_cla24_or111_y0;
  wire h_u_cla24_or112_y0;
  wire h_u_cla24_or113_y0;
  wire h_u_cla24_or114_y0;
  wire h_u_cla24_or115_y0;
  wire h_u_cla24_or116_y0;
  wire h_u_cla24_or117_y0;
  wire h_u_cla24_or118_y0;
  wire h_u_cla24_or119_y0;
  wire h_u_cla24_pg_logic15_y0;
  wire h_u_cla24_pg_logic15_y1;
  wire h_u_cla24_pg_logic15_y2;
  wire h_u_cla24_xor15_y0;
  wire h_u_cla24_and1240_y0;
  wire h_u_cla24_and1241_y0;
  wire h_u_cla24_and1242_y0;
  wire h_u_cla24_and1243_y0;
  wire h_u_cla24_and1244_y0;
  wire h_u_cla24_and1245_y0;
  wire h_u_cla24_and1246_y0;
  wire h_u_cla24_and1247_y0;
  wire h_u_cla24_and1248_y0;
  wire h_u_cla24_and1249_y0;
  wire h_u_cla24_and1250_y0;
  wire h_u_cla24_and1251_y0;
  wire h_u_cla24_and1252_y0;
  wire h_u_cla24_and1253_y0;
  wire h_u_cla24_and1254_y0;
  wire h_u_cla24_and1255_y0;
  wire h_u_cla24_and1256_y0;
  wire h_u_cla24_and1257_y0;
  wire h_u_cla24_and1258_y0;
  wire h_u_cla24_and1259_y0;
  wire h_u_cla24_and1260_y0;
  wire h_u_cla24_and1261_y0;
  wire h_u_cla24_and1262_y0;
  wire h_u_cla24_and1263_y0;
  wire h_u_cla24_and1264_y0;
  wire h_u_cla24_and1265_y0;
  wire h_u_cla24_and1266_y0;
  wire h_u_cla24_and1267_y0;
  wire h_u_cla24_and1268_y0;
  wire h_u_cla24_and1269_y0;
  wire h_u_cla24_and1270_y0;
  wire h_u_cla24_and1271_y0;
  wire h_u_cla24_and1272_y0;
  wire h_u_cla24_and1273_y0;
  wire h_u_cla24_and1274_y0;
  wire h_u_cla24_and1275_y0;
  wire h_u_cla24_and1276_y0;
  wire h_u_cla24_and1277_y0;
  wire h_u_cla24_and1278_y0;
  wire h_u_cla24_and1279_y0;
  wire h_u_cla24_and1280_y0;
  wire h_u_cla24_and1281_y0;
  wire h_u_cla24_and1282_y0;
  wire h_u_cla24_and1283_y0;
  wire h_u_cla24_and1284_y0;
  wire h_u_cla24_and1285_y0;
  wire h_u_cla24_and1286_y0;
  wire h_u_cla24_and1287_y0;
  wire h_u_cla24_and1288_y0;
  wire h_u_cla24_and1289_y0;
  wire h_u_cla24_and1290_y0;
  wire h_u_cla24_and1291_y0;
  wire h_u_cla24_and1292_y0;
  wire h_u_cla24_and1293_y0;
  wire h_u_cla24_and1294_y0;
  wire h_u_cla24_and1295_y0;
  wire h_u_cla24_and1296_y0;
  wire h_u_cla24_and1297_y0;
  wire h_u_cla24_and1298_y0;
  wire h_u_cla24_and1299_y0;
  wire h_u_cla24_and1300_y0;
  wire h_u_cla24_and1301_y0;
  wire h_u_cla24_and1302_y0;
  wire h_u_cla24_and1303_y0;
  wire h_u_cla24_and1304_y0;
  wire h_u_cla24_and1305_y0;
  wire h_u_cla24_and1306_y0;
  wire h_u_cla24_and1307_y0;
  wire h_u_cla24_and1308_y0;
  wire h_u_cla24_and1309_y0;
  wire h_u_cla24_and1310_y0;
  wire h_u_cla24_and1311_y0;
  wire h_u_cla24_and1312_y0;
  wire h_u_cla24_and1313_y0;
  wire h_u_cla24_and1314_y0;
  wire h_u_cla24_and1315_y0;
  wire h_u_cla24_and1316_y0;
  wire h_u_cla24_and1317_y0;
  wire h_u_cla24_and1318_y0;
  wire h_u_cla24_and1319_y0;
  wire h_u_cla24_and1320_y0;
  wire h_u_cla24_and1321_y0;
  wire h_u_cla24_and1322_y0;
  wire h_u_cla24_and1323_y0;
  wire h_u_cla24_and1324_y0;
  wire h_u_cla24_and1325_y0;
  wire h_u_cla24_and1326_y0;
  wire h_u_cla24_and1327_y0;
  wire h_u_cla24_and1328_y0;
  wire h_u_cla24_and1329_y0;
  wire h_u_cla24_and1330_y0;
  wire h_u_cla24_and1331_y0;
  wire h_u_cla24_and1332_y0;
  wire h_u_cla24_and1333_y0;
  wire h_u_cla24_and1334_y0;
  wire h_u_cla24_and1335_y0;
  wire h_u_cla24_and1336_y0;
  wire h_u_cla24_and1337_y0;
  wire h_u_cla24_and1338_y0;
  wire h_u_cla24_and1339_y0;
  wire h_u_cla24_and1340_y0;
  wire h_u_cla24_and1341_y0;
  wire h_u_cla24_and1342_y0;
  wire h_u_cla24_and1343_y0;
  wire h_u_cla24_and1344_y0;
  wire h_u_cla24_and1345_y0;
  wire h_u_cla24_and1346_y0;
  wire h_u_cla24_and1347_y0;
  wire h_u_cla24_and1348_y0;
  wire h_u_cla24_and1349_y0;
  wire h_u_cla24_and1350_y0;
  wire h_u_cla24_and1351_y0;
  wire h_u_cla24_and1352_y0;
  wire h_u_cla24_and1353_y0;
  wire h_u_cla24_and1354_y0;
  wire h_u_cla24_and1355_y0;
  wire h_u_cla24_and1356_y0;
  wire h_u_cla24_and1357_y0;
  wire h_u_cla24_and1358_y0;
  wire h_u_cla24_and1359_y0;
  wire h_u_cla24_and1360_y0;
  wire h_u_cla24_and1361_y0;
  wire h_u_cla24_and1362_y0;
  wire h_u_cla24_and1363_y0;
  wire h_u_cla24_and1364_y0;
  wire h_u_cla24_and1365_y0;
  wire h_u_cla24_and1366_y0;
  wire h_u_cla24_and1367_y0;
  wire h_u_cla24_and1368_y0;
  wire h_u_cla24_and1369_y0;
  wire h_u_cla24_and1370_y0;
  wire h_u_cla24_and1371_y0;
  wire h_u_cla24_and1372_y0;
  wire h_u_cla24_and1373_y0;
  wire h_u_cla24_and1374_y0;
  wire h_u_cla24_and1375_y0;
  wire h_u_cla24_and1376_y0;
  wire h_u_cla24_and1377_y0;
  wire h_u_cla24_and1378_y0;
  wire h_u_cla24_and1379_y0;
  wire h_u_cla24_and1380_y0;
  wire h_u_cla24_and1381_y0;
  wire h_u_cla24_and1382_y0;
  wire h_u_cla24_and1383_y0;
  wire h_u_cla24_and1384_y0;
  wire h_u_cla24_and1385_y0;
  wire h_u_cla24_and1386_y0;
  wire h_u_cla24_and1387_y0;
  wire h_u_cla24_and1388_y0;
  wire h_u_cla24_and1389_y0;
  wire h_u_cla24_and1390_y0;
  wire h_u_cla24_and1391_y0;
  wire h_u_cla24_and1392_y0;
  wire h_u_cla24_and1393_y0;
  wire h_u_cla24_and1394_y0;
  wire h_u_cla24_and1395_y0;
  wire h_u_cla24_and1396_y0;
  wire h_u_cla24_and1397_y0;
  wire h_u_cla24_and1398_y0;
  wire h_u_cla24_and1399_y0;
  wire h_u_cla24_and1400_y0;
  wire h_u_cla24_and1401_y0;
  wire h_u_cla24_and1402_y0;
  wire h_u_cla24_and1403_y0;
  wire h_u_cla24_and1404_y0;
  wire h_u_cla24_and1405_y0;
  wire h_u_cla24_and1406_y0;
  wire h_u_cla24_and1407_y0;
  wire h_u_cla24_and1408_y0;
  wire h_u_cla24_and1409_y0;
  wire h_u_cla24_and1410_y0;
  wire h_u_cla24_and1411_y0;
  wire h_u_cla24_and1412_y0;
  wire h_u_cla24_and1413_y0;
  wire h_u_cla24_and1414_y0;
  wire h_u_cla24_and1415_y0;
  wire h_u_cla24_and1416_y0;
  wire h_u_cla24_and1417_y0;
  wire h_u_cla24_and1418_y0;
  wire h_u_cla24_and1419_y0;
  wire h_u_cla24_and1420_y0;
  wire h_u_cla24_and1421_y0;
  wire h_u_cla24_and1422_y0;
  wire h_u_cla24_and1423_y0;
  wire h_u_cla24_and1424_y0;
  wire h_u_cla24_and1425_y0;
  wire h_u_cla24_and1426_y0;
  wire h_u_cla24_and1427_y0;
  wire h_u_cla24_and1428_y0;
  wire h_u_cla24_and1429_y0;
  wire h_u_cla24_and1430_y0;
  wire h_u_cla24_and1431_y0;
  wire h_u_cla24_and1432_y0;
  wire h_u_cla24_and1433_y0;
  wire h_u_cla24_and1434_y0;
  wire h_u_cla24_and1435_y0;
  wire h_u_cla24_and1436_y0;
  wire h_u_cla24_and1437_y0;
  wire h_u_cla24_and1438_y0;
  wire h_u_cla24_and1439_y0;
  wire h_u_cla24_and1440_y0;
  wire h_u_cla24_and1441_y0;
  wire h_u_cla24_and1442_y0;
  wire h_u_cla24_and1443_y0;
  wire h_u_cla24_and1444_y0;
  wire h_u_cla24_and1445_y0;
  wire h_u_cla24_and1446_y0;
  wire h_u_cla24_and1447_y0;
  wire h_u_cla24_and1448_y0;
  wire h_u_cla24_and1449_y0;
  wire h_u_cla24_and1450_y0;
  wire h_u_cla24_and1451_y0;
  wire h_u_cla24_and1452_y0;
  wire h_u_cla24_and1453_y0;
  wire h_u_cla24_and1454_y0;
  wire h_u_cla24_and1455_y0;
  wire h_u_cla24_and1456_y0;
  wire h_u_cla24_and1457_y0;
  wire h_u_cla24_and1458_y0;
  wire h_u_cla24_and1459_y0;
  wire h_u_cla24_and1460_y0;
  wire h_u_cla24_and1461_y0;
  wire h_u_cla24_and1462_y0;
  wire h_u_cla24_and1463_y0;
  wire h_u_cla24_and1464_y0;
  wire h_u_cla24_and1465_y0;
  wire h_u_cla24_and1466_y0;
  wire h_u_cla24_and1467_y0;
  wire h_u_cla24_and1468_y0;
  wire h_u_cla24_and1469_y0;
  wire h_u_cla24_and1470_y0;
  wire h_u_cla24_and1471_y0;
  wire h_u_cla24_and1472_y0;
  wire h_u_cla24_and1473_y0;
  wire h_u_cla24_and1474_y0;
  wire h_u_cla24_and1475_y0;
  wire h_u_cla24_and1476_y0;
  wire h_u_cla24_and1477_y0;
  wire h_u_cla24_and1478_y0;
  wire h_u_cla24_and1479_y0;
  wire h_u_cla24_and1480_y0;
  wire h_u_cla24_and1481_y0;
  wire h_u_cla24_and1482_y0;
  wire h_u_cla24_and1483_y0;
  wire h_u_cla24_and1484_y0;
  wire h_u_cla24_and1485_y0;
  wire h_u_cla24_and1486_y0;
  wire h_u_cla24_and1487_y0;
  wire h_u_cla24_and1488_y0;
  wire h_u_cla24_and1489_y0;
  wire h_u_cla24_and1490_y0;
  wire h_u_cla24_and1491_y0;
  wire h_u_cla24_and1492_y0;
  wire h_u_cla24_and1493_y0;
  wire h_u_cla24_and1494_y0;
  wire h_u_cla24_and1495_y0;
  wire h_u_cla24_or120_y0;
  wire h_u_cla24_or121_y0;
  wire h_u_cla24_or122_y0;
  wire h_u_cla24_or123_y0;
  wire h_u_cla24_or124_y0;
  wire h_u_cla24_or125_y0;
  wire h_u_cla24_or126_y0;
  wire h_u_cla24_or127_y0;
  wire h_u_cla24_or128_y0;
  wire h_u_cla24_or129_y0;
  wire h_u_cla24_or130_y0;
  wire h_u_cla24_or131_y0;
  wire h_u_cla24_or132_y0;
  wire h_u_cla24_or133_y0;
  wire h_u_cla24_or134_y0;
  wire h_u_cla24_or135_y0;
  wire h_u_cla24_pg_logic16_y0;
  wire h_u_cla24_pg_logic16_y1;
  wire h_u_cla24_pg_logic16_y2;
  wire h_u_cla24_xor16_y0;
  wire h_u_cla24_and1496_y0;
  wire h_u_cla24_and1497_y0;
  wire h_u_cla24_and1498_y0;
  wire h_u_cla24_and1499_y0;
  wire h_u_cla24_and1500_y0;
  wire h_u_cla24_and1501_y0;
  wire h_u_cla24_and1502_y0;
  wire h_u_cla24_and1503_y0;
  wire h_u_cla24_and1504_y0;
  wire h_u_cla24_and1505_y0;
  wire h_u_cla24_and1506_y0;
  wire h_u_cla24_and1507_y0;
  wire h_u_cla24_and1508_y0;
  wire h_u_cla24_and1509_y0;
  wire h_u_cla24_and1510_y0;
  wire h_u_cla24_and1511_y0;
  wire h_u_cla24_and1512_y0;
  wire h_u_cla24_and1513_y0;
  wire h_u_cla24_and1514_y0;
  wire h_u_cla24_and1515_y0;
  wire h_u_cla24_and1516_y0;
  wire h_u_cla24_and1517_y0;
  wire h_u_cla24_and1518_y0;
  wire h_u_cla24_and1519_y0;
  wire h_u_cla24_and1520_y0;
  wire h_u_cla24_and1521_y0;
  wire h_u_cla24_and1522_y0;
  wire h_u_cla24_and1523_y0;
  wire h_u_cla24_and1524_y0;
  wire h_u_cla24_and1525_y0;
  wire h_u_cla24_and1526_y0;
  wire h_u_cla24_and1527_y0;
  wire h_u_cla24_and1528_y0;
  wire h_u_cla24_and1529_y0;
  wire h_u_cla24_and1530_y0;
  wire h_u_cla24_and1531_y0;
  wire h_u_cla24_and1532_y0;
  wire h_u_cla24_and1533_y0;
  wire h_u_cla24_and1534_y0;
  wire h_u_cla24_and1535_y0;
  wire h_u_cla24_and1536_y0;
  wire h_u_cla24_and1537_y0;
  wire h_u_cla24_and1538_y0;
  wire h_u_cla24_and1539_y0;
  wire h_u_cla24_and1540_y0;
  wire h_u_cla24_and1541_y0;
  wire h_u_cla24_and1542_y0;
  wire h_u_cla24_and1543_y0;
  wire h_u_cla24_and1544_y0;
  wire h_u_cla24_and1545_y0;
  wire h_u_cla24_and1546_y0;
  wire h_u_cla24_and1547_y0;
  wire h_u_cla24_and1548_y0;
  wire h_u_cla24_and1549_y0;
  wire h_u_cla24_and1550_y0;
  wire h_u_cla24_and1551_y0;
  wire h_u_cla24_and1552_y0;
  wire h_u_cla24_and1553_y0;
  wire h_u_cla24_and1554_y0;
  wire h_u_cla24_and1555_y0;
  wire h_u_cla24_and1556_y0;
  wire h_u_cla24_and1557_y0;
  wire h_u_cla24_and1558_y0;
  wire h_u_cla24_and1559_y0;
  wire h_u_cla24_and1560_y0;
  wire h_u_cla24_and1561_y0;
  wire h_u_cla24_and1562_y0;
  wire h_u_cla24_and1563_y0;
  wire h_u_cla24_and1564_y0;
  wire h_u_cla24_and1565_y0;
  wire h_u_cla24_and1566_y0;
  wire h_u_cla24_and1567_y0;
  wire h_u_cla24_and1568_y0;
  wire h_u_cla24_and1569_y0;
  wire h_u_cla24_and1570_y0;
  wire h_u_cla24_and1571_y0;
  wire h_u_cla24_and1572_y0;
  wire h_u_cla24_and1573_y0;
  wire h_u_cla24_and1574_y0;
  wire h_u_cla24_and1575_y0;
  wire h_u_cla24_and1576_y0;
  wire h_u_cla24_and1577_y0;
  wire h_u_cla24_and1578_y0;
  wire h_u_cla24_and1579_y0;
  wire h_u_cla24_and1580_y0;
  wire h_u_cla24_and1581_y0;
  wire h_u_cla24_and1582_y0;
  wire h_u_cla24_and1583_y0;
  wire h_u_cla24_and1584_y0;
  wire h_u_cla24_and1585_y0;
  wire h_u_cla24_and1586_y0;
  wire h_u_cla24_and1587_y0;
  wire h_u_cla24_and1588_y0;
  wire h_u_cla24_and1589_y0;
  wire h_u_cla24_and1590_y0;
  wire h_u_cla24_and1591_y0;
  wire h_u_cla24_and1592_y0;
  wire h_u_cla24_and1593_y0;
  wire h_u_cla24_and1594_y0;
  wire h_u_cla24_and1595_y0;
  wire h_u_cla24_and1596_y0;
  wire h_u_cla24_and1597_y0;
  wire h_u_cla24_and1598_y0;
  wire h_u_cla24_and1599_y0;
  wire h_u_cla24_and1600_y0;
  wire h_u_cla24_and1601_y0;
  wire h_u_cla24_and1602_y0;
  wire h_u_cla24_and1603_y0;
  wire h_u_cla24_and1604_y0;
  wire h_u_cla24_and1605_y0;
  wire h_u_cla24_and1606_y0;
  wire h_u_cla24_and1607_y0;
  wire h_u_cla24_and1608_y0;
  wire h_u_cla24_and1609_y0;
  wire h_u_cla24_and1610_y0;
  wire h_u_cla24_and1611_y0;
  wire h_u_cla24_and1612_y0;
  wire h_u_cla24_and1613_y0;
  wire h_u_cla24_and1614_y0;
  wire h_u_cla24_and1615_y0;
  wire h_u_cla24_and1616_y0;
  wire h_u_cla24_and1617_y0;
  wire h_u_cla24_and1618_y0;
  wire h_u_cla24_and1619_y0;
  wire h_u_cla24_and1620_y0;
  wire h_u_cla24_and1621_y0;
  wire h_u_cla24_and1622_y0;
  wire h_u_cla24_and1623_y0;
  wire h_u_cla24_and1624_y0;
  wire h_u_cla24_and1625_y0;
  wire h_u_cla24_and1626_y0;
  wire h_u_cla24_and1627_y0;
  wire h_u_cla24_and1628_y0;
  wire h_u_cla24_and1629_y0;
  wire h_u_cla24_and1630_y0;
  wire h_u_cla24_and1631_y0;
  wire h_u_cla24_and1632_y0;
  wire h_u_cla24_and1633_y0;
  wire h_u_cla24_and1634_y0;
  wire h_u_cla24_and1635_y0;
  wire h_u_cla24_and1636_y0;
  wire h_u_cla24_and1637_y0;
  wire h_u_cla24_and1638_y0;
  wire h_u_cla24_and1639_y0;
  wire h_u_cla24_and1640_y0;
  wire h_u_cla24_and1641_y0;
  wire h_u_cla24_and1642_y0;
  wire h_u_cla24_and1643_y0;
  wire h_u_cla24_and1644_y0;
  wire h_u_cla24_and1645_y0;
  wire h_u_cla24_and1646_y0;
  wire h_u_cla24_and1647_y0;
  wire h_u_cla24_and1648_y0;
  wire h_u_cla24_and1649_y0;
  wire h_u_cla24_and1650_y0;
  wire h_u_cla24_and1651_y0;
  wire h_u_cla24_and1652_y0;
  wire h_u_cla24_and1653_y0;
  wire h_u_cla24_and1654_y0;
  wire h_u_cla24_and1655_y0;
  wire h_u_cla24_and1656_y0;
  wire h_u_cla24_and1657_y0;
  wire h_u_cla24_and1658_y0;
  wire h_u_cla24_and1659_y0;
  wire h_u_cla24_and1660_y0;
  wire h_u_cla24_and1661_y0;
  wire h_u_cla24_and1662_y0;
  wire h_u_cla24_and1663_y0;
  wire h_u_cla24_and1664_y0;
  wire h_u_cla24_and1665_y0;
  wire h_u_cla24_and1666_y0;
  wire h_u_cla24_and1667_y0;
  wire h_u_cla24_and1668_y0;
  wire h_u_cla24_and1669_y0;
  wire h_u_cla24_and1670_y0;
  wire h_u_cla24_and1671_y0;
  wire h_u_cla24_and1672_y0;
  wire h_u_cla24_and1673_y0;
  wire h_u_cla24_and1674_y0;
  wire h_u_cla24_and1675_y0;
  wire h_u_cla24_and1676_y0;
  wire h_u_cla24_and1677_y0;
  wire h_u_cla24_and1678_y0;
  wire h_u_cla24_and1679_y0;
  wire h_u_cla24_and1680_y0;
  wire h_u_cla24_and1681_y0;
  wire h_u_cla24_and1682_y0;
  wire h_u_cla24_and1683_y0;
  wire h_u_cla24_and1684_y0;
  wire h_u_cla24_and1685_y0;
  wire h_u_cla24_and1686_y0;
  wire h_u_cla24_and1687_y0;
  wire h_u_cla24_and1688_y0;
  wire h_u_cla24_and1689_y0;
  wire h_u_cla24_and1690_y0;
  wire h_u_cla24_and1691_y0;
  wire h_u_cla24_and1692_y0;
  wire h_u_cla24_and1693_y0;
  wire h_u_cla24_and1694_y0;
  wire h_u_cla24_and1695_y0;
  wire h_u_cla24_and1696_y0;
  wire h_u_cla24_and1697_y0;
  wire h_u_cla24_and1698_y0;
  wire h_u_cla24_and1699_y0;
  wire h_u_cla24_and1700_y0;
  wire h_u_cla24_and1701_y0;
  wire h_u_cla24_and1702_y0;
  wire h_u_cla24_and1703_y0;
  wire h_u_cla24_and1704_y0;
  wire h_u_cla24_and1705_y0;
  wire h_u_cla24_and1706_y0;
  wire h_u_cla24_and1707_y0;
  wire h_u_cla24_and1708_y0;
  wire h_u_cla24_and1709_y0;
  wire h_u_cla24_and1710_y0;
  wire h_u_cla24_and1711_y0;
  wire h_u_cla24_and1712_y0;
  wire h_u_cla24_and1713_y0;
  wire h_u_cla24_and1714_y0;
  wire h_u_cla24_and1715_y0;
  wire h_u_cla24_and1716_y0;
  wire h_u_cla24_and1717_y0;
  wire h_u_cla24_and1718_y0;
  wire h_u_cla24_and1719_y0;
  wire h_u_cla24_and1720_y0;
  wire h_u_cla24_and1721_y0;
  wire h_u_cla24_and1722_y0;
  wire h_u_cla24_and1723_y0;
  wire h_u_cla24_and1724_y0;
  wire h_u_cla24_and1725_y0;
  wire h_u_cla24_and1726_y0;
  wire h_u_cla24_and1727_y0;
  wire h_u_cla24_and1728_y0;
  wire h_u_cla24_and1729_y0;
  wire h_u_cla24_and1730_y0;
  wire h_u_cla24_and1731_y0;
  wire h_u_cla24_and1732_y0;
  wire h_u_cla24_and1733_y0;
  wire h_u_cla24_and1734_y0;
  wire h_u_cla24_and1735_y0;
  wire h_u_cla24_and1736_y0;
  wire h_u_cla24_and1737_y0;
  wire h_u_cla24_and1738_y0;
  wire h_u_cla24_and1739_y0;
  wire h_u_cla24_and1740_y0;
  wire h_u_cla24_and1741_y0;
  wire h_u_cla24_and1742_y0;
  wire h_u_cla24_and1743_y0;
  wire h_u_cla24_and1744_y0;
  wire h_u_cla24_and1745_y0;
  wire h_u_cla24_and1746_y0;
  wire h_u_cla24_and1747_y0;
  wire h_u_cla24_and1748_y0;
  wire h_u_cla24_and1749_y0;
  wire h_u_cla24_and1750_y0;
  wire h_u_cla24_and1751_y0;
  wire h_u_cla24_and1752_y0;
  wire h_u_cla24_and1753_y0;
  wire h_u_cla24_and1754_y0;
  wire h_u_cla24_and1755_y0;
  wire h_u_cla24_and1756_y0;
  wire h_u_cla24_and1757_y0;
  wire h_u_cla24_and1758_y0;
  wire h_u_cla24_and1759_y0;
  wire h_u_cla24_and1760_y0;
  wire h_u_cla24_and1761_y0;
  wire h_u_cla24_and1762_y0;
  wire h_u_cla24_and1763_y0;
  wire h_u_cla24_and1764_y0;
  wire h_u_cla24_and1765_y0;
  wire h_u_cla24_and1766_y0;
  wire h_u_cla24_and1767_y0;
  wire h_u_cla24_and1768_y0;
  wire h_u_cla24_and1769_y0;
  wire h_u_cla24_and1770_y0;
  wire h_u_cla24_and1771_y0;
  wire h_u_cla24_and1772_y0;
  wire h_u_cla24_and1773_y0;
  wire h_u_cla24_and1774_y0;
  wire h_u_cla24_and1775_y0;
  wire h_u_cla24_and1776_y0;
  wire h_u_cla24_and1777_y0;
  wire h_u_cla24_and1778_y0;
  wire h_u_cla24_and1779_y0;
  wire h_u_cla24_and1780_y0;
  wire h_u_cla24_and1781_y0;
  wire h_u_cla24_and1782_y0;
  wire h_u_cla24_and1783_y0;
  wire h_u_cla24_and1784_y0;
  wire h_u_cla24_or136_y0;
  wire h_u_cla24_or137_y0;
  wire h_u_cla24_or138_y0;
  wire h_u_cla24_or139_y0;
  wire h_u_cla24_or140_y0;
  wire h_u_cla24_or141_y0;
  wire h_u_cla24_or142_y0;
  wire h_u_cla24_or143_y0;
  wire h_u_cla24_or144_y0;
  wire h_u_cla24_or145_y0;
  wire h_u_cla24_or146_y0;
  wire h_u_cla24_or147_y0;
  wire h_u_cla24_or148_y0;
  wire h_u_cla24_or149_y0;
  wire h_u_cla24_or150_y0;
  wire h_u_cla24_or151_y0;
  wire h_u_cla24_or152_y0;
  wire h_u_cla24_pg_logic17_y0;
  wire h_u_cla24_pg_logic17_y1;
  wire h_u_cla24_pg_logic17_y2;
  wire h_u_cla24_xor17_y0;
  wire h_u_cla24_and1785_y0;
  wire h_u_cla24_and1786_y0;
  wire h_u_cla24_and1787_y0;
  wire h_u_cla24_and1788_y0;
  wire h_u_cla24_and1789_y0;
  wire h_u_cla24_and1790_y0;
  wire h_u_cla24_and1791_y0;
  wire h_u_cla24_and1792_y0;
  wire h_u_cla24_and1793_y0;
  wire h_u_cla24_and1794_y0;
  wire h_u_cla24_and1795_y0;
  wire h_u_cla24_and1796_y0;
  wire h_u_cla24_and1797_y0;
  wire h_u_cla24_and1798_y0;
  wire h_u_cla24_and1799_y0;
  wire h_u_cla24_and1800_y0;
  wire h_u_cla24_and1801_y0;
  wire h_u_cla24_and1802_y0;
  wire h_u_cla24_and1803_y0;
  wire h_u_cla24_and1804_y0;
  wire h_u_cla24_and1805_y0;
  wire h_u_cla24_and1806_y0;
  wire h_u_cla24_and1807_y0;
  wire h_u_cla24_and1808_y0;
  wire h_u_cla24_and1809_y0;
  wire h_u_cla24_and1810_y0;
  wire h_u_cla24_and1811_y0;
  wire h_u_cla24_and1812_y0;
  wire h_u_cla24_and1813_y0;
  wire h_u_cla24_and1814_y0;
  wire h_u_cla24_and1815_y0;
  wire h_u_cla24_and1816_y0;
  wire h_u_cla24_and1817_y0;
  wire h_u_cla24_and1818_y0;
  wire h_u_cla24_and1819_y0;
  wire h_u_cla24_and1820_y0;
  wire h_u_cla24_and1821_y0;
  wire h_u_cla24_and1822_y0;
  wire h_u_cla24_and1823_y0;
  wire h_u_cla24_and1824_y0;
  wire h_u_cla24_and1825_y0;
  wire h_u_cla24_and1826_y0;
  wire h_u_cla24_and1827_y0;
  wire h_u_cla24_and1828_y0;
  wire h_u_cla24_and1829_y0;
  wire h_u_cla24_and1830_y0;
  wire h_u_cla24_and1831_y0;
  wire h_u_cla24_and1832_y0;
  wire h_u_cla24_and1833_y0;
  wire h_u_cla24_and1834_y0;
  wire h_u_cla24_and1835_y0;
  wire h_u_cla24_and1836_y0;
  wire h_u_cla24_and1837_y0;
  wire h_u_cla24_and1838_y0;
  wire h_u_cla24_and1839_y0;
  wire h_u_cla24_and1840_y0;
  wire h_u_cla24_and1841_y0;
  wire h_u_cla24_and1842_y0;
  wire h_u_cla24_and1843_y0;
  wire h_u_cla24_and1844_y0;
  wire h_u_cla24_and1845_y0;
  wire h_u_cla24_and1846_y0;
  wire h_u_cla24_and1847_y0;
  wire h_u_cla24_and1848_y0;
  wire h_u_cla24_and1849_y0;
  wire h_u_cla24_and1850_y0;
  wire h_u_cla24_and1851_y0;
  wire h_u_cla24_and1852_y0;
  wire h_u_cla24_and1853_y0;
  wire h_u_cla24_and1854_y0;
  wire h_u_cla24_and1855_y0;
  wire h_u_cla24_and1856_y0;
  wire h_u_cla24_and1857_y0;
  wire h_u_cla24_and1858_y0;
  wire h_u_cla24_and1859_y0;
  wire h_u_cla24_and1860_y0;
  wire h_u_cla24_and1861_y0;
  wire h_u_cla24_and1862_y0;
  wire h_u_cla24_and1863_y0;
  wire h_u_cla24_and1864_y0;
  wire h_u_cla24_and1865_y0;
  wire h_u_cla24_and1866_y0;
  wire h_u_cla24_and1867_y0;
  wire h_u_cla24_and1868_y0;
  wire h_u_cla24_and1869_y0;
  wire h_u_cla24_and1870_y0;
  wire h_u_cla24_and1871_y0;
  wire h_u_cla24_and1872_y0;
  wire h_u_cla24_and1873_y0;
  wire h_u_cla24_and1874_y0;
  wire h_u_cla24_and1875_y0;
  wire h_u_cla24_and1876_y0;
  wire h_u_cla24_and1877_y0;
  wire h_u_cla24_and1878_y0;
  wire h_u_cla24_and1879_y0;
  wire h_u_cla24_and1880_y0;
  wire h_u_cla24_and1881_y0;
  wire h_u_cla24_and1882_y0;
  wire h_u_cla24_and1883_y0;
  wire h_u_cla24_and1884_y0;
  wire h_u_cla24_and1885_y0;
  wire h_u_cla24_and1886_y0;
  wire h_u_cla24_and1887_y0;
  wire h_u_cla24_and1888_y0;
  wire h_u_cla24_and1889_y0;
  wire h_u_cla24_and1890_y0;
  wire h_u_cla24_and1891_y0;
  wire h_u_cla24_and1892_y0;
  wire h_u_cla24_and1893_y0;
  wire h_u_cla24_and1894_y0;
  wire h_u_cla24_and1895_y0;
  wire h_u_cla24_and1896_y0;
  wire h_u_cla24_and1897_y0;
  wire h_u_cla24_and1898_y0;
  wire h_u_cla24_and1899_y0;
  wire h_u_cla24_and1900_y0;
  wire h_u_cla24_and1901_y0;
  wire h_u_cla24_and1902_y0;
  wire h_u_cla24_and1903_y0;
  wire h_u_cla24_and1904_y0;
  wire h_u_cla24_and1905_y0;
  wire h_u_cla24_and1906_y0;
  wire h_u_cla24_and1907_y0;
  wire h_u_cla24_and1908_y0;
  wire h_u_cla24_and1909_y0;
  wire h_u_cla24_and1910_y0;
  wire h_u_cla24_and1911_y0;
  wire h_u_cla24_and1912_y0;
  wire h_u_cla24_and1913_y0;
  wire h_u_cla24_and1914_y0;
  wire h_u_cla24_and1915_y0;
  wire h_u_cla24_and1916_y0;
  wire h_u_cla24_and1917_y0;
  wire h_u_cla24_and1918_y0;
  wire h_u_cla24_and1919_y0;
  wire h_u_cla24_and1920_y0;
  wire h_u_cla24_and1921_y0;
  wire h_u_cla24_and1922_y0;
  wire h_u_cla24_and1923_y0;
  wire h_u_cla24_and1924_y0;
  wire h_u_cla24_and1925_y0;
  wire h_u_cla24_and1926_y0;
  wire h_u_cla24_and1927_y0;
  wire h_u_cla24_and1928_y0;
  wire h_u_cla24_and1929_y0;
  wire h_u_cla24_and1930_y0;
  wire h_u_cla24_and1931_y0;
  wire h_u_cla24_and1932_y0;
  wire h_u_cla24_and1933_y0;
  wire h_u_cla24_and1934_y0;
  wire h_u_cla24_and1935_y0;
  wire h_u_cla24_and1936_y0;
  wire h_u_cla24_and1937_y0;
  wire h_u_cla24_and1938_y0;
  wire h_u_cla24_and1939_y0;
  wire h_u_cla24_and1940_y0;
  wire h_u_cla24_and1941_y0;
  wire h_u_cla24_and1942_y0;
  wire h_u_cla24_and1943_y0;
  wire h_u_cla24_and1944_y0;
  wire h_u_cla24_and1945_y0;
  wire h_u_cla24_and1946_y0;
  wire h_u_cla24_and1947_y0;
  wire h_u_cla24_and1948_y0;
  wire h_u_cla24_and1949_y0;
  wire h_u_cla24_and1950_y0;
  wire h_u_cla24_and1951_y0;
  wire h_u_cla24_and1952_y0;
  wire h_u_cla24_and1953_y0;
  wire h_u_cla24_and1954_y0;
  wire h_u_cla24_and1955_y0;
  wire h_u_cla24_and1956_y0;
  wire h_u_cla24_and1957_y0;
  wire h_u_cla24_and1958_y0;
  wire h_u_cla24_and1959_y0;
  wire h_u_cla24_and1960_y0;
  wire h_u_cla24_and1961_y0;
  wire h_u_cla24_and1962_y0;
  wire h_u_cla24_and1963_y0;
  wire h_u_cla24_and1964_y0;
  wire h_u_cla24_and1965_y0;
  wire h_u_cla24_and1966_y0;
  wire h_u_cla24_and1967_y0;
  wire h_u_cla24_and1968_y0;
  wire h_u_cla24_and1969_y0;
  wire h_u_cla24_and1970_y0;
  wire h_u_cla24_and1971_y0;
  wire h_u_cla24_and1972_y0;
  wire h_u_cla24_and1973_y0;
  wire h_u_cla24_and1974_y0;
  wire h_u_cla24_and1975_y0;
  wire h_u_cla24_and1976_y0;
  wire h_u_cla24_and1977_y0;
  wire h_u_cla24_and1978_y0;
  wire h_u_cla24_and1979_y0;
  wire h_u_cla24_and1980_y0;
  wire h_u_cla24_and1981_y0;
  wire h_u_cla24_and1982_y0;
  wire h_u_cla24_and1983_y0;
  wire h_u_cla24_and1984_y0;
  wire h_u_cla24_and1985_y0;
  wire h_u_cla24_and1986_y0;
  wire h_u_cla24_and1987_y0;
  wire h_u_cla24_and1988_y0;
  wire h_u_cla24_and1989_y0;
  wire h_u_cla24_and1990_y0;
  wire h_u_cla24_and1991_y0;
  wire h_u_cla24_and1992_y0;
  wire h_u_cla24_and1993_y0;
  wire h_u_cla24_and1994_y0;
  wire h_u_cla24_and1995_y0;
  wire h_u_cla24_and1996_y0;
  wire h_u_cla24_and1997_y0;
  wire h_u_cla24_and1998_y0;
  wire h_u_cla24_and1999_y0;
  wire h_u_cla24_and2000_y0;
  wire h_u_cla24_and2001_y0;
  wire h_u_cla24_and2002_y0;
  wire h_u_cla24_and2003_y0;
  wire h_u_cla24_and2004_y0;
  wire h_u_cla24_and2005_y0;
  wire h_u_cla24_and2006_y0;
  wire h_u_cla24_and2007_y0;
  wire h_u_cla24_and2008_y0;
  wire h_u_cla24_and2009_y0;
  wire h_u_cla24_and2010_y0;
  wire h_u_cla24_and2011_y0;
  wire h_u_cla24_and2012_y0;
  wire h_u_cla24_and2013_y0;
  wire h_u_cla24_and2014_y0;
  wire h_u_cla24_and2015_y0;
  wire h_u_cla24_and2016_y0;
  wire h_u_cla24_and2017_y0;
  wire h_u_cla24_and2018_y0;
  wire h_u_cla24_and2019_y0;
  wire h_u_cla24_and2020_y0;
  wire h_u_cla24_and2021_y0;
  wire h_u_cla24_and2022_y0;
  wire h_u_cla24_and2023_y0;
  wire h_u_cla24_and2024_y0;
  wire h_u_cla24_and2025_y0;
  wire h_u_cla24_and2026_y0;
  wire h_u_cla24_and2027_y0;
  wire h_u_cla24_and2028_y0;
  wire h_u_cla24_and2029_y0;
  wire h_u_cla24_and2030_y0;
  wire h_u_cla24_and2031_y0;
  wire h_u_cla24_and2032_y0;
  wire h_u_cla24_and2033_y0;
  wire h_u_cla24_and2034_y0;
  wire h_u_cla24_and2035_y0;
  wire h_u_cla24_and2036_y0;
  wire h_u_cla24_and2037_y0;
  wire h_u_cla24_and2038_y0;
  wire h_u_cla24_and2039_y0;
  wire h_u_cla24_and2040_y0;
  wire h_u_cla24_and2041_y0;
  wire h_u_cla24_and2042_y0;
  wire h_u_cla24_and2043_y0;
  wire h_u_cla24_and2044_y0;
  wire h_u_cla24_and2045_y0;
  wire h_u_cla24_and2046_y0;
  wire h_u_cla24_and2047_y0;
  wire h_u_cla24_and2048_y0;
  wire h_u_cla24_and2049_y0;
  wire h_u_cla24_and2050_y0;
  wire h_u_cla24_and2051_y0;
  wire h_u_cla24_and2052_y0;
  wire h_u_cla24_and2053_y0;
  wire h_u_cla24_and2054_y0;
  wire h_u_cla24_and2055_y0;
  wire h_u_cla24_and2056_y0;
  wire h_u_cla24_and2057_y0;
  wire h_u_cla24_and2058_y0;
  wire h_u_cla24_and2059_y0;
  wire h_u_cla24_and2060_y0;
  wire h_u_cla24_and2061_y0;
  wire h_u_cla24_and2062_y0;
  wire h_u_cla24_and2063_y0;
  wire h_u_cla24_and2064_y0;
  wire h_u_cla24_and2065_y0;
  wire h_u_cla24_and2066_y0;
  wire h_u_cla24_and2067_y0;
  wire h_u_cla24_and2068_y0;
  wire h_u_cla24_and2069_y0;
  wire h_u_cla24_and2070_y0;
  wire h_u_cla24_and2071_y0;
  wire h_u_cla24_and2072_y0;
  wire h_u_cla24_and2073_y0;
  wire h_u_cla24_and2074_y0;
  wire h_u_cla24_and2075_y0;
  wire h_u_cla24_and2076_y0;
  wire h_u_cla24_and2077_y0;
  wire h_u_cla24_and2078_y0;
  wire h_u_cla24_and2079_y0;
  wire h_u_cla24_and2080_y0;
  wire h_u_cla24_and2081_y0;
  wire h_u_cla24_and2082_y0;
  wire h_u_cla24_and2083_y0;
  wire h_u_cla24_and2084_y0;
  wire h_u_cla24_and2085_y0;
  wire h_u_cla24_and2086_y0;
  wire h_u_cla24_and2087_y0;
  wire h_u_cla24_and2088_y0;
  wire h_u_cla24_and2089_y0;
  wire h_u_cla24_and2090_y0;
  wire h_u_cla24_and2091_y0;
  wire h_u_cla24_and2092_y0;
  wire h_u_cla24_and2093_y0;
  wire h_u_cla24_and2094_y0;
  wire h_u_cla24_and2095_y0;
  wire h_u_cla24_and2096_y0;
  wire h_u_cla24_and2097_y0;
  wire h_u_cla24_and2098_y0;
  wire h_u_cla24_and2099_y0;
  wire h_u_cla24_and2100_y0;
  wire h_u_cla24_and2101_y0;
  wire h_u_cla24_and2102_y0;
  wire h_u_cla24_and2103_y0;
  wire h_u_cla24_and2104_y0;
  wire h_u_cla24_and2105_y0;
  wire h_u_cla24_and2106_y0;
  wire h_u_cla24_and2107_y0;
  wire h_u_cla24_and2108_y0;
  wire h_u_cla24_or153_y0;
  wire h_u_cla24_or154_y0;
  wire h_u_cla24_or155_y0;
  wire h_u_cla24_or156_y0;
  wire h_u_cla24_or157_y0;
  wire h_u_cla24_or158_y0;
  wire h_u_cla24_or159_y0;
  wire h_u_cla24_or160_y0;
  wire h_u_cla24_or161_y0;
  wire h_u_cla24_or162_y0;
  wire h_u_cla24_or163_y0;
  wire h_u_cla24_or164_y0;
  wire h_u_cla24_or165_y0;
  wire h_u_cla24_or166_y0;
  wire h_u_cla24_or167_y0;
  wire h_u_cla24_or168_y0;
  wire h_u_cla24_or169_y0;
  wire h_u_cla24_or170_y0;
  wire h_u_cla24_pg_logic18_y0;
  wire h_u_cla24_pg_logic18_y1;
  wire h_u_cla24_pg_logic18_y2;
  wire h_u_cla24_xor18_y0;
  wire h_u_cla24_and2109_y0;
  wire h_u_cla24_and2110_y0;
  wire h_u_cla24_and2111_y0;
  wire h_u_cla24_and2112_y0;
  wire h_u_cla24_and2113_y0;
  wire h_u_cla24_and2114_y0;
  wire h_u_cla24_and2115_y0;
  wire h_u_cla24_and2116_y0;
  wire h_u_cla24_and2117_y0;
  wire h_u_cla24_and2118_y0;
  wire h_u_cla24_and2119_y0;
  wire h_u_cla24_and2120_y0;
  wire h_u_cla24_and2121_y0;
  wire h_u_cla24_and2122_y0;
  wire h_u_cla24_and2123_y0;
  wire h_u_cla24_and2124_y0;
  wire h_u_cla24_and2125_y0;
  wire h_u_cla24_and2126_y0;
  wire h_u_cla24_and2127_y0;
  wire h_u_cla24_and2128_y0;
  wire h_u_cla24_and2129_y0;
  wire h_u_cla24_and2130_y0;
  wire h_u_cla24_and2131_y0;
  wire h_u_cla24_and2132_y0;
  wire h_u_cla24_and2133_y0;
  wire h_u_cla24_and2134_y0;
  wire h_u_cla24_and2135_y0;
  wire h_u_cla24_and2136_y0;
  wire h_u_cla24_and2137_y0;
  wire h_u_cla24_and2138_y0;
  wire h_u_cla24_and2139_y0;
  wire h_u_cla24_and2140_y0;
  wire h_u_cla24_and2141_y0;
  wire h_u_cla24_and2142_y0;
  wire h_u_cla24_and2143_y0;
  wire h_u_cla24_and2144_y0;
  wire h_u_cla24_and2145_y0;
  wire h_u_cla24_and2146_y0;
  wire h_u_cla24_and2147_y0;
  wire h_u_cla24_and2148_y0;
  wire h_u_cla24_and2149_y0;
  wire h_u_cla24_and2150_y0;
  wire h_u_cla24_and2151_y0;
  wire h_u_cla24_and2152_y0;
  wire h_u_cla24_and2153_y0;
  wire h_u_cla24_and2154_y0;
  wire h_u_cla24_and2155_y0;
  wire h_u_cla24_and2156_y0;
  wire h_u_cla24_and2157_y0;
  wire h_u_cla24_and2158_y0;
  wire h_u_cla24_and2159_y0;
  wire h_u_cla24_and2160_y0;
  wire h_u_cla24_and2161_y0;
  wire h_u_cla24_and2162_y0;
  wire h_u_cla24_and2163_y0;
  wire h_u_cla24_and2164_y0;
  wire h_u_cla24_and2165_y0;
  wire h_u_cla24_and2166_y0;
  wire h_u_cla24_and2167_y0;
  wire h_u_cla24_and2168_y0;
  wire h_u_cla24_and2169_y0;
  wire h_u_cla24_and2170_y0;
  wire h_u_cla24_and2171_y0;
  wire h_u_cla24_and2172_y0;
  wire h_u_cla24_and2173_y0;
  wire h_u_cla24_and2174_y0;
  wire h_u_cla24_and2175_y0;
  wire h_u_cla24_and2176_y0;
  wire h_u_cla24_and2177_y0;
  wire h_u_cla24_and2178_y0;
  wire h_u_cla24_and2179_y0;
  wire h_u_cla24_and2180_y0;
  wire h_u_cla24_and2181_y0;
  wire h_u_cla24_and2182_y0;
  wire h_u_cla24_and2183_y0;
  wire h_u_cla24_and2184_y0;
  wire h_u_cla24_and2185_y0;
  wire h_u_cla24_and2186_y0;
  wire h_u_cla24_and2187_y0;
  wire h_u_cla24_and2188_y0;
  wire h_u_cla24_and2189_y0;
  wire h_u_cla24_and2190_y0;
  wire h_u_cla24_and2191_y0;
  wire h_u_cla24_and2192_y0;
  wire h_u_cla24_and2193_y0;
  wire h_u_cla24_and2194_y0;
  wire h_u_cla24_and2195_y0;
  wire h_u_cla24_and2196_y0;
  wire h_u_cla24_and2197_y0;
  wire h_u_cla24_and2198_y0;
  wire h_u_cla24_and2199_y0;
  wire h_u_cla24_and2200_y0;
  wire h_u_cla24_and2201_y0;
  wire h_u_cla24_and2202_y0;
  wire h_u_cla24_and2203_y0;
  wire h_u_cla24_and2204_y0;
  wire h_u_cla24_and2205_y0;
  wire h_u_cla24_and2206_y0;
  wire h_u_cla24_and2207_y0;
  wire h_u_cla24_and2208_y0;
  wire h_u_cla24_and2209_y0;
  wire h_u_cla24_and2210_y0;
  wire h_u_cla24_and2211_y0;
  wire h_u_cla24_and2212_y0;
  wire h_u_cla24_and2213_y0;
  wire h_u_cla24_and2214_y0;
  wire h_u_cla24_and2215_y0;
  wire h_u_cla24_and2216_y0;
  wire h_u_cla24_and2217_y0;
  wire h_u_cla24_and2218_y0;
  wire h_u_cla24_and2219_y0;
  wire h_u_cla24_and2220_y0;
  wire h_u_cla24_and2221_y0;
  wire h_u_cla24_and2222_y0;
  wire h_u_cla24_and2223_y0;
  wire h_u_cla24_and2224_y0;
  wire h_u_cla24_and2225_y0;
  wire h_u_cla24_and2226_y0;
  wire h_u_cla24_and2227_y0;
  wire h_u_cla24_and2228_y0;
  wire h_u_cla24_and2229_y0;
  wire h_u_cla24_and2230_y0;
  wire h_u_cla24_and2231_y0;
  wire h_u_cla24_and2232_y0;
  wire h_u_cla24_and2233_y0;
  wire h_u_cla24_and2234_y0;
  wire h_u_cla24_and2235_y0;
  wire h_u_cla24_and2236_y0;
  wire h_u_cla24_and2237_y0;
  wire h_u_cla24_and2238_y0;
  wire h_u_cla24_and2239_y0;
  wire h_u_cla24_and2240_y0;
  wire h_u_cla24_and2241_y0;
  wire h_u_cla24_and2242_y0;
  wire h_u_cla24_and2243_y0;
  wire h_u_cla24_and2244_y0;
  wire h_u_cla24_and2245_y0;
  wire h_u_cla24_and2246_y0;
  wire h_u_cla24_and2247_y0;
  wire h_u_cla24_and2248_y0;
  wire h_u_cla24_and2249_y0;
  wire h_u_cla24_and2250_y0;
  wire h_u_cla24_and2251_y0;
  wire h_u_cla24_and2252_y0;
  wire h_u_cla24_and2253_y0;
  wire h_u_cla24_and2254_y0;
  wire h_u_cla24_and2255_y0;
  wire h_u_cla24_and2256_y0;
  wire h_u_cla24_and2257_y0;
  wire h_u_cla24_and2258_y0;
  wire h_u_cla24_and2259_y0;
  wire h_u_cla24_and2260_y0;
  wire h_u_cla24_and2261_y0;
  wire h_u_cla24_and2262_y0;
  wire h_u_cla24_and2263_y0;
  wire h_u_cla24_and2264_y0;
  wire h_u_cla24_and2265_y0;
  wire h_u_cla24_and2266_y0;
  wire h_u_cla24_and2267_y0;
  wire h_u_cla24_and2268_y0;
  wire h_u_cla24_and2269_y0;
  wire h_u_cla24_and2270_y0;
  wire h_u_cla24_and2271_y0;
  wire h_u_cla24_and2272_y0;
  wire h_u_cla24_and2273_y0;
  wire h_u_cla24_and2274_y0;
  wire h_u_cla24_and2275_y0;
  wire h_u_cla24_and2276_y0;
  wire h_u_cla24_and2277_y0;
  wire h_u_cla24_and2278_y0;
  wire h_u_cla24_and2279_y0;
  wire h_u_cla24_and2280_y0;
  wire h_u_cla24_and2281_y0;
  wire h_u_cla24_and2282_y0;
  wire h_u_cla24_and2283_y0;
  wire h_u_cla24_and2284_y0;
  wire h_u_cla24_and2285_y0;
  wire h_u_cla24_and2286_y0;
  wire h_u_cla24_and2287_y0;
  wire h_u_cla24_and2288_y0;
  wire h_u_cla24_and2289_y0;
  wire h_u_cla24_and2290_y0;
  wire h_u_cla24_and2291_y0;
  wire h_u_cla24_and2292_y0;
  wire h_u_cla24_and2293_y0;
  wire h_u_cla24_and2294_y0;
  wire h_u_cla24_and2295_y0;
  wire h_u_cla24_and2296_y0;
  wire h_u_cla24_and2297_y0;
  wire h_u_cla24_and2298_y0;
  wire h_u_cla24_and2299_y0;
  wire h_u_cla24_and2300_y0;
  wire h_u_cla24_and2301_y0;
  wire h_u_cla24_and2302_y0;
  wire h_u_cla24_and2303_y0;
  wire h_u_cla24_and2304_y0;
  wire h_u_cla24_and2305_y0;
  wire h_u_cla24_and2306_y0;
  wire h_u_cla24_and2307_y0;
  wire h_u_cla24_and2308_y0;
  wire h_u_cla24_and2309_y0;
  wire h_u_cla24_and2310_y0;
  wire h_u_cla24_and2311_y0;
  wire h_u_cla24_and2312_y0;
  wire h_u_cla24_and2313_y0;
  wire h_u_cla24_and2314_y0;
  wire h_u_cla24_and2315_y0;
  wire h_u_cla24_and2316_y0;
  wire h_u_cla24_and2317_y0;
  wire h_u_cla24_and2318_y0;
  wire h_u_cla24_and2319_y0;
  wire h_u_cla24_and2320_y0;
  wire h_u_cla24_and2321_y0;
  wire h_u_cla24_and2322_y0;
  wire h_u_cla24_and2323_y0;
  wire h_u_cla24_and2324_y0;
  wire h_u_cla24_and2325_y0;
  wire h_u_cla24_and2326_y0;
  wire h_u_cla24_and2327_y0;
  wire h_u_cla24_and2328_y0;
  wire h_u_cla24_and2329_y0;
  wire h_u_cla24_and2330_y0;
  wire h_u_cla24_and2331_y0;
  wire h_u_cla24_and2332_y0;
  wire h_u_cla24_and2333_y0;
  wire h_u_cla24_and2334_y0;
  wire h_u_cla24_and2335_y0;
  wire h_u_cla24_and2336_y0;
  wire h_u_cla24_and2337_y0;
  wire h_u_cla24_and2338_y0;
  wire h_u_cla24_and2339_y0;
  wire h_u_cla24_and2340_y0;
  wire h_u_cla24_and2341_y0;
  wire h_u_cla24_and2342_y0;
  wire h_u_cla24_and2343_y0;
  wire h_u_cla24_and2344_y0;
  wire h_u_cla24_and2345_y0;
  wire h_u_cla24_and2346_y0;
  wire h_u_cla24_and2347_y0;
  wire h_u_cla24_and2348_y0;
  wire h_u_cla24_and2349_y0;
  wire h_u_cla24_and2350_y0;
  wire h_u_cla24_and2351_y0;
  wire h_u_cla24_and2352_y0;
  wire h_u_cla24_and2353_y0;
  wire h_u_cla24_and2354_y0;
  wire h_u_cla24_and2355_y0;
  wire h_u_cla24_and2356_y0;
  wire h_u_cla24_and2357_y0;
  wire h_u_cla24_and2358_y0;
  wire h_u_cla24_and2359_y0;
  wire h_u_cla24_and2360_y0;
  wire h_u_cla24_and2361_y0;
  wire h_u_cla24_and2362_y0;
  wire h_u_cla24_and2363_y0;
  wire h_u_cla24_and2364_y0;
  wire h_u_cla24_and2365_y0;
  wire h_u_cla24_and2366_y0;
  wire h_u_cla24_and2367_y0;
  wire h_u_cla24_and2368_y0;
  wire h_u_cla24_and2369_y0;
  wire h_u_cla24_and2370_y0;
  wire h_u_cla24_and2371_y0;
  wire h_u_cla24_and2372_y0;
  wire h_u_cla24_and2373_y0;
  wire h_u_cla24_and2374_y0;
  wire h_u_cla24_and2375_y0;
  wire h_u_cla24_and2376_y0;
  wire h_u_cla24_and2377_y0;
  wire h_u_cla24_and2378_y0;
  wire h_u_cla24_and2379_y0;
  wire h_u_cla24_and2380_y0;
  wire h_u_cla24_and2381_y0;
  wire h_u_cla24_and2382_y0;
  wire h_u_cla24_and2383_y0;
  wire h_u_cla24_and2384_y0;
  wire h_u_cla24_and2385_y0;
  wire h_u_cla24_and2386_y0;
  wire h_u_cla24_and2387_y0;
  wire h_u_cla24_and2388_y0;
  wire h_u_cla24_and2389_y0;
  wire h_u_cla24_and2390_y0;
  wire h_u_cla24_and2391_y0;
  wire h_u_cla24_and2392_y0;
  wire h_u_cla24_and2393_y0;
  wire h_u_cla24_and2394_y0;
  wire h_u_cla24_and2395_y0;
  wire h_u_cla24_and2396_y0;
  wire h_u_cla24_and2397_y0;
  wire h_u_cla24_and2398_y0;
  wire h_u_cla24_and2399_y0;
  wire h_u_cla24_and2400_y0;
  wire h_u_cla24_and2401_y0;
  wire h_u_cla24_and2402_y0;
  wire h_u_cla24_and2403_y0;
  wire h_u_cla24_and2404_y0;
  wire h_u_cla24_and2405_y0;
  wire h_u_cla24_and2406_y0;
  wire h_u_cla24_and2407_y0;
  wire h_u_cla24_and2408_y0;
  wire h_u_cla24_and2409_y0;
  wire h_u_cla24_and2410_y0;
  wire h_u_cla24_and2411_y0;
  wire h_u_cla24_and2412_y0;
  wire h_u_cla24_and2413_y0;
  wire h_u_cla24_and2414_y0;
  wire h_u_cla24_and2415_y0;
  wire h_u_cla24_and2416_y0;
  wire h_u_cla24_and2417_y0;
  wire h_u_cla24_and2418_y0;
  wire h_u_cla24_and2419_y0;
  wire h_u_cla24_and2420_y0;
  wire h_u_cla24_and2421_y0;
  wire h_u_cla24_and2422_y0;
  wire h_u_cla24_and2423_y0;
  wire h_u_cla24_and2424_y0;
  wire h_u_cla24_and2425_y0;
  wire h_u_cla24_and2426_y0;
  wire h_u_cla24_and2427_y0;
  wire h_u_cla24_and2428_y0;
  wire h_u_cla24_and2429_y0;
  wire h_u_cla24_and2430_y0;
  wire h_u_cla24_and2431_y0;
  wire h_u_cla24_and2432_y0;
  wire h_u_cla24_and2433_y0;
  wire h_u_cla24_and2434_y0;
  wire h_u_cla24_and2435_y0;
  wire h_u_cla24_and2436_y0;
  wire h_u_cla24_and2437_y0;
  wire h_u_cla24_and2438_y0;
  wire h_u_cla24_and2439_y0;
  wire h_u_cla24_and2440_y0;
  wire h_u_cla24_and2441_y0;
  wire h_u_cla24_and2442_y0;
  wire h_u_cla24_and2443_y0;
  wire h_u_cla24_and2444_y0;
  wire h_u_cla24_and2445_y0;
  wire h_u_cla24_and2446_y0;
  wire h_u_cla24_and2447_y0;
  wire h_u_cla24_and2448_y0;
  wire h_u_cla24_and2449_y0;
  wire h_u_cla24_and2450_y0;
  wire h_u_cla24_and2451_y0;
  wire h_u_cla24_and2452_y0;
  wire h_u_cla24_and2453_y0;
  wire h_u_cla24_and2454_y0;
  wire h_u_cla24_and2455_y0;
  wire h_u_cla24_and2456_y0;
  wire h_u_cla24_and2457_y0;
  wire h_u_cla24_and2458_y0;
  wire h_u_cla24_and2459_y0;
  wire h_u_cla24_and2460_y0;
  wire h_u_cla24_and2461_y0;
  wire h_u_cla24_and2462_y0;
  wire h_u_cla24_and2463_y0;
  wire h_u_cla24_and2464_y0;
  wire h_u_cla24_and2465_y0;
  wire h_u_cla24_and2466_y0;
  wire h_u_cla24_and2467_y0;
  wire h_u_cla24_and2468_y0;
  wire h_u_cla24_and2469_y0;
  wire h_u_cla24_or171_y0;
  wire h_u_cla24_or172_y0;
  wire h_u_cla24_or173_y0;
  wire h_u_cla24_or174_y0;
  wire h_u_cla24_or175_y0;
  wire h_u_cla24_or176_y0;
  wire h_u_cla24_or177_y0;
  wire h_u_cla24_or178_y0;
  wire h_u_cla24_or179_y0;
  wire h_u_cla24_or180_y0;
  wire h_u_cla24_or181_y0;
  wire h_u_cla24_or182_y0;
  wire h_u_cla24_or183_y0;
  wire h_u_cla24_or184_y0;
  wire h_u_cla24_or185_y0;
  wire h_u_cla24_or186_y0;
  wire h_u_cla24_or187_y0;
  wire h_u_cla24_or188_y0;
  wire h_u_cla24_or189_y0;
  wire h_u_cla24_pg_logic19_y0;
  wire h_u_cla24_pg_logic19_y1;
  wire h_u_cla24_pg_logic19_y2;
  wire h_u_cla24_xor19_y0;
  wire h_u_cla24_and2470_y0;
  wire h_u_cla24_and2471_y0;
  wire h_u_cla24_and2472_y0;
  wire h_u_cla24_and2473_y0;
  wire h_u_cla24_and2474_y0;
  wire h_u_cla24_and2475_y0;
  wire h_u_cla24_and2476_y0;
  wire h_u_cla24_and2477_y0;
  wire h_u_cla24_and2478_y0;
  wire h_u_cla24_and2479_y0;
  wire h_u_cla24_and2480_y0;
  wire h_u_cla24_and2481_y0;
  wire h_u_cla24_and2482_y0;
  wire h_u_cla24_and2483_y0;
  wire h_u_cla24_and2484_y0;
  wire h_u_cla24_and2485_y0;
  wire h_u_cla24_and2486_y0;
  wire h_u_cla24_and2487_y0;
  wire h_u_cla24_and2488_y0;
  wire h_u_cla24_and2489_y0;
  wire h_u_cla24_and2490_y0;
  wire h_u_cla24_and2491_y0;
  wire h_u_cla24_and2492_y0;
  wire h_u_cla24_and2493_y0;
  wire h_u_cla24_and2494_y0;
  wire h_u_cla24_and2495_y0;
  wire h_u_cla24_and2496_y0;
  wire h_u_cla24_and2497_y0;
  wire h_u_cla24_and2498_y0;
  wire h_u_cla24_and2499_y0;
  wire h_u_cla24_and2500_y0;
  wire h_u_cla24_and2501_y0;
  wire h_u_cla24_and2502_y0;
  wire h_u_cla24_and2503_y0;
  wire h_u_cla24_and2504_y0;
  wire h_u_cla24_and2505_y0;
  wire h_u_cla24_and2506_y0;
  wire h_u_cla24_and2507_y0;
  wire h_u_cla24_and2508_y0;
  wire h_u_cla24_and2509_y0;
  wire h_u_cla24_and2510_y0;
  wire h_u_cla24_and2511_y0;
  wire h_u_cla24_and2512_y0;
  wire h_u_cla24_and2513_y0;
  wire h_u_cla24_and2514_y0;
  wire h_u_cla24_and2515_y0;
  wire h_u_cla24_and2516_y0;
  wire h_u_cla24_and2517_y0;
  wire h_u_cla24_and2518_y0;
  wire h_u_cla24_and2519_y0;
  wire h_u_cla24_and2520_y0;
  wire h_u_cla24_and2521_y0;
  wire h_u_cla24_and2522_y0;
  wire h_u_cla24_and2523_y0;
  wire h_u_cla24_and2524_y0;
  wire h_u_cla24_and2525_y0;
  wire h_u_cla24_and2526_y0;
  wire h_u_cla24_and2527_y0;
  wire h_u_cla24_and2528_y0;
  wire h_u_cla24_and2529_y0;
  wire h_u_cla24_and2530_y0;
  wire h_u_cla24_and2531_y0;
  wire h_u_cla24_and2532_y0;
  wire h_u_cla24_and2533_y0;
  wire h_u_cla24_and2534_y0;
  wire h_u_cla24_and2535_y0;
  wire h_u_cla24_and2536_y0;
  wire h_u_cla24_and2537_y0;
  wire h_u_cla24_and2538_y0;
  wire h_u_cla24_and2539_y0;
  wire h_u_cla24_and2540_y0;
  wire h_u_cla24_and2541_y0;
  wire h_u_cla24_and2542_y0;
  wire h_u_cla24_and2543_y0;
  wire h_u_cla24_and2544_y0;
  wire h_u_cla24_and2545_y0;
  wire h_u_cla24_and2546_y0;
  wire h_u_cla24_and2547_y0;
  wire h_u_cla24_and2548_y0;
  wire h_u_cla24_and2549_y0;
  wire h_u_cla24_and2550_y0;
  wire h_u_cla24_and2551_y0;
  wire h_u_cla24_and2552_y0;
  wire h_u_cla24_and2553_y0;
  wire h_u_cla24_and2554_y0;
  wire h_u_cla24_and2555_y0;
  wire h_u_cla24_and2556_y0;
  wire h_u_cla24_and2557_y0;
  wire h_u_cla24_and2558_y0;
  wire h_u_cla24_and2559_y0;
  wire h_u_cla24_and2560_y0;
  wire h_u_cla24_and2561_y0;
  wire h_u_cla24_and2562_y0;
  wire h_u_cla24_and2563_y0;
  wire h_u_cla24_and2564_y0;
  wire h_u_cla24_and2565_y0;
  wire h_u_cla24_and2566_y0;
  wire h_u_cla24_and2567_y0;
  wire h_u_cla24_and2568_y0;
  wire h_u_cla24_and2569_y0;
  wire h_u_cla24_and2570_y0;
  wire h_u_cla24_and2571_y0;
  wire h_u_cla24_and2572_y0;
  wire h_u_cla24_and2573_y0;
  wire h_u_cla24_and2574_y0;
  wire h_u_cla24_and2575_y0;
  wire h_u_cla24_and2576_y0;
  wire h_u_cla24_and2577_y0;
  wire h_u_cla24_and2578_y0;
  wire h_u_cla24_and2579_y0;
  wire h_u_cla24_and2580_y0;
  wire h_u_cla24_and2581_y0;
  wire h_u_cla24_and2582_y0;
  wire h_u_cla24_and2583_y0;
  wire h_u_cla24_and2584_y0;
  wire h_u_cla24_and2585_y0;
  wire h_u_cla24_and2586_y0;
  wire h_u_cla24_and2587_y0;
  wire h_u_cla24_and2588_y0;
  wire h_u_cla24_and2589_y0;
  wire h_u_cla24_and2590_y0;
  wire h_u_cla24_and2591_y0;
  wire h_u_cla24_and2592_y0;
  wire h_u_cla24_and2593_y0;
  wire h_u_cla24_and2594_y0;
  wire h_u_cla24_and2595_y0;
  wire h_u_cla24_and2596_y0;
  wire h_u_cla24_and2597_y0;
  wire h_u_cla24_and2598_y0;
  wire h_u_cla24_and2599_y0;
  wire h_u_cla24_and2600_y0;
  wire h_u_cla24_and2601_y0;
  wire h_u_cla24_and2602_y0;
  wire h_u_cla24_and2603_y0;
  wire h_u_cla24_and2604_y0;
  wire h_u_cla24_and2605_y0;
  wire h_u_cla24_and2606_y0;
  wire h_u_cla24_and2607_y0;
  wire h_u_cla24_and2608_y0;
  wire h_u_cla24_and2609_y0;
  wire h_u_cla24_and2610_y0;
  wire h_u_cla24_and2611_y0;
  wire h_u_cla24_and2612_y0;
  wire h_u_cla24_and2613_y0;
  wire h_u_cla24_and2614_y0;
  wire h_u_cla24_and2615_y0;
  wire h_u_cla24_and2616_y0;
  wire h_u_cla24_and2617_y0;
  wire h_u_cla24_and2618_y0;
  wire h_u_cla24_and2619_y0;
  wire h_u_cla24_and2620_y0;
  wire h_u_cla24_and2621_y0;
  wire h_u_cla24_and2622_y0;
  wire h_u_cla24_and2623_y0;
  wire h_u_cla24_and2624_y0;
  wire h_u_cla24_and2625_y0;
  wire h_u_cla24_and2626_y0;
  wire h_u_cla24_and2627_y0;
  wire h_u_cla24_and2628_y0;
  wire h_u_cla24_and2629_y0;
  wire h_u_cla24_and2630_y0;
  wire h_u_cla24_and2631_y0;
  wire h_u_cla24_and2632_y0;
  wire h_u_cla24_and2633_y0;
  wire h_u_cla24_and2634_y0;
  wire h_u_cla24_and2635_y0;
  wire h_u_cla24_and2636_y0;
  wire h_u_cla24_and2637_y0;
  wire h_u_cla24_and2638_y0;
  wire h_u_cla24_and2639_y0;
  wire h_u_cla24_and2640_y0;
  wire h_u_cla24_and2641_y0;
  wire h_u_cla24_and2642_y0;
  wire h_u_cla24_and2643_y0;
  wire h_u_cla24_and2644_y0;
  wire h_u_cla24_and2645_y0;
  wire h_u_cla24_and2646_y0;
  wire h_u_cla24_and2647_y0;
  wire h_u_cla24_and2648_y0;
  wire h_u_cla24_and2649_y0;
  wire h_u_cla24_and2650_y0;
  wire h_u_cla24_and2651_y0;
  wire h_u_cla24_and2652_y0;
  wire h_u_cla24_and2653_y0;
  wire h_u_cla24_and2654_y0;
  wire h_u_cla24_and2655_y0;
  wire h_u_cla24_and2656_y0;
  wire h_u_cla24_and2657_y0;
  wire h_u_cla24_and2658_y0;
  wire h_u_cla24_and2659_y0;
  wire h_u_cla24_and2660_y0;
  wire h_u_cla24_and2661_y0;
  wire h_u_cla24_and2662_y0;
  wire h_u_cla24_and2663_y0;
  wire h_u_cla24_and2664_y0;
  wire h_u_cla24_and2665_y0;
  wire h_u_cla24_and2666_y0;
  wire h_u_cla24_and2667_y0;
  wire h_u_cla24_and2668_y0;
  wire h_u_cla24_and2669_y0;
  wire h_u_cla24_and2670_y0;
  wire h_u_cla24_and2671_y0;
  wire h_u_cla24_and2672_y0;
  wire h_u_cla24_and2673_y0;
  wire h_u_cla24_and2674_y0;
  wire h_u_cla24_and2675_y0;
  wire h_u_cla24_and2676_y0;
  wire h_u_cla24_and2677_y0;
  wire h_u_cla24_and2678_y0;
  wire h_u_cla24_and2679_y0;
  wire h_u_cla24_and2680_y0;
  wire h_u_cla24_and2681_y0;
  wire h_u_cla24_and2682_y0;
  wire h_u_cla24_and2683_y0;
  wire h_u_cla24_and2684_y0;
  wire h_u_cla24_and2685_y0;
  wire h_u_cla24_and2686_y0;
  wire h_u_cla24_and2687_y0;
  wire h_u_cla24_and2688_y0;
  wire h_u_cla24_and2689_y0;
  wire h_u_cla24_and2690_y0;
  wire h_u_cla24_and2691_y0;
  wire h_u_cla24_and2692_y0;
  wire h_u_cla24_and2693_y0;
  wire h_u_cla24_and2694_y0;
  wire h_u_cla24_and2695_y0;
  wire h_u_cla24_and2696_y0;
  wire h_u_cla24_and2697_y0;
  wire h_u_cla24_and2698_y0;
  wire h_u_cla24_and2699_y0;
  wire h_u_cla24_and2700_y0;
  wire h_u_cla24_and2701_y0;
  wire h_u_cla24_and2702_y0;
  wire h_u_cla24_and2703_y0;
  wire h_u_cla24_and2704_y0;
  wire h_u_cla24_and2705_y0;
  wire h_u_cla24_and2706_y0;
  wire h_u_cla24_and2707_y0;
  wire h_u_cla24_and2708_y0;
  wire h_u_cla24_and2709_y0;
  wire h_u_cla24_and2710_y0;
  wire h_u_cla24_and2711_y0;
  wire h_u_cla24_and2712_y0;
  wire h_u_cla24_and2713_y0;
  wire h_u_cla24_and2714_y0;
  wire h_u_cla24_and2715_y0;
  wire h_u_cla24_and2716_y0;
  wire h_u_cla24_and2717_y0;
  wire h_u_cla24_and2718_y0;
  wire h_u_cla24_and2719_y0;
  wire h_u_cla24_and2720_y0;
  wire h_u_cla24_and2721_y0;
  wire h_u_cla24_and2722_y0;
  wire h_u_cla24_and2723_y0;
  wire h_u_cla24_and2724_y0;
  wire h_u_cla24_and2725_y0;
  wire h_u_cla24_and2726_y0;
  wire h_u_cla24_and2727_y0;
  wire h_u_cla24_and2728_y0;
  wire h_u_cla24_and2729_y0;
  wire h_u_cla24_and2730_y0;
  wire h_u_cla24_and2731_y0;
  wire h_u_cla24_and2732_y0;
  wire h_u_cla24_and2733_y0;
  wire h_u_cla24_and2734_y0;
  wire h_u_cla24_and2735_y0;
  wire h_u_cla24_and2736_y0;
  wire h_u_cla24_and2737_y0;
  wire h_u_cla24_and2738_y0;
  wire h_u_cla24_and2739_y0;
  wire h_u_cla24_and2740_y0;
  wire h_u_cla24_and2741_y0;
  wire h_u_cla24_and2742_y0;
  wire h_u_cla24_and2743_y0;
  wire h_u_cla24_and2744_y0;
  wire h_u_cla24_and2745_y0;
  wire h_u_cla24_and2746_y0;
  wire h_u_cla24_and2747_y0;
  wire h_u_cla24_and2748_y0;
  wire h_u_cla24_and2749_y0;
  wire h_u_cla24_and2750_y0;
  wire h_u_cla24_and2751_y0;
  wire h_u_cla24_and2752_y0;
  wire h_u_cla24_and2753_y0;
  wire h_u_cla24_and2754_y0;
  wire h_u_cla24_and2755_y0;
  wire h_u_cla24_and2756_y0;
  wire h_u_cla24_and2757_y0;
  wire h_u_cla24_and2758_y0;
  wire h_u_cla24_and2759_y0;
  wire h_u_cla24_and2760_y0;
  wire h_u_cla24_and2761_y0;
  wire h_u_cla24_and2762_y0;
  wire h_u_cla24_and2763_y0;
  wire h_u_cla24_and2764_y0;
  wire h_u_cla24_and2765_y0;
  wire h_u_cla24_and2766_y0;
  wire h_u_cla24_and2767_y0;
  wire h_u_cla24_and2768_y0;
  wire h_u_cla24_and2769_y0;
  wire h_u_cla24_and2770_y0;
  wire h_u_cla24_and2771_y0;
  wire h_u_cla24_and2772_y0;
  wire h_u_cla24_and2773_y0;
  wire h_u_cla24_and2774_y0;
  wire h_u_cla24_and2775_y0;
  wire h_u_cla24_and2776_y0;
  wire h_u_cla24_and2777_y0;
  wire h_u_cla24_and2778_y0;
  wire h_u_cla24_and2779_y0;
  wire h_u_cla24_and2780_y0;
  wire h_u_cla24_and2781_y0;
  wire h_u_cla24_and2782_y0;
  wire h_u_cla24_and2783_y0;
  wire h_u_cla24_and2784_y0;
  wire h_u_cla24_and2785_y0;
  wire h_u_cla24_and2786_y0;
  wire h_u_cla24_and2787_y0;
  wire h_u_cla24_and2788_y0;
  wire h_u_cla24_and2789_y0;
  wire h_u_cla24_and2790_y0;
  wire h_u_cla24_and2791_y0;
  wire h_u_cla24_and2792_y0;
  wire h_u_cla24_and2793_y0;
  wire h_u_cla24_and2794_y0;
  wire h_u_cla24_and2795_y0;
  wire h_u_cla24_and2796_y0;
  wire h_u_cla24_and2797_y0;
  wire h_u_cla24_and2798_y0;
  wire h_u_cla24_and2799_y0;
  wire h_u_cla24_and2800_y0;
  wire h_u_cla24_and2801_y0;
  wire h_u_cla24_and2802_y0;
  wire h_u_cla24_and2803_y0;
  wire h_u_cla24_and2804_y0;
  wire h_u_cla24_and2805_y0;
  wire h_u_cla24_and2806_y0;
  wire h_u_cla24_and2807_y0;
  wire h_u_cla24_and2808_y0;
  wire h_u_cla24_and2809_y0;
  wire h_u_cla24_and2810_y0;
  wire h_u_cla24_and2811_y0;
  wire h_u_cla24_and2812_y0;
  wire h_u_cla24_and2813_y0;
  wire h_u_cla24_and2814_y0;
  wire h_u_cla24_and2815_y0;
  wire h_u_cla24_and2816_y0;
  wire h_u_cla24_and2817_y0;
  wire h_u_cla24_and2818_y0;
  wire h_u_cla24_and2819_y0;
  wire h_u_cla24_and2820_y0;
  wire h_u_cla24_and2821_y0;
  wire h_u_cla24_and2822_y0;
  wire h_u_cla24_and2823_y0;
  wire h_u_cla24_and2824_y0;
  wire h_u_cla24_and2825_y0;
  wire h_u_cla24_and2826_y0;
  wire h_u_cla24_and2827_y0;
  wire h_u_cla24_and2828_y0;
  wire h_u_cla24_and2829_y0;
  wire h_u_cla24_and2830_y0;
  wire h_u_cla24_and2831_y0;
  wire h_u_cla24_and2832_y0;
  wire h_u_cla24_and2833_y0;
  wire h_u_cla24_and2834_y0;
  wire h_u_cla24_and2835_y0;
  wire h_u_cla24_and2836_y0;
  wire h_u_cla24_and2837_y0;
  wire h_u_cla24_and2838_y0;
  wire h_u_cla24_and2839_y0;
  wire h_u_cla24_and2840_y0;
  wire h_u_cla24_and2841_y0;
  wire h_u_cla24_and2842_y0;
  wire h_u_cla24_and2843_y0;
  wire h_u_cla24_and2844_y0;
  wire h_u_cla24_and2845_y0;
  wire h_u_cla24_and2846_y0;
  wire h_u_cla24_and2847_y0;
  wire h_u_cla24_and2848_y0;
  wire h_u_cla24_and2849_y0;
  wire h_u_cla24_and2850_y0;
  wire h_u_cla24_and2851_y0;
  wire h_u_cla24_and2852_y0;
  wire h_u_cla24_and2853_y0;
  wire h_u_cla24_and2854_y0;
  wire h_u_cla24_and2855_y0;
  wire h_u_cla24_and2856_y0;
  wire h_u_cla24_and2857_y0;
  wire h_u_cla24_and2858_y0;
  wire h_u_cla24_and2859_y0;
  wire h_u_cla24_and2860_y0;
  wire h_u_cla24_and2861_y0;
  wire h_u_cla24_and2862_y0;
  wire h_u_cla24_and2863_y0;
  wire h_u_cla24_and2864_y0;
  wire h_u_cla24_and2865_y0;
  wire h_u_cla24_and2866_y0;
  wire h_u_cla24_and2867_y0;
  wire h_u_cla24_and2868_y0;
  wire h_u_cla24_and2869_y0;
  wire h_u_cla24_or190_y0;
  wire h_u_cla24_or191_y0;
  wire h_u_cla24_or192_y0;
  wire h_u_cla24_or193_y0;
  wire h_u_cla24_or194_y0;
  wire h_u_cla24_or195_y0;
  wire h_u_cla24_or196_y0;
  wire h_u_cla24_or197_y0;
  wire h_u_cla24_or198_y0;
  wire h_u_cla24_or199_y0;
  wire h_u_cla24_or200_y0;
  wire h_u_cla24_or201_y0;
  wire h_u_cla24_or202_y0;
  wire h_u_cla24_or203_y0;
  wire h_u_cla24_or204_y0;
  wire h_u_cla24_or205_y0;
  wire h_u_cla24_or206_y0;
  wire h_u_cla24_or207_y0;
  wire h_u_cla24_or208_y0;
  wire h_u_cla24_or209_y0;
  wire h_u_cla24_pg_logic20_y0;
  wire h_u_cla24_pg_logic20_y1;
  wire h_u_cla24_pg_logic20_y2;
  wire h_u_cla24_xor20_y0;
  wire h_u_cla24_and2870_y0;
  wire h_u_cla24_and2871_y0;
  wire h_u_cla24_and2872_y0;
  wire h_u_cla24_and2873_y0;
  wire h_u_cla24_and2874_y0;
  wire h_u_cla24_and2875_y0;
  wire h_u_cla24_and2876_y0;
  wire h_u_cla24_and2877_y0;
  wire h_u_cla24_and2878_y0;
  wire h_u_cla24_and2879_y0;
  wire h_u_cla24_and2880_y0;
  wire h_u_cla24_and2881_y0;
  wire h_u_cla24_and2882_y0;
  wire h_u_cla24_and2883_y0;
  wire h_u_cla24_and2884_y0;
  wire h_u_cla24_and2885_y0;
  wire h_u_cla24_and2886_y0;
  wire h_u_cla24_and2887_y0;
  wire h_u_cla24_and2888_y0;
  wire h_u_cla24_and2889_y0;
  wire h_u_cla24_and2890_y0;
  wire h_u_cla24_and2891_y0;
  wire h_u_cla24_and2892_y0;
  wire h_u_cla24_and2893_y0;
  wire h_u_cla24_and2894_y0;
  wire h_u_cla24_and2895_y0;
  wire h_u_cla24_and2896_y0;
  wire h_u_cla24_and2897_y0;
  wire h_u_cla24_and2898_y0;
  wire h_u_cla24_and2899_y0;
  wire h_u_cla24_and2900_y0;
  wire h_u_cla24_and2901_y0;
  wire h_u_cla24_and2902_y0;
  wire h_u_cla24_and2903_y0;
  wire h_u_cla24_and2904_y0;
  wire h_u_cla24_and2905_y0;
  wire h_u_cla24_and2906_y0;
  wire h_u_cla24_and2907_y0;
  wire h_u_cla24_and2908_y0;
  wire h_u_cla24_and2909_y0;
  wire h_u_cla24_and2910_y0;
  wire h_u_cla24_and2911_y0;
  wire h_u_cla24_and2912_y0;
  wire h_u_cla24_and2913_y0;
  wire h_u_cla24_and2914_y0;
  wire h_u_cla24_and2915_y0;
  wire h_u_cla24_and2916_y0;
  wire h_u_cla24_and2917_y0;
  wire h_u_cla24_and2918_y0;
  wire h_u_cla24_and2919_y0;
  wire h_u_cla24_and2920_y0;
  wire h_u_cla24_and2921_y0;
  wire h_u_cla24_and2922_y0;
  wire h_u_cla24_and2923_y0;
  wire h_u_cla24_and2924_y0;
  wire h_u_cla24_and2925_y0;
  wire h_u_cla24_and2926_y0;
  wire h_u_cla24_and2927_y0;
  wire h_u_cla24_and2928_y0;
  wire h_u_cla24_and2929_y0;
  wire h_u_cla24_and2930_y0;
  wire h_u_cla24_and2931_y0;
  wire h_u_cla24_and2932_y0;
  wire h_u_cla24_and2933_y0;
  wire h_u_cla24_and2934_y0;
  wire h_u_cla24_and2935_y0;
  wire h_u_cla24_and2936_y0;
  wire h_u_cla24_and2937_y0;
  wire h_u_cla24_and2938_y0;
  wire h_u_cla24_and2939_y0;
  wire h_u_cla24_and2940_y0;
  wire h_u_cla24_and2941_y0;
  wire h_u_cla24_and2942_y0;
  wire h_u_cla24_and2943_y0;
  wire h_u_cla24_and2944_y0;
  wire h_u_cla24_and2945_y0;
  wire h_u_cla24_and2946_y0;
  wire h_u_cla24_and2947_y0;
  wire h_u_cla24_and2948_y0;
  wire h_u_cla24_and2949_y0;
  wire h_u_cla24_and2950_y0;
  wire h_u_cla24_and2951_y0;
  wire h_u_cla24_and2952_y0;
  wire h_u_cla24_and2953_y0;
  wire h_u_cla24_and2954_y0;
  wire h_u_cla24_and2955_y0;
  wire h_u_cla24_and2956_y0;
  wire h_u_cla24_and2957_y0;
  wire h_u_cla24_and2958_y0;
  wire h_u_cla24_and2959_y0;
  wire h_u_cla24_and2960_y0;
  wire h_u_cla24_and2961_y0;
  wire h_u_cla24_and2962_y0;
  wire h_u_cla24_and2963_y0;
  wire h_u_cla24_and2964_y0;
  wire h_u_cla24_and2965_y0;
  wire h_u_cla24_and2966_y0;
  wire h_u_cla24_and2967_y0;
  wire h_u_cla24_and2968_y0;
  wire h_u_cla24_and2969_y0;
  wire h_u_cla24_and2970_y0;
  wire h_u_cla24_and2971_y0;
  wire h_u_cla24_and2972_y0;
  wire h_u_cla24_and2973_y0;
  wire h_u_cla24_and2974_y0;
  wire h_u_cla24_and2975_y0;
  wire h_u_cla24_and2976_y0;
  wire h_u_cla24_and2977_y0;
  wire h_u_cla24_and2978_y0;
  wire h_u_cla24_and2979_y0;
  wire h_u_cla24_and2980_y0;
  wire h_u_cla24_and2981_y0;
  wire h_u_cla24_and2982_y0;
  wire h_u_cla24_and2983_y0;
  wire h_u_cla24_and2984_y0;
  wire h_u_cla24_and2985_y0;
  wire h_u_cla24_and2986_y0;
  wire h_u_cla24_and2987_y0;
  wire h_u_cla24_and2988_y0;
  wire h_u_cla24_and2989_y0;
  wire h_u_cla24_and2990_y0;
  wire h_u_cla24_and2991_y0;
  wire h_u_cla24_and2992_y0;
  wire h_u_cla24_and2993_y0;
  wire h_u_cla24_and2994_y0;
  wire h_u_cla24_and2995_y0;
  wire h_u_cla24_and2996_y0;
  wire h_u_cla24_and2997_y0;
  wire h_u_cla24_and2998_y0;
  wire h_u_cla24_and2999_y0;
  wire h_u_cla24_and3000_y0;
  wire h_u_cla24_and3001_y0;
  wire h_u_cla24_and3002_y0;
  wire h_u_cla24_and3003_y0;
  wire h_u_cla24_and3004_y0;
  wire h_u_cla24_and3005_y0;
  wire h_u_cla24_and3006_y0;
  wire h_u_cla24_and3007_y0;
  wire h_u_cla24_and3008_y0;
  wire h_u_cla24_and3009_y0;
  wire h_u_cla24_and3010_y0;
  wire h_u_cla24_and3011_y0;
  wire h_u_cla24_and3012_y0;
  wire h_u_cla24_and3013_y0;
  wire h_u_cla24_and3014_y0;
  wire h_u_cla24_and3015_y0;
  wire h_u_cla24_and3016_y0;
  wire h_u_cla24_and3017_y0;
  wire h_u_cla24_and3018_y0;
  wire h_u_cla24_and3019_y0;
  wire h_u_cla24_and3020_y0;
  wire h_u_cla24_and3021_y0;
  wire h_u_cla24_and3022_y0;
  wire h_u_cla24_and3023_y0;
  wire h_u_cla24_and3024_y0;
  wire h_u_cla24_and3025_y0;
  wire h_u_cla24_and3026_y0;
  wire h_u_cla24_and3027_y0;
  wire h_u_cla24_and3028_y0;
  wire h_u_cla24_and3029_y0;
  wire h_u_cla24_and3030_y0;
  wire h_u_cla24_and3031_y0;
  wire h_u_cla24_and3032_y0;
  wire h_u_cla24_and3033_y0;
  wire h_u_cla24_and3034_y0;
  wire h_u_cla24_and3035_y0;
  wire h_u_cla24_and3036_y0;
  wire h_u_cla24_and3037_y0;
  wire h_u_cla24_and3038_y0;
  wire h_u_cla24_and3039_y0;
  wire h_u_cla24_and3040_y0;
  wire h_u_cla24_and3041_y0;
  wire h_u_cla24_and3042_y0;
  wire h_u_cla24_and3043_y0;
  wire h_u_cla24_and3044_y0;
  wire h_u_cla24_and3045_y0;
  wire h_u_cla24_and3046_y0;
  wire h_u_cla24_and3047_y0;
  wire h_u_cla24_and3048_y0;
  wire h_u_cla24_and3049_y0;
  wire h_u_cla24_and3050_y0;
  wire h_u_cla24_and3051_y0;
  wire h_u_cla24_and3052_y0;
  wire h_u_cla24_and3053_y0;
  wire h_u_cla24_and3054_y0;
  wire h_u_cla24_and3055_y0;
  wire h_u_cla24_and3056_y0;
  wire h_u_cla24_and3057_y0;
  wire h_u_cla24_and3058_y0;
  wire h_u_cla24_and3059_y0;
  wire h_u_cla24_and3060_y0;
  wire h_u_cla24_and3061_y0;
  wire h_u_cla24_and3062_y0;
  wire h_u_cla24_and3063_y0;
  wire h_u_cla24_and3064_y0;
  wire h_u_cla24_and3065_y0;
  wire h_u_cla24_and3066_y0;
  wire h_u_cla24_and3067_y0;
  wire h_u_cla24_and3068_y0;
  wire h_u_cla24_and3069_y0;
  wire h_u_cla24_and3070_y0;
  wire h_u_cla24_and3071_y0;
  wire h_u_cla24_and3072_y0;
  wire h_u_cla24_and3073_y0;
  wire h_u_cla24_and3074_y0;
  wire h_u_cla24_and3075_y0;
  wire h_u_cla24_and3076_y0;
  wire h_u_cla24_and3077_y0;
  wire h_u_cla24_and3078_y0;
  wire h_u_cla24_and3079_y0;
  wire h_u_cla24_and3080_y0;
  wire h_u_cla24_and3081_y0;
  wire h_u_cla24_and3082_y0;
  wire h_u_cla24_and3083_y0;
  wire h_u_cla24_and3084_y0;
  wire h_u_cla24_and3085_y0;
  wire h_u_cla24_and3086_y0;
  wire h_u_cla24_and3087_y0;
  wire h_u_cla24_and3088_y0;
  wire h_u_cla24_and3089_y0;
  wire h_u_cla24_and3090_y0;
  wire h_u_cla24_and3091_y0;
  wire h_u_cla24_and3092_y0;
  wire h_u_cla24_and3093_y0;
  wire h_u_cla24_and3094_y0;
  wire h_u_cla24_and3095_y0;
  wire h_u_cla24_and3096_y0;
  wire h_u_cla24_and3097_y0;
  wire h_u_cla24_and3098_y0;
  wire h_u_cla24_and3099_y0;
  wire h_u_cla24_and3100_y0;
  wire h_u_cla24_and3101_y0;
  wire h_u_cla24_and3102_y0;
  wire h_u_cla24_and3103_y0;
  wire h_u_cla24_and3104_y0;
  wire h_u_cla24_and3105_y0;
  wire h_u_cla24_and3106_y0;
  wire h_u_cla24_and3107_y0;
  wire h_u_cla24_and3108_y0;
  wire h_u_cla24_and3109_y0;
  wire h_u_cla24_and3110_y0;
  wire h_u_cla24_and3111_y0;
  wire h_u_cla24_and3112_y0;
  wire h_u_cla24_and3113_y0;
  wire h_u_cla24_and3114_y0;
  wire h_u_cla24_and3115_y0;
  wire h_u_cla24_and3116_y0;
  wire h_u_cla24_and3117_y0;
  wire h_u_cla24_and3118_y0;
  wire h_u_cla24_and3119_y0;
  wire h_u_cla24_and3120_y0;
  wire h_u_cla24_and3121_y0;
  wire h_u_cla24_and3122_y0;
  wire h_u_cla24_and3123_y0;
  wire h_u_cla24_and3124_y0;
  wire h_u_cla24_and3125_y0;
  wire h_u_cla24_and3126_y0;
  wire h_u_cla24_and3127_y0;
  wire h_u_cla24_and3128_y0;
  wire h_u_cla24_and3129_y0;
  wire h_u_cla24_and3130_y0;
  wire h_u_cla24_and3131_y0;
  wire h_u_cla24_and3132_y0;
  wire h_u_cla24_and3133_y0;
  wire h_u_cla24_and3134_y0;
  wire h_u_cla24_and3135_y0;
  wire h_u_cla24_and3136_y0;
  wire h_u_cla24_and3137_y0;
  wire h_u_cla24_and3138_y0;
  wire h_u_cla24_and3139_y0;
  wire h_u_cla24_and3140_y0;
  wire h_u_cla24_and3141_y0;
  wire h_u_cla24_and3142_y0;
  wire h_u_cla24_and3143_y0;
  wire h_u_cla24_and3144_y0;
  wire h_u_cla24_and3145_y0;
  wire h_u_cla24_and3146_y0;
  wire h_u_cla24_and3147_y0;
  wire h_u_cla24_and3148_y0;
  wire h_u_cla24_and3149_y0;
  wire h_u_cla24_and3150_y0;
  wire h_u_cla24_and3151_y0;
  wire h_u_cla24_and3152_y0;
  wire h_u_cla24_and3153_y0;
  wire h_u_cla24_and3154_y0;
  wire h_u_cla24_and3155_y0;
  wire h_u_cla24_and3156_y0;
  wire h_u_cla24_and3157_y0;
  wire h_u_cla24_and3158_y0;
  wire h_u_cla24_and3159_y0;
  wire h_u_cla24_and3160_y0;
  wire h_u_cla24_and3161_y0;
  wire h_u_cla24_and3162_y0;
  wire h_u_cla24_and3163_y0;
  wire h_u_cla24_and3164_y0;
  wire h_u_cla24_and3165_y0;
  wire h_u_cla24_and3166_y0;
  wire h_u_cla24_and3167_y0;
  wire h_u_cla24_and3168_y0;
  wire h_u_cla24_and3169_y0;
  wire h_u_cla24_and3170_y0;
  wire h_u_cla24_and3171_y0;
  wire h_u_cla24_and3172_y0;
  wire h_u_cla24_and3173_y0;
  wire h_u_cla24_and3174_y0;
  wire h_u_cla24_and3175_y0;
  wire h_u_cla24_and3176_y0;
  wire h_u_cla24_and3177_y0;
  wire h_u_cla24_and3178_y0;
  wire h_u_cla24_and3179_y0;
  wire h_u_cla24_and3180_y0;
  wire h_u_cla24_and3181_y0;
  wire h_u_cla24_and3182_y0;
  wire h_u_cla24_and3183_y0;
  wire h_u_cla24_and3184_y0;
  wire h_u_cla24_and3185_y0;
  wire h_u_cla24_and3186_y0;
  wire h_u_cla24_and3187_y0;
  wire h_u_cla24_and3188_y0;
  wire h_u_cla24_and3189_y0;
  wire h_u_cla24_and3190_y0;
  wire h_u_cla24_and3191_y0;
  wire h_u_cla24_and3192_y0;
  wire h_u_cla24_and3193_y0;
  wire h_u_cla24_and3194_y0;
  wire h_u_cla24_and3195_y0;
  wire h_u_cla24_and3196_y0;
  wire h_u_cla24_and3197_y0;
  wire h_u_cla24_and3198_y0;
  wire h_u_cla24_and3199_y0;
  wire h_u_cla24_and3200_y0;
  wire h_u_cla24_and3201_y0;
  wire h_u_cla24_and3202_y0;
  wire h_u_cla24_and3203_y0;
  wire h_u_cla24_and3204_y0;
  wire h_u_cla24_and3205_y0;
  wire h_u_cla24_and3206_y0;
  wire h_u_cla24_and3207_y0;
  wire h_u_cla24_and3208_y0;
  wire h_u_cla24_and3209_y0;
  wire h_u_cla24_and3210_y0;
  wire h_u_cla24_and3211_y0;
  wire h_u_cla24_and3212_y0;
  wire h_u_cla24_and3213_y0;
  wire h_u_cla24_and3214_y0;
  wire h_u_cla24_and3215_y0;
  wire h_u_cla24_and3216_y0;
  wire h_u_cla24_and3217_y0;
  wire h_u_cla24_and3218_y0;
  wire h_u_cla24_and3219_y0;
  wire h_u_cla24_and3220_y0;
  wire h_u_cla24_and3221_y0;
  wire h_u_cla24_and3222_y0;
  wire h_u_cla24_and3223_y0;
  wire h_u_cla24_and3224_y0;
  wire h_u_cla24_and3225_y0;
  wire h_u_cla24_and3226_y0;
  wire h_u_cla24_and3227_y0;
  wire h_u_cla24_and3228_y0;
  wire h_u_cla24_and3229_y0;
  wire h_u_cla24_and3230_y0;
  wire h_u_cla24_and3231_y0;
  wire h_u_cla24_and3232_y0;
  wire h_u_cla24_and3233_y0;
  wire h_u_cla24_and3234_y0;
  wire h_u_cla24_and3235_y0;
  wire h_u_cla24_and3236_y0;
  wire h_u_cla24_and3237_y0;
  wire h_u_cla24_and3238_y0;
  wire h_u_cla24_and3239_y0;
  wire h_u_cla24_and3240_y0;
  wire h_u_cla24_and3241_y0;
  wire h_u_cla24_and3242_y0;
  wire h_u_cla24_and3243_y0;
  wire h_u_cla24_and3244_y0;
  wire h_u_cla24_and3245_y0;
  wire h_u_cla24_and3246_y0;
  wire h_u_cla24_and3247_y0;
  wire h_u_cla24_and3248_y0;
  wire h_u_cla24_and3249_y0;
  wire h_u_cla24_and3250_y0;
  wire h_u_cla24_and3251_y0;
  wire h_u_cla24_and3252_y0;
  wire h_u_cla24_and3253_y0;
  wire h_u_cla24_and3254_y0;
  wire h_u_cla24_and3255_y0;
  wire h_u_cla24_and3256_y0;
  wire h_u_cla24_and3257_y0;
  wire h_u_cla24_and3258_y0;
  wire h_u_cla24_and3259_y0;
  wire h_u_cla24_and3260_y0;
  wire h_u_cla24_and3261_y0;
  wire h_u_cla24_and3262_y0;
  wire h_u_cla24_and3263_y0;
  wire h_u_cla24_and3264_y0;
  wire h_u_cla24_and3265_y0;
  wire h_u_cla24_and3266_y0;
  wire h_u_cla24_and3267_y0;
  wire h_u_cla24_and3268_y0;
  wire h_u_cla24_and3269_y0;
  wire h_u_cla24_and3270_y0;
  wire h_u_cla24_and3271_y0;
  wire h_u_cla24_and3272_y0;
  wire h_u_cla24_and3273_y0;
  wire h_u_cla24_and3274_y0;
  wire h_u_cla24_and3275_y0;
  wire h_u_cla24_and3276_y0;
  wire h_u_cla24_and3277_y0;
  wire h_u_cla24_and3278_y0;
  wire h_u_cla24_and3279_y0;
  wire h_u_cla24_and3280_y0;
  wire h_u_cla24_and3281_y0;
  wire h_u_cla24_and3282_y0;
  wire h_u_cla24_and3283_y0;
  wire h_u_cla24_and3284_y0;
  wire h_u_cla24_and3285_y0;
  wire h_u_cla24_and3286_y0;
  wire h_u_cla24_and3287_y0;
  wire h_u_cla24_and3288_y0;
  wire h_u_cla24_and3289_y0;
  wire h_u_cla24_and3290_y0;
  wire h_u_cla24_and3291_y0;
  wire h_u_cla24_and3292_y0;
  wire h_u_cla24_and3293_y0;
  wire h_u_cla24_and3294_y0;
  wire h_u_cla24_and3295_y0;
  wire h_u_cla24_and3296_y0;
  wire h_u_cla24_and3297_y0;
  wire h_u_cla24_and3298_y0;
  wire h_u_cla24_and3299_y0;
  wire h_u_cla24_and3300_y0;
  wire h_u_cla24_and3301_y0;
  wire h_u_cla24_and3302_y0;
  wire h_u_cla24_and3303_y0;
  wire h_u_cla24_and3304_y0;
  wire h_u_cla24_and3305_y0;
  wire h_u_cla24_and3306_y0;
  wire h_u_cla24_and3307_y0;
  wire h_u_cla24_and3308_y0;
  wire h_u_cla24_and3309_y0;
  wire h_u_cla24_and3310_y0;
  wire h_u_cla24_or210_y0;
  wire h_u_cla24_or211_y0;
  wire h_u_cla24_or212_y0;
  wire h_u_cla24_or213_y0;
  wire h_u_cla24_or214_y0;
  wire h_u_cla24_or215_y0;
  wire h_u_cla24_or216_y0;
  wire h_u_cla24_or217_y0;
  wire h_u_cla24_or218_y0;
  wire h_u_cla24_or219_y0;
  wire h_u_cla24_or220_y0;
  wire h_u_cla24_or221_y0;
  wire h_u_cla24_or222_y0;
  wire h_u_cla24_or223_y0;
  wire h_u_cla24_or224_y0;
  wire h_u_cla24_or225_y0;
  wire h_u_cla24_or226_y0;
  wire h_u_cla24_or227_y0;
  wire h_u_cla24_or228_y0;
  wire h_u_cla24_or229_y0;
  wire h_u_cla24_or230_y0;
  wire h_u_cla24_pg_logic21_y0;
  wire h_u_cla24_pg_logic21_y1;
  wire h_u_cla24_pg_logic21_y2;
  wire h_u_cla24_xor21_y0;
  wire h_u_cla24_and3311_y0;
  wire h_u_cla24_and3312_y0;
  wire h_u_cla24_and3313_y0;
  wire h_u_cla24_and3314_y0;
  wire h_u_cla24_and3315_y0;
  wire h_u_cla24_and3316_y0;
  wire h_u_cla24_and3317_y0;
  wire h_u_cla24_and3318_y0;
  wire h_u_cla24_and3319_y0;
  wire h_u_cla24_and3320_y0;
  wire h_u_cla24_and3321_y0;
  wire h_u_cla24_and3322_y0;
  wire h_u_cla24_and3323_y0;
  wire h_u_cla24_and3324_y0;
  wire h_u_cla24_and3325_y0;
  wire h_u_cla24_and3326_y0;
  wire h_u_cla24_and3327_y0;
  wire h_u_cla24_and3328_y0;
  wire h_u_cla24_and3329_y0;
  wire h_u_cla24_and3330_y0;
  wire h_u_cla24_and3331_y0;
  wire h_u_cla24_and3332_y0;
  wire h_u_cla24_and3333_y0;
  wire h_u_cla24_and3334_y0;
  wire h_u_cla24_and3335_y0;
  wire h_u_cla24_and3336_y0;
  wire h_u_cla24_and3337_y0;
  wire h_u_cla24_and3338_y0;
  wire h_u_cla24_and3339_y0;
  wire h_u_cla24_and3340_y0;
  wire h_u_cla24_and3341_y0;
  wire h_u_cla24_and3342_y0;
  wire h_u_cla24_and3343_y0;
  wire h_u_cla24_and3344_y0;
  wire h_u_cla24_and3345_y0;
  wire h_u_cla24_and3346_y0;
  wire h_u_cla24_and3347_y0;
  wire h_u_cla24_and3348_y0;
  wire h_u_cla24_and3349_y0;
  wire h_u_cla24_and3350_y0;
  wire h_u_cla24_and3351_y0;
  wire h_u_cla24_and3352_y0;
  wire h_u_cla24_and3353_y0;
  wire h_u_cla24_and3354_y0;
  wire h_u_cla24_and3355_y0;
  wire h_u_cla24_and3356_y0;
  wire h_u_cla24_and3357_y0;
  wire h_u_cla24_and3358_y0;
  wire h_u_cla24_and3359_y0;
  wire h_u_cla24_and3360_y0;
  wire h_u_cla24_and3361_y0;
  wire h_u_cla24_and3362_y0;
  wire h_u_cla24_and3363_y0;
  wire h_u_cla24_and3364_y0;
  wire h_u_cla24_and3365_y0;
  wire h_u_cla24_and3366_y0;
  wire h_u_cla24_and3367_y0;
  wire h_u_cla24_and3368_y0;
  wire h_u_cla24_and3369_y0;
  wire h_u_cla24_and3370_y0;
  wire h_u_cla24_and3371_y0;
  wire h_u_cla24_and3372_y0;
  wire h_u_cla24_and3373_y0;
  wire h_u_cla24_and3374_y0;
  wire h_u_cla24_and3375_y0;
  wire h_u_cla24_and3376_y0;
  wire h_u_cla24_and3377_y0;
  wire h_u_cla24_and3378_y0;
  wire h_u_cla24_and3379_y0;
  wire h_u_cla24_and3380_y0;
  wire h_u_cla24_and3381_y0;
  wire h_u_cla24_and3382_y0;
  wire h_u_cla24_and3383_y0;
  wire h_u_cla24_and3384_y0;
  wire h_u_cla24_and3385_y0;
  wire h_u_cla24_and3386_y0;
  wire h_u_cla24_and3387_y0;
  wire h_u_cla24_and3388_y0;
  wire h_u_cla24_and3389_y0;
  wire h_u_cla24_and3390_y0;
  wire h_u_cla24_and3391_y0;
  wire h_u_cla24_and3392_y0;
  wire h_u_cla24_and3393_y0;
  wire h_u_cla24_and3394_y0;
  wire h_u_cla24_and3395_y0;
  wire h_u_cla24_and3396_y0;
  wire h_u_cla24_and3397_y0;
  wire h_u_cla24_and3398_y0;
  wire h_u_cla24_and3399_y0;
  wire h_u_cla24_and3400_y0;
  wire h_u_cla24_and3401_y0;
  wire h_u_cla24_and3402_y0;
  wire h_u_cla24_and3403_y0;
  wire h_u_cla24_and3404_y0;
  wire h_u_cla24_and3405_y0;
  wire h_u_cla24_and3406_y0;
  wire h_u_cla24_and3407_y0;
  wire h_u_cla24_and3408_y0;
  wire h_u_cla24_and3409_y0;
  wire h_u_cla24_and3410_y0;
  wire h_u_cla24_and3411_y0;
  wire h_u_cla24_and3412_y0;
  wire h_u_cla24_and3413_y0;
  wire h_u_cla24_and3414_y0;
  wire h_u_cla24_and3415_y0;
  wire h_u_cla24_and3416_y0;
  wire h_u_cla24_and3417_y0;
  wire h_u_cla24_and3418_y0;
  wire h_u_cla24_and3419_y0;
  wire h_u_cla24_and3420_y0;
  wire h_u_cla24_and3421_y0;
  wire h_u_cla24_and3422_y0;
  wire h_u_cla24_and3423_y0;
  wire h_u_cla24_and3424_y0;
  wire h_u_cla24_and3425_y0;
  wire h_u_cla24_and3426_y0;
  wire h_u_cla24_and3427_y0;
  wire h_u_cla24_and3428_y0;
  wire h_u_cla24_and3429_y0;
  wire h_u_cla24_and3430_y0;
  wire h_u_cla24_and3431_y0;
  wire h_u_cla24_and3432_y0;
  wire h_u_cla24_and3433_y0;
  wire h_u_cla24_and3434_y0;
  wire h_u_cla24_and3435_y0;
  wire h_u_cla24_and3436_y0;
  wire h_u_cla24_and3437_y0;
  wire h_u_cla24_and3438_y0;
  wire h_u_cla24_and3439_y0;
  wire h_u_cla24_and3440_y0;
  wire h_u_cla24_and3441_y0;
  wire h_u_cla24_and3442_y0;
  wire h_u_cla24_and3443_y0;
  wire h_u_cla24_and3444_y0;
  wire h_u_cla24_and3445_y0;
  wire h_u_cla24_and3446_y0;
  wire h_u_cla24_and3447_y0;
  wire h_u_cla24_and3448_y0;
  wire h_u_cla24_and3449_y0;
  wire h_u_cla24_and3450_y0;
  wire h_u_cla24_and3451_y0;
  wire h_u_cla24_and3452_y0;
  wire h_u_cla24_and3453_y0;
  wire h_u_cla24_and3454_y0;
  wire h_u_cla24_and3455_y0;
  wire h_u_cla24_and3456_y0;
  wire h_u_cla24_and3457_y0;
  wire h_u_cla24_and3458_y0;
  wire h_u_cla24_and3459_y0;
  wire h_u_cla24_and3460_y0;
  wire h_u_cla24_and3461_y0;
  wire h_u_cla24_and3462_y0;
  wire h_u_cla24_and3463_y0;
  wire h_u_cla24_and3464_y0;
  wire h_u_cla24_and3465_y0;
  wire h_u_cla24_and3466_y0;
  wire h_u_cla24_and3467_y0;
  wire h_u_cla24_and3468_y0;
  wire h_u_cla24_and3469_y0;
  wire h_u_cla24_and3470_y0;
  wire h_u_cla24_and3471_y0;
  wire h_u_cla24_and3472_y0;
  wire h_u_cla24_and3473_y0;
  wire h_u_cla24_and3474_y0;
  wire h_u_cla24_and3475_y0;
  wire h_u_cla24_and3476_y0;
  wire h_u_cla24_and3477_y0;
  wire h_u_cla24_and3478_y0;
  wire h_u_cla24_and3479_y0;
  wire h_u_cla24_and3480_y0;
  wire h_u_cla24_and3481_y0;
  wire h_u_cla24_and3482_y0;
  wire h_u_cla24_and3483_y0;
  wire h_u_cla24_and3484_y0;
  wire h_u_cla24_and3485_y0;
  wire h_u_cla24_and3486_y0;
  wire h_u_cla24_and3487_y0;
  wire h_u_cla24_and3488_y0;
  wire h_u_cla24_and3489_y0;
  wire h_u_cla24_and3490_y0;
  wire h_u_cla24_and3491_y0;
  wire h_u_cla24_and3492_y0;
  wire h_u_cla24_and3493_y0;
  wire h_u_cla24_and3494_y0;
  wire h_u_cla24_and3495_y0;
  wire h_u_cla24_and3496_y0;
  wire h_u_cla24_and3497_y0;
  wire h_u_cla24_and3498_y0;
  wire h_u_cla24_and3499_y0;
  wire h_u_cla24_and3500_y0;
  wire h_u_cla24_and3501_y0;
  wire h_u_cla24_and3502_y0;
  wire h_u_cla24_and3503_y0;
  wire h_u_cla24_and3504_y0;
  wire h_u_cla24_and3505_y0;
  wire h_u_cla24_and3506_y0;
  wire h_u_cla24_and3507_y0;
  wire h_u_cla24_and3508_y0;
  wire h_u_cla24_and3509_y0;
  wire h_u_cla24_and3510_y0;
  wire h_u_cla24_and3511_y0;
  wire h_u_cla24_and3512_y0;
  wire h_u_cla24_and3513_y0;
  wire h_u_cla24_and3514_y0;
  wire h_u_cla24_and3515_y0;
  wire h_u_cla24_and3516_y0;
  wire h_u_cla24_and3517_y0;
  wire h_u_cla24_and3518_y0;
  wire h_u_cla24_and3519_y0;
  wire h_u_cla24_and3520_y0;
  wire h_u_cla24_and3521_y0;
  wire h_u_cla24_and3522_y0;
  wire h_u_cla24_and3523_y0;
  wire h_u_cla24_and3524_y0;
  wire h_u_cla24_and3525_y0;
  wire h_u_cla24_and3526_y0;
  wire h_u_cla24_and3527_y0;
  wire h_u_cla24_and3528_y0;
  wire h_u_cla24_and3529_y0;
  wire h_u_cla24_and3530_y0;
  wire h_u_cla24_and3531_y0;
  wire h_u_cla24_and3532_y0;
  wire h_u_cla24_and3533_y0;
  wire h_u_cla24_and3534_y0;
  wire h_u_cla24_and3535_y0;
  wire h_u_cla24_and3536_y0;
  wire h_u_cla24_and3537_y0;
  wire h_u_cla24_and3538_y0;
  wire h_u_cla24_and3539_y0;
  wire h_u_cla24_and3540_y0;
  wire h_u_cla24_and3541_y0;
  wire h_u_cla24_and3542_y0;
  wire h_u_cla24_and3543_y0;
  wire h_u_cla24_and3544_y0;
  wire h_u_cla24_and3545_y0;
  wire h_u_cla24_and3546_y0;
  wire h_u_cla24_and3547_y0;
  wire h_u_cla24_and3548_y0;
  wire h_u_cla24_and3549_y0;
  wire h_u_cla24_and3550_y0;
  wire h_u_cla24_and3551_y0;
  wire h_u_cla24_and3552_y0;
  wire h_u_cla24_and3553_y0;
  wire h_u_cla24_and3554_y0;
  wire h_u_cla24_and3555_y0;
  wire h_u_cla24_and3556_y0;
  wire h_u_cla24_and3557_y0;
  wire h_u_cla24_and3558_y0;
  wire h_u_cla24_and3559_y0;
  wire h_u_cla24_and3560_y0;
  wire h_u_cla24_and3561_y0;
  wire h_u_cla24_and3562_y0;
  wire h_u_cla24_and3563_y0;
  wire h_u_cla24_and3564_y0;
  wire h_u_cla24_and3565_y0;
  wire h_u_cla24_and3566_y0;
  wire h_u_cla24_and3567_y0;
  wire h_u_cla24_and3568_y0;
  wire h_u_cla24_and3569_y0;
  wire h_u_cla24_and3570_y0;
  wire h_u_cla24_and3571_y0;
  wire h_u_cla24_and3572_y0;
  wire h_u_cla24_and3573_y0;
  wire h_u_cla24_and3574_y0;
  wire h_u_cla24_and3575_y0;
  wire h_u_cla24_and3576_y0;
  wire h_u_cla24_and3577_y0;
  wire h_u_cla24_and3578_y0;
  wire h_u_cla24_and3579_y0;
  wire h_u_cla24_and3580_y0;
  wire h_u_cla24_and3581_y0;
  wire h_u_cla24_and3582_y0;
  wire h_u_cla24_and3583_y0;
  wire h_u_cla24_and3584_y0;
  wire h_u_cla24_and3585_y0;
  wire h_u_cla24_and3586_y0;
  wire h_u_cla24_and3587_y0;
  wire h_u_cla24_and3588_y0;
  wire h_u_cla24_and3589_y0;
  wire h_u_cla24_and3590_y0;
  wire h_u_cla24_and3591_y0;
  wire h_u_cla24_and3592_y0;
  wire h_u_cla24_and3593_y0;
  wire h_u_cla24_and3594_y0;
  wire h_u_cla24_and3595_y0;
  wire h_u_cla24_and3596_y0;
  wire h_u_cla24_and3597_y0;
  wire h_u_cla24_and3598_y0;
  wire h_u_cla24_and3599_y0;
  wire h_u_cla24_and3600_y0;
  wire h_u_cla24_and3601_y0;
  wire h_u_cla24_and3602_y0;
  wire h_u_cla24_and3603_y0;
  wire h_u_cla24_and3604_y0;
  wire h_u_cla24_and3605_y0;
  wire h_u_cla24_and3606_y0;
  wire h_u_cla24_and3607_y0;
  wire h_u_cla24_and3608_y0;
  wire h_u_cla24_and3609_y0;
  wire h_u_cla24_and3610_y0;
  wire h_u_cla24_and3611_y0;
  wire h_u_cla24_and3612_y0;
  wire h_u_cla24_and3613_y0;
  wire h_u_cla24_and3614_y0;
  wire h_u_cla24_and3615_y0;
  wire h_u_cla24_and3616_y0;
  wire h_u_cla24_and3617_y0;
  wire h_u_cla24_and3618_y0;
  wire h_u_cla24_and3619_y0;
  wire h_u_cla24_and3620_y0;
  wire h_u_cla24_and3621_y0;
  wire h_u_cla24_and3622_y0;
  wire h_u_cla24_and3623_y0;
  wire h_u_cla24_and3624_y0;
  wire h_u_cla24_and3625_y0;
  wire h_u_cla24_and3626_y0;
  wire h_u_cla24_and3627_y0;
  wire h_u_cla24_and3628_y0;
  wire h_u_cla24_and3629_y0;
  wire h_u_cla24_and3630_y0;
  wire h_u_cla24_and3631_y0;
  wire h_u_cla24_and3632_y0;
  wire h_u_cla24_and3633_y0;
  wire h_u_cla24_and3634_y0;
  wire h_u_cla24_and3635_y0;
  wire h_u_cla24_and3636_y0;
  wire h_u_cla24_and3637_y0;
  wire h_u_cla24_and3638_y0;
  wire h_u_cla24_and3639_y0;
  wire h_u_cla24_and3640_y0;
  wire h_u_cla24_and3641_y0;
  wire h_u_cla24_and3642_y0;
  wire h_u_cla24_and3643_y0;
  wire h_u_cla24_and3644_y0;
  wire h_u_cla24_and3645_y0;
  wire h_u_cla24_and3646_y0;
  wire h_u_cla24_and3647_y0;
  wire h_u_cla24_and3648_y0;
  wire h_u_cla24_and3649_y0;
  wire h_u_cla24_and3650_y0;
  wire h_u_cla24_and3651_y0;
  wire h_u_cla24_and3652_y0;
  wire h_u_cla24_and3653_y0;
  wire h_u_cla24_and3654_y0;
  wire h_u_cla24_and3655_y0;
  wire h_u_cla24_and3656_y0;
  wire h_u_cla24_and3657_y0;
  wire h_u_cla24_and3658_y0;
  wire h_u_cla24_and3659_y0;
  wire h_u_cla24_and3660_y0;
  wire h_u_cla24_and3661_y0;
  wire h_u_cla24_and3662_y0;
  wire h_u_cla24_and3663_y0;
  wire h_u_cla24_and3664_y0;
  wire h_u_cla24_and3665_y0;
  wire h_u_cla24_and3666_y0;
  wire h_u_cla24_and3667_y0;
  wire h_u_cla24_and3668_y0;
  wire h_u_cla24_and3669_y0;
  wire h_u_cla24_and3670_y0;
  wire h_u_cla24_and3671_y0;
  wire h_u_cla24_and3672_y0;
  wire h_u_cla24_and3673_y0;
  wire h_u_cla24_and3674_y0;
  wire h_u_cla24_and3675_y0;
  wire h_u_cla24_and3676_y0;
  wire h_u_cla24_and3677_y0;
  wire h_u_cla24_and3678_y0;
  wire h_u_cla24_and3679_y0;
  wire h_u_cla24_and3680_y0;
  wire h_u_cla24_and3681_y0;
  wire h_u_cla24_and3682_y0;
  wire h_u_cla24_and3683_y0;
  wire h_u_cla24_and3684_y0;
  wire h_u_cla24_and3685_y0;
  wire h_u_cla24_and3686_y0;
  wire h_u_cla24_and3687_y0;
  wire h_u_cla24_and3688_y0;
  wire h_u_cla24_and3689_y0;
  wire h_u_cla24_and3690_y0;
  wire h_u_cla24_and3691_y0;
  wire h_u_cla24_and3692_y0;
  wire h_u_cla24_and3693_y0;
  wire h_u_cla24_and3694_y0;
  wire h_u_cla24_and3695_y0;
  wire h_u_cla24_and3696_y0;
  wire h_u_cla24_and3697_y0;
  wire h_u_cla24_and3698_y0;
  wire h_u_cla24_and3699_y0;
  wire h_u_cla24_and3700_y0;
  wire h_u_cla24_and3701_y0;
  wire h_u_cla24_and3702_y0;
  wire h_u_cla24_and3703_y0;
  wire h_u_cla24_and3704_y0;
  wire h_u_cla24_and3705_y0;
  wire h_u_cla24_and3706_y0;
  wire h_u_cla24_and3707_y0;
  wire h_u_cla24_and3708_y0;
  wire h_u_cla24_and3709_y0;
  wire h_u_cla24_and3710_y0;
  wire h_u_cla24_and3711_y0;
  wire h_u_cla24_and3712_y0;
  wire h_u_cla24_and3713_y0;
  wire h_u_cla24_and3714_y0;
  wire h_u_cla24_and3715_y0;
  wire h_u_cla24_and3716_y0;
  wire h_u_cla24_and3717_y0;
  wire h_u_cla24_and3718_y0;
  wire h_u_cla24_and3719_y0;
  wire h_u_cla24_and3720_y0;
  wire h_u_cla24_and3721_y0;
  wire h_u_cla24_and3722_y0;
  wire h_u_cla24_and3723_y0;
  wire h_u_cla24_and3724_y0;
  wire h_u_cla24_and3725_y0;
  wire h_u_cla24_and3726_y0;
  wire h_u_cla24_and3727_y0;
  wire h_u_cla24_and3728_y0;
  wire h_u_cla24_and3729_y0;
  wire h_u_cla24_and3730_y0;
  wire h_u_cla24_and3731_y0;
  wire h_u_cla24_and3732_y0;
  wire h_u_cla24_and3733_y0;
  wire h_u_cla24_and3734_y0;
  wire h_u_cla24_and3735_y0;
  wire h_u_cla24_and3736_y0;
  wire h_u_cla24_and3737_y0;
  wire h_u_cla24_and3738_y0;
  wire h_u_cla24_and3739_y0;
  wire h_u_cla24_and3740_y0;
  wire h_u_cla24_and3741_y0;
  wire h_u_cla24_and3742_y0;
  wire h_u_cla24_and3743_y0;
  wire h_u_cla24_and3744_y0;
  wire h_u_cla24_and3745_y0;
  wire h_u_cla24_and3746_y0;
  wire h_u_cla24_and3747_y0;
  wire h_u_cla24_and3748_y0;
  wire h_u_cla24_and3749_y0;
  wire h_u_cla24_and3750_y0;
  wire h_u_cla24_and3751_y0;
  wire h_u_cla24_and3752_y0;
  wire h_u_cla24_and3753_y0;
  wire h_u_cla24_and3754_y0;
  wire h_u_cla24_and3755_y0;
  wire h_u_cla24_and3756_y0;
  wire h_u_cla24_and3757_y0;
  wire h_u_cla24_and3758_y0;
  wire h_u_cla24_and3759_y0;
  wire h_u_cla24_and3760_y0;
  wire h_u_cla24_and3761_y0;
  wire h_u_cla24_and3762_y0;
  wire h_u_cla24_and3763_y0;
  wire h_u_cla24_and3764_y0;
  wire h_u_cla24_and3765_y0;
  wire h_u_cla24_and3766_y0;
  wire h_u_cla24_and3767_y0;
  wire h_u_cla24_and3768_y0;
  wire h_u_cla24_and3769_y0;
  wire h_u_cla24_and3770_y0;
  wire h_u_cla24_and3771_y0;
  wire h_u_cla24_and3772_y0;
  wire h_u_cla24_and3773_y0;
  wire h_u_cla24_and3774_y0;
  wire h_u_cla24_and3775_y0;
  wire h_u_cla24_and3776_y0;
  wire h_u_cla24_and3777_y0;
  wire h_u_cla24_and3778_y0;
  wire h_u_cla24_and3779_y0;
  wire h_u_cla24_and3780_y0;
  wire h_u_cla24_and3781_y0;
  wire h_u_cla24_and3782_y0;
  wire h_u_cla24_and3783_y0;
  wire h_u_cla24_and3784_y0;
  wire h_u_cla24_and3785_y0;
  wire h_u_cla24_and3786_y0;
  wire h_u_cla24_and3787_y0;
  wire h_u_cla24_and3788_y0;
  wire h_u_cla24_and3789_y0;
  wire h_u_cla24_and3790_y0;
  wire h_u_cla24_and3791_y0;
  wire h_u_cla24_and3792_y0;
  wire h_u_cla24_and3793_y0;
  wire h_u_cla24_and3794_y0;
  wire h_u_cla24_or231_y0;
  wire h_u_cla24_or232_y0;
  wire h_u_cla24_or233_y0;
  wire h_u_cla24_or234_y0;
  wire h_u_cla24_or235_y0;
  wire h_u_cla24_or236_y0;
  wire h_u_cla24_or237_y0;
  wire h_u_cla24_or238_y0;
  wire h_u_cla24_or239_y0;
  wire h_u_cla24_or240_y0;
  wire h_u_cla24_or241_y0;
  wire h_u_cla24_or242_y0;
  wire h_u_cla24_or243_y0;
  wire h_u_cla24_or244_y0;
  wire h_u_cla24_or245_y0;
  wire h_u_cla24_or246_y0;
  wire h_u_cla24_or247_y0;
  wire h_u_cla24_or248_y0;
  wire h_u_cla24_or249_y0;
  wire h_u_cla24_or250_y0;
  wire h_u_cla24_or251_y0;
  wire h_u_cla24_or252_y0;
  wire h_u_cla24_pg_logic22_y0;
  wire h_u_cla24_pg_logic22_y1;
  wire h_u_cla24_pg_logic22_y2;
  wire h_u_cla24_xor22_y0;
  wire h_u_cla24_and3795_y0;
  wire h_u_cla24_and3796_y0;
  wire h_u_cla24_and3797_y0;
  wire h_u_cla24_and3798_y0;
  wire h_u_cla24_and3799_y0;
  wire h_u_cla24_and3800_y0;
  wire h_u_cla24_and3801_y0;
  wire h_u_cla24_and3802_y0;
  wire h_u_cla24_and3803_y0;
  wire h_u_cla24_and3804_y0;
  wire h_u_cla24_and3805_y0;
  wire h_u_cla24_and3806_y0;
  wire h_u_cla24_and3807_y0;
  wire h_u_cla24_and3808_y0;
  wire h_u_cla24_and3809_y0;
  wire h_u_cla24_and3810_y0;
  wire h_u_cla24_and3811_y0;
  wire h_u_cla24_and3812_y0;
  wire h_u_cla24_and3813_y0;
  wire h_u_cla24_and3814_y0;
  wire h_u_cla24_and3815_y0;
  wire h_u_cla24_and3816_y0;
  wire h_u_cla24_and3817_y0;
  wire h_u_cla24_and3818_y0;
  wire h_u_cla24_and3819_y0;
  wire h_u_cla24_and3820_y0;
  wire h_u_cla24_and3821_y0;
  wire h_u_cla24_and3822_y0;
  wire h_u_cla24_and3823_y0;
  wire h_u_cla24_and3824_y0;
  wire h_u_cla24_and3825_y0;
  wire h_u_cla24_and3826_y0;
  wire h_u_cla24_and3827_y0;
  wire h_u_cla24_and3828_y0;
  wire h_u_cla24_and3829_y0;
  wire h_u_cla24_and3830_y0;
  wire h_u_cla24_and3831_y0;
  wire h_u_cla24_and3832_y0;
  wire h_u_cla24_and3833_y0;
  wire h_u_cla24_and3834_y0;
  wire h_u_cla24_and3835_y0;
  wire h_u_cla24_and3836_y0;
  wire h_u_cla24_and3837_y0;
  wire h_u_cla24_and3838_y0;
  wire h_u_cla24_and3839_y0;
  wire h_u_cla24_and3840_y0;
  wire h_u_cla24_and3841_y0;
  wire h_u_cla24_and3842_y0;
  wire h_u_cla24_and3843_y0;
  wire h_u_cla24_and3844_y0;
  wire h_u_cla24_and3845_y0;
  wire h_u_cla24_and3846_y0;
  wire h_u_cla24_and3847_y0;
  wire h_u_cla24_and3848_y0;
  wire h_u_cla24_and3849_y0;
  wire h_u_cla24_and3850_y0;
  wire h_u_cla24_and3851_y0;
  wire h_u_cla24_and3852_y0;
  wire h_u_cla24_and3853_y0;
  wire h_u_cla24_and3854_y0;
  wire h_u_cla24_and3855_y0;
  wire h_u_cla24_and3856_y0;
  wire h_u_cla24_and3857_y0;
  wire h_u_cla24_and3858_y0;
  wire h_u_cla24_and3859_y0;
  wire h_u_cla24_and3860_y0;
  wire h_u_cla24_and3861_y0;
  wire h_u_cla24_and3862_y0;
  wire h_u_cla24_and3863_y0;
  wire h_u_cla24_and3864_y0;
  wire h_u_cla24_and3865_y0;
  wire h_u_cla24_and3866_y0;
  wire h_u_cla24_and3867_y0;
  wire h_u_cla24_and3868_y0;
  wire h_u_cla24_and3869_y0;
  wire h_u_cla24_and3870_y0;
  wire h_u_cla24_and3871_y0;
  wire h_u_cla24_and3872_y0;
  wire h_u_cla24_and3873_y0;
  wire h_u_cla24_and3874_y0;
  wire h_u_cla24_and3875_y0;
  wire h_u_cla24_and3876_y0;
  wire h_u_cla24_and3877_y0;
  wire h_u_cla24_and3878_y0;
  wire h_u_cla24_and3879_y0;
  wire h_u_cla24_and3880_y0;
  wire h_u_cla24_and3881_y0;
  wire h_u_cla24_and3882_y0;
  wire h_u_cla24_and3883_y0;
  wire h_u_cla24_and3884_y0;
  wire h_u_cla24_and3885_y0;
  wire h_u_cla24_and3886_y0;
  wire h_u_cla24_and3887_y0;
  wire h_u_cla24_and3888_y0;
  wire h_u_cla24_and3889_y0;
  wire h_u_cla24_and3890_y0;
  wire h_u_cla24_and3891_y0;
  wire h_u_cla24_and3892_y0;
  wire h_u_cla24_and3893_y0;
  wire h_u_cla24_and3894_y0;
  wire h_u_cla24_and3895_y0;
  wire h_u_cla24_and3896_y0;
  wire h_u_cla24_and3897_y0;
  wire h_u_cla24_and3898_y0;
  wire h_u_cla24_and3899_y0;
  wire h_u_cla24_and3900_y0;
  wire h_u_cla24_and3901_y0;
  wire h_u_cla24_and3902_y0;
  wire h_u_cla24_and3903_y0;
  wire h_u_cla24_and3904_y0;
  wire h_u_cla24_and3905_y0;
  wire h_u_cla24_and3906_y0;
  wire h_u_cla24_and3907_y0;
  wire h_u_cla24_and3908_y0;
  wire h_u_cla24_and3909_y0;
  wire h_u_cla24_and3910_y0;
  wire h_u_cla24_and3911_y0;
  wire h_u_cla24_and3912_y0;
  wire h_u_cla24_and3913_y0;
  wire h_u_cla24_and3914_y0;
  wire h_u_cla24_and3915_y0;
  wire h_u_cla24_and3916_y0;
  wire h_u_cla24_and3917_y0;
  wire h_u_cla24_and3918_y0;
  wire h_u_cla24_and3919_y0;
  wire h_u_cla24_and3920_y0;
  wire h_u_cla24_and3921_y0;
  wire h_u_cla24_and3922_y0;
  wire h_u_cla24_and3923_y0;
  wire h_u_cla24_and3924_y0;
  wire h_u_cla24_and3925_y0;
  wire h_u_cla24_and3926_y0;
  wire h_u_cla24_and3927_y0;
  wire h_u_cla24_and3928_y0;
  wire h_u_cla24_and3929_y0;
  wire h_u_cla24_and3930_y0;
  wire h_u_cla24_and3931_y0;
  wire h_u_cla24_and3932_y0;
  wire h_u_cla24_and3933_y0;
  wire h_u_cla24_and3934_y0;
  wire h_u_cla24_and3935_y0;
  wire h_u_cla24_and3936_y0;
  wire h_u_cla24_and3937_y0;
  wire h_u_cla24_and3938_y0;
  wire h_u_cla24_and3939_y0;
  wire h_u_cla24_and3940_y0;
  wire h_u_cla24_and3941_y0;
  wire h_u_cla24_and3942_y0;
  wire h_u_cla24_and3943_y0;
  wire h_u_cla24_and3944_y0;
  wire h_u_cla24_and3945_y0;
  wire h_u_cla24_and3946_y0;
  wire h_u_cla24_and3947_y0;
  wire h_u_cla24_and3948_y0;
  wire h_u_cla24_and3949_y0;
  wire h_u_cla24_and3950_y0;
  wire h_u_cla24_and3951_y0;
  wire h_u_cla24_and3952_y0;
  wire h_u_cla24_and3953_y0;
  wire h_u_cla24_and3954_y0;
  wire h_u_cla24_and3955_y0;
  wire h_u_cla24_and3956_y0;
  wire h_u_cla24_and3957_y0;
  wire h_u_cla24_and3958_y0;
  wire h_u_cla24_and3959_y0;
  wire h_u_cla24_and3960_y0;
  wire h_u_cla24_and3961_y0;
  wire h_u_cla24_and3962_y0;
  wire h_u_cla24_and3963_y0;
  wire h_u_cla24_and3964_y0;
  wire h_u_cla24_and3965_y0;
  wire h_u_cla24_and3966_y0;
  wire h_u_cla24_and3967_y0;
  wire h_u_cla24_and3968_y0;
  wire h_u_cla24_and3969_y0;
  wire h_u_cla24_and3970_y0;
  wire h_u_cla24_and3971_y0;
  wire h_u_cla24_and3972_y0;
  wire h_u_cla24_and3973_y0;
  wire h_u_cla24_and3974_y0;
  wire h_u_cla24_and3975_y0;
  wire h_u_cla24_and3976_y0;
  wire h_u_cla24_and3977_y0;
  wire h_u_cla24_and3978_y0;
  wire h_u_cla24_and3979_y0;
  wire h_u_cla24_and3980_y0;
  wire h_u_cla24_and3981_y0;
  wire h_u_cla24_and3982_y0;
  wire h_u_cla24_and3983_y0;
  wire h_u_cla24_and3984_y0;
  wire h_u_cla24_and3985_y0;
  wire h_u_cla24_and3986_y0;
  wire h_u_cla24_and3987_y0;
  wire h_u_cla24_and3988_y0;
  wire h_u_cla24_and3989_y0;
  wire h_u_cla24_and3990_y0;
  wire h_u_cla24_and3991_y0;
  wire h_u_cla24_and3992_y0;
  wire h_u_cla24_and3993_y0;
  wire h_u_cla24_and3994_y0;
  wire h_u_cla24_and3995_y0;
  wire h_u_cla24_and3996_y0;
  wire h_u_cla24_and3997_y0;
  wire h_u_cla24_and3998_y0;
  wire h_u_cla24_and3999_y0;
  wire h_u_cla24_and4000_y0;
  wire h_u_cla24_and4001_y0;
  wire h_u_cla24_and4002_y0;
  wire h_u_cla24_and4003_y0;
  wire h_u_cla24_and4004_y0;
  wire h_u_cla24_and4005_y0;
  wire h_u_cla24_and4006_y0;
  wire h_u_cla24_and4007_y0;
  wire h_u_cla24_and4008_y0;
  wire h_u_cla24_and4009_y0;
  wire h_u_cla24_and4010_y0;
  wire h_u_cla24_and4011_y0;
  wire h_u_cla24_and4012_y0;
  wire h_u_cla24_and4013_y0;
  wire h_u_cla24_and4014_y0;
  wire h_u_cla24_and4015_y0;
  wire h_u_cla24_and4016_y0;
  wire h_u_cla24_and4017_y0;
  wire h_u_cla24_and4018_y0;
  wire h_u_cla24_and4019_y0;
  wire h_u_cla24_and4020_y0;
  wire h_u_cla24_and4021_y0;
  wire h_u_cla24_and4022_y0;
  wire h_u_cla24_and4023_y0;
  wire h_u_cla24_and4024_y0;
  wire h_u_cla24_and4025_y0;
  wire h_u_cla24_and4026_y0;
  wire h_u_cla24_and4027_y0;
  wire h_u_cla24_and4028_y0;
  wire h_u_cla24_and4029_y0;
  wire h_u_cla24_and4030_y0;
  wire h_u_cla24_and4031_y0;
  wire h_u_cla24_and4032_y0;
  wire h_u_cla24_and4033_y0;
  wire h_u_cla24_and4034_y0;
  wire h_u_cla24_and4035_y0;
  wire h_u_cla24_and4036_y0;
  wire h_u_cla24_and4037_y0;
  wire h_u_cla24_and4038_y0;
  wire h_u_cla24_and4039_y0;
  wire h_u_cla24_and4040_y0;
  wire h_u_cla24_and4041_y0;
  wire h_u_cla24_and4042_y0;
  wire h_u_cla24_and4043_y0;
  wire h_u_cla24_and4044_y0;
  wire h_u_cla24_and4045_y0;
  wire h_u_cla24_and4046_y0;
  wire h_u_cla24_and4047_y0;
  wire h_u_cla24_and4048_y0;
  wire h_u_cla24_and4049_y0;
  wire h_u_cla24_and4050_y0;
  wire h_u_cla24_and4051_y0;
  wire h_u_cla24_and4052_y0;
  wire h_u_cla24_and4053_y0;
  wire h_u_cla24_and4054_y0;
  wire h_u_cla24_and4055_y0;
  wire h_u_cla24_and4056_y0;
  wire h_u_cla24_and4057_y0;
  wire h_u_cla24_and4058_y0;
  wire h_u_cla24_and4059_y0;
  wire h_u_cla24_and4060_y0;
  wire h_u_cla24_and4061_y0;
  wire h_u_cla24_and4062_y0;
  wire h_u_cla24_and4063_y0;
  wire h_u_cla24_and4064_y0;
  wire h_u_cla24_and4065_y0;
  wire h_u_cla24_and4066_y0;
  wire h_u_cla24_and4067_y0;
  wire h_u_cla24_and4068_y0;
  wire h_u_cla24_and4069_y0;
  wire h_u_cla24_and4070_y0;
  wire h_u_cla24_and4071_y0;
  wire h_u_cla24_and4072_y0;
  wire h_u_cla24_and4073_y0;
  wire h_u_cla24_and4074_y0;
  wire h_u_cla24_and4075_y0;
  wire h_u_cla24_and4076_y0;
  wire h_u_cla24_and4077_y0;
  wire h_u_cla24_and4078_y0;
  wire h_u_cla24_and4079_y0;
  wire h_u_cla24_and4080_y0;
  wire h_u_cla24_and4081_y0;
  wire h_u_cla24_and4082_y0;
  wire h_u_cla24_and4083_y0;
  wire h_u_cla24_and4084_y0;
  wire h_u_cla24_and4085_y0;
  wire h_u_cla24_and4086_y0;
  wire h_u_cla24_and4087_y0;
  wire h_u_cla24_and4088_y0;
  wire h_u_cla24_and4089_y0;
  wire h_u_cla24_and4090_y0;
  wire h_u_cla24_and4091_y0;
  wire h_u_cla24_and4092_y0;
  wire h_u_cla24_and4093_y0;
  wire h_u_cla24_and4094_y0;
  wire h_u_cla24_and4095_y0;
  wire h_u_cla24_and4096_y0;
  wire h_u_cla24_and4097_y0;
  wire h_u_cla24_and4098_y0;
  wire h_u_cla24_and4099_y0;
  wire h_u_cla24_and4100_y0;
  wire h_u_cla24_and4101_y0;
  wire h_u_cla24_and4102_y0;
  wire h_u_cla24_and4103_y0;
  wire h_u_cla24_and4104_y0;
  wire h_u_cla24_and4105_y0;
  wire h_u_cla24_and4106_y0;
  wire h_u_cla24_and4107_y0;
  wire h_u_cla24_and4108_y0;
  wire h_u_cla24_and4109_y0;
  wire h_u_cla24_and4110_y0;
  wire h_u_cla24_and4111_y0;
  wire h_u_cla24_and4112_y0;
  wire h_u_cla24_and4113_y0;
  wire h_u_cla24_and4114_y0;
  wire h_u_cla24_and4115_y0;
  wire h_u_cla24_and4116_y0;
  wire h_u_cla24_and4117_y0;
  wire h_u_cla24_and4118_y0;
  wire h_u_cla24_and4119_y0;
  wire h_u_cla24_and4120_y0;
  wire h_u_cla24_and4121_y0;
  wire h_u_cla24_and4122_y0;
  wire h_u_cla24_and4123_y0;
  wire h_u_cla24_and4124_y0;
  wire h_u_cla24_and4125_y0;
  wire h_u_cla24_and4126_y0;
  wire h_u_cla24_and4127_y0;
  wire h_u_cla24_and4128_y0;
  wire h_u_cla24_and4129_y0;
  wire h_u_cla24_and4130_y0;
  wire h_u_cla24_and4131_y0;
  wire h_u_cla24_and4132_y0;
  wire h_u_cla24_and4133_y0;
  wire h_u_cla24_and4134_y0;
  wire h_u_cla24_and4135_y0;
  wire h_u_cla24_and4136_y0;
  wire h_u_cla24_and4137_y0;
  wire h_u_cla24_and4138_y0;
  wire h_u_cla24_and4139_y0;
  wire h_u_cla24_and4140_y0;
  wire h_u_cla24_and4141_y0;
  wire h_u_cla24_and4142_y0;
  wire h_u_cla24_and4143_y0;
  wire h_u_cla24_and4144_y0;
  wire h_u_cla24_and4145_y0;
  wire h_u_cla24_and4146_y0;
  wire h_u_cla24_and4147_y0;
  wire h_u_cla24_and4148_y0;
  wire h_u_cla24_and4149_y0;
  wire h_u_cla24_and4150_y0;
  wire h_u_cla24_and4151_y0;
  wire h_u_cla24_and4152_y0;
  wire h_u_cla24_and4153_y0;
  wire h_u_cla24_and4154_y0;
  wire h_u_cla24_and4155_y0;
  wire h_u_cla24_and4156_y0;
  wire h_u_cla24_and4157_y0;
  wire h_u_cla24_and4158_y0;
  wire h_u_cla24_and4159_y0;
  wire h_u_cla24_and4160_y0;
  wire h_u_cla24_and4161_y0;
  wire h_u_cla24_and4162_y0;
  wire h_u_cla24_and4163_y0;
  wire h_u_cla24_and4164_y0;
  wire h_u_cla24_and4165_y0;
  wire h_u_cla24_and4166_y0;
  wire h_u_cla24_and4167_y0;
  wire h_u_cla24_and4168_y0;
  wire h_u_cla24_and4169_y0;
  wire h_u_cla24_and4170_y0;
  wire h_u_cla24_and4171_y0;
  wire h_u_cla24_and4172_y0;
  wire h_u_cla24_and4173_y0;
  wire h_u_cla24_and4174_y0;
  wire h_u_cla24_and4175_y0;
  wire h_u_cla24_and4176_y0;
  wire h_u_cla24_and4177_y0;
  wire h_u_cla24_and4178_y0;
  wire h_u_cla24_and4179_y0;
  wire h_u_cla24_and4180_y0;
  wire h_u_cla24_and4181_y0;
  wire h_u_cla24_and4182_y0;
  wire h_u_cla24_and4183_y0;
  wire h_u_cla24_and4184_y0;
  wire h_u_cla24_and4185_y0;
  wire h_u_cla24_and4186_y0;
  wire h_u_cla24_and4187_y0;
  wire h_u_cla24_and4188_y0;
  wire h_u_cla24_and4189_y0;
  wire h_u_cla24_and4190_y0;
  wire h_u_cla24_and4191_y0;
  wire h_u_cla24_and4192_y0;
  wire h_u_cla24_and4193_y0;
  wire h_u_cla24_and4194_y0;
  wire h_u_cla24_and4195_y0;
  wire h_u_cla24_and4196_y0;
  wire h_u_cla24_and4197_y0;
  wire h_u_cla24_and4198_y0;
  wire h_u_cla24_and4199_y0;
  wire h_u_cla24_and4200_y0;
  wire h_u_cla24_and4201_y0;
  wire h_u_cla24_and4202_y0;
  wire h_u_cla24_and4203_y0;
  wire h_u_cla24_and4204_y0;
  wire h_u_cla24_and4205_y0;
  wire h_u_cla24_and4206_y0;
  wire h_u_cla24_and4207_y0;
  wire h_u_cla24_and4208_y0;
  wire h_u_cla24_and4209_y0;
  wire h_u_cla24_and4210_y0;
  wire h_u_cla24_and4211_y0;
  wire h_u_cla24_and4212_y0;
  wire h_u_cla24_and4213_y0;
  wire h_u_cla24_and4214_y0;
  wire h_u_cla24_and4215_y0;
  wire h_u_cla24_and4216_y0;
  wire h_u_cla24_and4217_y0;
  wire h_u_cla24_and4218_y0;
  wire h_u_cla24_and4219_y0;
  wire h_u_cla24_and4220_y0;
  wire h_u_cla24_and4221_y0;
  wire h_u_cla24_and4222_y0;
  wire h_u_cla24_and4223_y0;
  wire h_u_cla24_and4224_y0;
  wire h_u_cla24_and4225_y0;
  wire h_u_cla24_and4226_y0;
  wire h_u_cla24_and4227_y0;
  wire h_u_cla24_and4228_y0;
  wire h_u_cla24_and4229_y0;
  wire h_u_cla24_and4230_y0;
  wire h_u_cla24_and4231_y0;
  wire h_u_cla24_and4232_y0;
  wire h_u_cla24_and4233_y0;
  wire h_u_cla24_and4234_y0;
  wire h_u_cla24_and4235_y0;
  wire h_u_cla24_and4236_y0;
  wire h_u_cla24_and4237_y0;
  wire h_u_cla24_and4238_y0;
  wire h_u_cla24_and4239_y0;
  wire h_u_cla24_and4240_y0;
  wire h_u_cla24_and4241_y0;
  wire h_u_cla24_and4242_y0;
  wire h_u_cla24_and4243_y0;
  wire h_u_cla24_and4244_y0;
  wire h_u_cla24_and4245_y0;
  wire h_u_cla24_and4246_y0;
  wire h_u_cla24_and4247_y0;
  wire h_u_cla24_and4248_y0;
  wire h_u_cla24_and4249_y0;
  wire h_u_cla24_and4250_y0;
  wire h_u_cla24_and4251_y0;
  wire h_u_cla24_and4252_y0;
  wire h_u_cla24_and4253_y0;
  wire h_u_cla24_and4254_y0;
  wire h_u_cla24_and4255_y0;
  wire h_u_cla24_and4256_y0;
  wire h_u_cla24_and4257_y0;
  wire h_u_cla24_and4258_y0;
  wire h_u_cla24_and4259_y0;
  wire h_u_cla24_and4260_y0;
  wire h_u_cla24_and4261_y0;
  wire h_u_cla24_and4262_y0;
  wire h_u_cla24_and4263_y0;
  wire h_u_cla24_and4264_y0;
  wire h_u_cla24_and4265_y0;
  wire h_u_cla24_and4266_y0;
  wire h_u_cla24_and4267_y0;
  wire h_u_cla24_and4268_y0;
  wire h_u_cla24_and4269_y0;
  wire h_u_cla24_and4270_y0;
  wire h_u_cla24_and4271_y0;
  wire h_u_cla24_and4272_y0;
  wire h_u_cla24_and4273_y0;
  wire h_u_cla24_and4274_y0;
  wire h_u_cla24_and4275_y0;
  wire h_u_cla24_and4276_y0;
  wire h_u_cla24_and4277_y0;
  wire h_u_cla24_and4278_y0;
  wire h_u_cla24_and4279_y0;
  wire h_u_cla24_and4280_y0;
  wire h_u_cla24_and4281_y0;
  wire h_u_cla24_and4282_y0;
  wire h_u_cla24_and4283_y0;
  wire h_u_cla24_and4284_y0;
  wire h_u_cla24_and4285_y0;
  wire h_u_cla24_and4286_y0;
  wire h_u_cla24_and4287_y0;
  wire h_u_cla24_and4288_y0;
  wire h_u_cla24_and4289_y0;
  wire h_u_cla24_and4290_y0;
  wire h_u_cla24_and4291_y0;
  wire h_u_cla24_and4292_y0;
  wire h_u_cla24_and4293_y0;
  wire h_u_cla24_and4294_y0;
  wire h_u_cla24_and4295_y0;
  wire h_u_cla24_and4296_y0;
  wire h_u_cla24_and4297_y0;
  wire h_u_cla24_and4298_y0;
  wire h_u_cla24_and4299_y0;
  wire h_u_cla24_and4300_y0;
  wire h_u_cla24_and4301_y0;
  wire h_u_cla24_and4302_y0;
  wire h_u_cla24_and4303_y0;
  wire h_u_cla24_and4304_y0;
  wire h_u_cla24_and4305_y0;
  wire h_u_cla24_and4306_y0;
  wire h_u_cla24_and4307_y0;
  wire h_u_cla24_and4308_y0;
  wire h_u_cla24_and4309_y0;
  wire h_u_cla24_and4310_y0;
  wire h_u_cla24_and4311_y0;
  wire h_u_cla24_and4312_y0;
  wire h_u_cla24_and4313_y0;
  wire h_u_cla24_and4314_y0;
  wire h_u_cla24_and4315_y0;
  wire h_u_cla24_and4316_y0;
  wire h_u_cla24_and4317_y0;
  wire h_u_cla24_and4318_y0;
  wire h_u_cla24_and4319_y0;
  wire h_u_cla24_and4320_y0;
  wire h_u_cla24_and4321_y0;
  wire h_u_cla24_and4322_y0;
  wire h_u_cla24_and4323_y0;
  wire h_u_cla24_or253_y0;
  wire h_u_cla24_or254_y0;
  wire h_u_cla24_or255_y0;
  wire h_u_cla24_or256_y0;
  wire h_u_cla24_or257_y0;
  wire h_u_cla24_or258_y0;
  wire h_u_cla24_or259_y0;
  wire h_u_cla24_or260_y0;
  wire h_u_cla24_or261_y0;
  wire h_u_cla24_or262_y0;
  wire h_u_cla24_or263_y0;
  wire h_u_cla24_or264_y0;
  wire h_u_cla24_or265_y0;
  wire h_u_cla24_or266_y0;
  wire h_u_cla24_or267_y0;
  wire h_u_cla24_or268_y0;
  wire h_u_cla24_or269_y0;
  wire h_u_cla24_or270_y0;
  wire h_u_cla24_or271_y0;
  wire h_u_cla24_or272_y0;
  wire h_u_cla24_or273_y0;
  wire h_u_cla24_or274_y0;
  wire h_u_cla24_or275_y0;
  wire h_u_cla24_pg_logic23_y0;
  wire h_u_cla24_pg_logic23_y1;
  wire h_u_cla24_pg_logic23_y2;
  wire h_u_cla24_xor23_y0;
  wire h_u_cla24_and4324_y0;
  wire h_u_cla24_and4325_y0;
  wire h_u_cla24_and4326_y0;
  wire h_u_cla24_and4327_y0;
  wire h_u_cla24_and4328_y0;
  wire h_u_cla24_and4329_y0;
  wire h_u_cla24_and4330_y0;
  wire h_u_cla24_and4331_y0;
  wire h_u_cla24_and4332_y0;
  wire h_u_cla24_and4333_y0;
  wire h_u_cla24_and4334_y0;
  wire h_u_cla24_and4335_y0;
  wire h_u_cla24_and4336_y0;
  wire h_u_cla24_and4337_y0;
  wire h_u_cla24_and4338_y0;
  wire h_u_cla24_and4339_y0;
  wire h_u_cla24_and4340_y0;
  wire h_u_cla24_and4341_y0;
  wire h_u_cla24_and4342_y0;
  wire h_u_cla24_and4343_y0;
  wire h_u_cla24_and4344_y0;
  wire h_u_cla24_and4345_y0;
  wire h_u_cla24_and4346_y0;
  wire h_u_cla24_and4347_y0;
  wire h_u_cla24_and4348_y0;
  wire h_u_cla24_and4349_y0;
  wire h_u_cla24_and4350_y0;
  wire h_u_cla24_and4351_y0;
  wire h_u_cla24_and4352_y0;
  wire h_u_cla24_and4353_y0;
  wire h_u_cla24_and4354_y0;
  wire h_u_cla24_and4355_y0;
  wire h_u_cla24_and4356_y0;
  wire h_u_cla24_and4357_y0;
  wire h_u_cla24_and4358_y0;
  wire h_u_cla24_and4359_y0;
  wire h_u_cla24_and4360_y0;
  wire h_u_cla24_and4361_y0;
  wire h_u_cla24_and4362_y0;
  wire h_u_cla24_and4363_y0;
  wire h_u_cla24_and4364_y0;
  wire h_u_cla24_and4365_y0;
  wire h_u_cla24_and4366_y0;
  wire h_u_cla24_and4367_y0;
  wire h_u_cla24_and4368_y0;
  wire h_u_cla24_and4369_y0;
  wire h_u_cla24_and4370_y0;
  wire h_u_cla24_and4371_y0;
  wire h_u_cla24_and4372_y0;
  wire h_u_cla24_and4373_y0;
  wire h_u_cla24_and4374_y0;
  wire h_u_cla24_and4375_y0;
  wire h_u_cla24_and4376_y0;
  wire h_u_cla24_and4377_y0;
  wire h_u_cla24_and4378_y0;
  wire h_u_cla24_and4379_y0;
  wire h_u_cla24_and4380_y0;
  wire h_u_cla24_and4381_y0;
  wire h_u_cla24_and4382_y0;
  wire h_u_cla24_and4383_y0;
  wire h_u_cla24_and4384_y0;
  wire h_u_cla24_and4385_y0;
  wire h_u_cla24_and4386_y0;
  wire h_u_cla24_and4387_y0;
  wire h_u_cla24_and4388_y0;
  wire h_u_cla24_and4389_y0;
  wire h_u_cla24_and4390_y0;
  wire h_u_cla24_and4391_y0;
  wire h_u_cla24_and4392_y0;
  wire h_u_cla24_and4393_y0;
  wire h_u_cla24_and4394_y0;
  wire h_u_cla24_and4395_y0;
  wire h_u_cla24_and4396_y0;
  wire h_u_cla24_and4397_y0;
  wire h_u_cla24_and4398_y0;
  wire h_u_cla24_and4399_y0;
  wire h_u_cla24_and4400_y0;
  wire h_u_cla24_and4401_y0;
  wire h_u_cla24_and4402_y0;
  wire h_u_cla24_and4403_y0;
  wire h_u_cla24_and4404_y0;
  wire h_u_cla24_and4405_y0;
  wire h_u_cla24_and4406_y0;
  wire h_u_cla24_and4407_y0;
  wire h_u_cla24_and4408_y0;
  wire h_u_cla24_and4409_y0;
  wire h_u_cla24_and4410_y0;
  wire h_u_cla24_and4411_y0;
  wire h_u_cla24_and4412_y0;
  wire h_u_cla24_and4413_y0;
  wire h_u_cla24_and4414_y0;
  wire h_u_cla24_and4415_y0;
  wire h_u_cla24_and4416_y0;
  wire h_u_cla24_and4417_y0;
  wire h_u_cla24_and4418_y0;
  wire h_u_cla24_and4419_y0;
  wire h_u_cla24_and4420_y0;
  wire h_u_cla24_and4421_y0;
  wire h_u_cla24_and4422_y0;
  wire h_u_cla24_and4423_y0;
  wire h_u_cla24_and4424_y0;
  wire h_u_cla24_and4425_y0;
  wire h_u_cla24_and4426_y0;
  wire h_u_cla24_and4427_y0;
  wire h_u_cla24_and4428_y0;
  wire h_u_cla24_and4429_y0;
  wire h_u_cla24_and4430_y0;
  wire h_u_cla24_and4431_y0;
  wire h_u_cla24_and4432_y0;
  wire h_u_cla24_and4433_y0;
  wire h_u_cla24_and4434_y0;
  wire h_u_cla24_and4435_y0;
  wire h_u_cla24_and4436_y0;
  wire h_u_cla24_and4437_y0;
  wire h_u_cla24_and4438_y0;
  wire h_u_cla24_and4439_y0;
  wire h_u_cla24_and4440_y0;
  wire h_u_cla24_and4441_y0;
  wire h_u_cla24_and4442_y0;
  wire h_u_cla24_and4443_y0;
  wire h_u_cla24_and4444_y0;
  wire h_u_cla24_and4445_y0;
  wire h_u_cla24_and4446_y0;
  wire h_u_cla24_and4447_y0;
  wire h_u_cla24_and4448_y0;
  wire h_u_cla24_and4449_y0;
  wire h_u_cla24_and4450_y0;
  wire h_u_cla24_and4451_y0;
  wire h_u_cla24_and4452_y0;
  wire h_u_cla24_and4453_y0;
  wire h_u_cla24_and4454_y0;
  wire h_u_cla24_and4455_y0;
  wire h_u_cla24_and4456_y0;
  wire h_u_cla24_and4457_y0;
  wire h_u_cla24_and4458_y0;
  wire h_u_cla24_and4459_y0;
  wire h_u_cla24_and4460_y0;
  wire h_u_cla24_and4461_y0;
  wire h_u_cla24_and4462_y0;
  wire h_u_cla24_and4463_y0;
  wire h_u_cla24_and4464_y0;
  wire h_u_cla24_and4465_y0;
  wire h_u_cla24_and4466_y0;
  wire h_u_cla24_and4467_y0;
  wire h_u_cla24_and4468_y0;
  wire h_u_cla24_and4469_y0;
  wire h_u_cla24_and4470_y0;
  wire h_u_cla24_and4471_y0;
  wire h_u_cla24_and4472_y0;
  wire h_u_cla24_and4473_y0;
  wire h_u_cla24_and4474_y0;
  wire h_u_cla24_and4475_y0;
  wire h_u_cla24_and4476_y0;
  wire h_u_cla24_and4477_y0;
  wire h_u_cla24_and4478_y0;
  wire h_u_cla24_and4479_y0;
  wire h_u_cla24_and4480_y0;
  wire h_u_cla24_and4481_y0;
  wire h_u_cla24_and4482_y0;
  wire h_u_cla24_and4483_y0;
  wire h_u_cla24_and4484_y0;
  wire h_u_cla24_and4485_y0;
  wire h_u_cla24_and4486_y0;
  wire h_u_cla24_and4487_y0;
  wire h_u_cla24_and4488_y0;
  wire h_u_cla24_and4489_y0;
  wire h_u_cla24_and4490_y0;
  wire h_u_cla24_and4491_y0;
  wire h_u_cla24_and4492_y0;
  wire h_u_cla24_and4493_y0;
  wire h_u_cla24_and4494_y0;
  wire h_u_cla24_and4495_y0;
  wire h_u_cla24_and4496_y0;
  wire h_u_cla24_and4497_y0;
  wire h_u_cla24_and4498_y0;
  wire h_u_cla24_and4499_y0;
  wire h_u_cla24_and4500_y0;
  wire h_u_cla24_and4501_y0;
  wire h_u_cla24_and4502_y0;
  wire h_u_cla24_and4503_y0;
  wire h_u_cla24_and4504_y0;
  wire h_u_cla24_and4505_y0;
  wire h_u_cla24_and4506_y0;
  wire h_u_cla24_and4507_y0;
  wire h_u_cla24_and4508_y0;
  wire h_u_cla24_and4509_y0;
  wire h_u_cla24_and4510_y0;
  wire h_u_cla24_and4511_y0;
  wire h_u_cla24_and4512_y0;
  wire h_u_cla24_and4513_y0;
  wire h_u_cla24_and4514_y0;
  wire h_u_cla24_and4515_y0;
  wire h_u_cla24_and4516_y0;
  wire h_u_cla24_and4517_y0;
  wire h_u_cla24_and4518_y0;
  wire h_u_cla24_and4519_y0;
  wire h_u_cla24_and4520_y0;
  wire h_u_cla24_and4521_y0;
  wire h_u_cla24_and4522_y0;
  wire h_u_cla24_and4523_y0;
  wire h_u_cla24_and4524_y0;
  wire h_u_cla24_and4525_y0;
  wire h_u_cla24_and4526_y0;
  wire h_u_cla24_and4527_y0;
  wire h_u_cla24_and4528_y0;
  wire h_u_cla24_and4529_y0;
  wire h_u_cla24_and4530_y0;
  wire h_u_cla24_and4531_y0;
  wire h_u_cla24_and4532_y0;
  wire h_u_cla24_and4533_y0;
  wire h_u_cla24_and4534_y0;
  wire h_u_cla24_and4535_y0;
  wire h_u_cla24_and4536_y0;
  wire h_u_cla24_and4537_y0;
  wire h_u_cla24_and4538_y0;
  wire h_u_cla24_and4539_y0;
  wire h_u_cla24_and4540_y0;
  wire h_u_cla24_and4541_y0;
  wire h_u_cla24_and4542_y0;
  wire h_u_cla24_and4543_y0;
  wire h_u_cla24_and4544_y0;
  wire h_u_cla24_and4545_y0;
  wire h_u_cla24_and4546_y0;
  wire h_u_cla24_and4547_y0;
  wire h_u_cla24_and4548_y0;
  wire h_u_cla24_and4549_y0;
  wire h_u_cla24_and4550_y0;
  wire h_u_cla24_and4551_y0;
  wire h_u_cla24_and4552_y0;
  wire h_u_cla24_and4553_y0;
  wire h_u_cla24_and4554_y0;
  wire h_u_cla24_and4555_y0;
  wire h_u_cla24_and4556_y0;
  wire h_u_cla24_and4557_y0;
  wire h_u_cla24_and4558_y0;
  wire h_u_cla24_and4559_y0;
  wire h_u_cla24_and4560_y0;
  wire h_u_cla24_and4561_y0;
  wire h_u_cla24_and4562_y0;
  wire h_u_cla24_and4563_y0;
  wire h_u_cla24_and4564_y0;
  wire h_u_cla24_and4565_y0;
  wire h_u_cla24_and4566_y0;
  wire h_u_cla24_and4567_y0;
  wire h_u_cla24_and4568_y0;
  wire h_u_cla24_and4569_y0;
  wire h_u_cla24_and4570_y0;
  wire h_u_cla24_and4571_y0;
  wire h_u_cla24_and4572_y0;
  wire h_u_cla24_and4573_y0;
  wire h_u_cla24_and4574_y0;
  wire h_u_cla24_and4575_y0;
  wire h_u_cla24_and4576_y0;
  wire h_u_cla24_and4577_y0;
  wire h_u_cla24_and4578_y0;
  wire h_u_cla24_and4579_y0;
  wire h_u_cla24_and4580_y0;
  wire h_u_cla24_and4581_y0;
  wire h_u_cla24_and4582_y0;
  wire h_u_cla24_and4583_y0;
  wire h_u_cla24_and4584_y0;
  wire h_u_cla24_and4585_y0;
  wire h_u_cla24_and4586_y0;
  wire h_u_cla24_and4587_y0;
  wire h_u_cla24_and4588_y0;
  wire h_u_cla24_and4589_y0;
  wire h_u_cla24_and4590_y0;
  wire h_u_cla24_and4591_y0;
  wire h_u_cla24_and4592_y0;
  wire h_u_cla24_and4593_y0;
  wire h_u_cla24_and4594_y0;
  wire h_u_cla24_and4595_y0;
  wire h_u_cla24_and4596_y0;
  wire h_u_cla24_and4597_y0;
  wire h_u_cla24_and4598_y0;
  wire h_u_cla24_and4599_y0;
  wire h_u_cla24_and4600_y0;
  wire h_u_cla24_and4601_y0;
  wire h_u_cla24_and4602_y0;
  wire h_u_cla24_and4603_y0;
  wire h_u_cla24_and4604_y0;
  wire h_u_cla24_and4605_y0;
  wire h_u_cla24_and4606_y0;
  wire h_u_cla24_and4607_y0;
  wire h_u_cla24_and4608_y0;
  wire h_u_cla24_and4609_y0;
  wire h_u_cla24_and4610_y0;
  wire h_u_cla24_and4611_y0;
  wire h_u_cla24_and4612_y0;
  wire h_u_cla24_and4613_y0;
  wire h_u_cla24_and4614_y0;
  wire h_u_cla24_and4615_y0;
  wire h_u_cla24_and4616_y0;
  wire h_u_cla24_and4617_y0;
  wire h_u_cla24_and4618_y0;
  wire h_u_cla24_and4619_y0;
  wire h_u_cla24_and4620_y0;
  wire h_u_cla24_and4621_y0;
  wire h_u_cla24_and4622_y0;
  wire h_u_cla24_and4623_y0;
  wire h_u_cla24_and4624_y0;
  wire h_u_cla24_and4625_y0;
  wire h_u_cla24_and4626_y0;
  wire h_u_cla24_and4627_y0;
  wire h_u_cla24_and4628_y0;
  wire h_u_cla24_and4629_y0;
  wire h_u_cla24_and4630_y0;
  wire h_u_cla24_and4631_y0;
  wire h_u_cla24_and4632_y0;
  wire h_u_cla24_and4633_y0;
  wire h_u_cla24_and4634_y0;
  wire h_u_cla24_and4635_y0;
  wire h_u_cla24_and4636_y0;
  wire h_u_cla24_and4637_y0;
  wire h_u_cla24_and4638_y0;
  wire h_u_cla24_and4639_y0;
  wire h_u_cla24_and4640_y0;
  wire h_u_cla24_and4641_y0;
  wire h_u_cla24_and4642_y0;
  wire h_u_cla24_and4643_y0;
  wire h_u_cla24_and4644_y0;
  wire h_u_cla24_and4645_y0;
  wire h_u_cla24_and4646_y0;
  wire h_u_cla24_and4647_y0;
  wire h_u_cla24_and4648_y0;
  wire h_u_cla24_and4649_y0;
  wire h_u_cla24_and4650_y0;
  wire h_u_cla24_and4651_y0;
  wire h_u_cla24_and4652_y0;
  wire h_u_cla24_and4653_y0;
  wire h_u_cla24_and4654_y0;
  wire h_u_cla24_and4655_y0;
  wire h_u_cla24_and4656_y0;
  wire h_u_cla24_and4657_y0;
  wire h_u_cla24_and4658_y0;
  wire h_u_cla24_and4659_y0;
  wire h_u_cla24_and4660_y0;
  wire h_u_cla24_and4661_y0;
  wire h_u_cla24_and4662_y0;
  wire h_u_cla24_and4663_y0;
  wire h_u_cla24_and4664_y0;
  wire h_u_cla24_and4665_y0;
  wire h_u_cla24_and4666_y0;
  wire h_u_cla24_and4667_y0;
  wire h_u_cla24_and4668_y0;
  wire h_u_cla24_and4669_y0;
  wire h_u_cla24_and4670_y0;
  wire h_u_cla24_and4671_y0;
  wire h_u_cla24_and4672_y0;
  wire h_u_cla24_and4673_y0;
  wire h_u_cla24_and4674_y0;
  wire h_u_cla24_and4675_y0;
  wire h_u_cla24_and4676_y0;
  wire h_u_cla24_and4677_y0;
  wire h_u_cla24_and4678_y0;
  wire h_u_cla24_and4679_y0;
  wire h_u_cla24_and4680_y0;
  wire h_u_cla24_and4681_y0;
  wire h_u_cla24_and4682_y0;
  wire h_u_cla24_and4683_y0;
  wire h_u_cla24_and4684_y0;
  wire h_u_cla24_and4685_y0;
  wire h_u_cla24_and4686_y0;
  wire h_u_cla24_and4687_y0;
  wire h_u_cla24_and4688_y0;
  wire h_u_cla24_and4689_y0;
  wire h_u_cla24_and4690_y0;
  wire h_u_cla24_and4691_y0;
  wire h_u_cla24_and4692_y0;
  wire h_u_cla24_and4693_y0;
  wire h_u_cla24_and4694_y0;
  wire h_u_cla24_and4695_y0;
  wire h_u_cla24_and4696_y0;
  wire h_u_cla24_and4697_y0;
  wire h_u_cla24_and4698_y0;
  wire h_u_cla24_and4699_y0;
  wire h_u_cla24_and4700_y0;
  wire h_u_cla24_and4701_y0;
  wire h_u_cla24_and4702_y0;
  wire h_u_cla24_and4703_y0;
  wire h_u_cla24_and4704_y0;
  wire h_u_cla24_and4705_y0;
  wire h_u_cla24_and4706_y0;
  wire h_u_cla24_and4707_y0;
  wire h_u_cla24_and4708_y0;
  wire h_u_cla24_and4709_y0;
  wire h_u_cla24_and4710_y0;
  wire h_u_cla24_and4711_y0;
  wire h_u_cla24_and4712_y0;
  wire h_u_cla24_and4713_y0;
  wire h_u_cla24_and4714_y0;
  wire h_u_cla24_and4715_y0;
  wire h_u_cla24_and4716_y0;
  wire h_u_cla24_and4717_y0;
  wire h_u_cla24_and4718_y0;
  wire h_u_cla24_and4719_y0;
  wire h_u_cla24_and4720_y0;
  wire h_u_cla24_and4721_y0;
  wire h_u_cla24_and4722_y0;
  wire h_u_cla24_and4723_y0;
  wire h_u_cla24_and4724_y0;
  wire h_u_cla24_and4725_y0;
  wire h_u_cla24_and4726_y0;
  wire h_u_cla24_and4727_y0;
  wire h_u_cla24_and4728_y0;
  wire h_u_cla24_and4729_y0;
  wire h_u_cla24_and4730_y0;
  wire h_u_cla24_and4731_y0;
  wire h_u_cla24_and4732_y0;
  wire h_u_cla24_and4733_y0;
  wire h_u_cla24_and4734_y0;
  wire h_u_cla24_and4735_y0;
  wire h_u_cla24_and4736_y0;
  wire h_u_cla24_and4737_y0;
  wire h_u_cla24_and4738_y0;
  wire h_u_cla24_and4739_y0;
  wire h_u_cla24_and4740_y0;
  wire h_u_cla24_and4741_y0;
  wire h_u_cla24_and4742_y0;
  wire h_u_cla24_and4743_y0;
  wire h_u_cla24_and4744_y0;
  wire h_u_cla24_and4745_y0;
  wire h_u_cla24_and4746_y0;
  wire h_u_cla24_and4747_y0;
  wire h_u_cla24_and4748_y0;
  wire h_u_cla24_and4749_y0;
  wire h_u_cla24_and4750_y0;
  wire h_u_cla24_and4751_y0;
  wire h_u_cla24_and4752_y0;
  wire h_u_cla24_and4753_y0;
  wire h_u_cla24_and4754_y0;
  wire h_u_cla24_and4755_y0;
  wire h_u_cla24_and4756_y0;
  wire h_u_cla24_and4757_y0;
  wire h_u_cla24_and4758_y0;
  wire h_u_cla24_and4759_y0;
  wire h_u_cla24_and4760_y0;
  wire h_u_cla24_and4761_y0;
  wire h_u_cla24_and4762_y0;
  wire h_u_cla24_and4763_y0;
  wire h_u_cla24_and4764_y0;
  wire h_u_cla24_and4765_y0;
  wire h_u_cla24_and4766_y0;
  wire h_u_cla24_and4767_y0;
  wire h_u_cla24_and4768_y0;
  wire h_u_cla24_and4769_y0;
  wire h_u_cla24_and4770_y0;
  wire h_u_cla24_and4771_y0;
  wire h_u_cla24_and4772_y0;
  wire h_u_cla24_and4773_y0;
  wire h_u_cla24_and4774_y0;
  wire h_u_cla24_and4775_y0;
  wire h_u_cla24_and4776_y0;
  wire h_u_cla24_and4777_y0;
  wire h_u_cla24_and4778_y0;
  wire h_u_cla24_and4779_y0;
  wire h_u_cla24_and4780_y0;
  wire h_u_cla24_and4781_y0;
  wire h_u_cla24_and4782_y0;
  wire h_u_cla24_and4783_y0;
  wire h_u_cla24_and4784_y0;
  wire h_u_cla24_and4785_y0;
  wire h_u_cla24_and4786_y0;
  wire h_u_cla24_and4787_y0;
  wire h_u_cla24_and4788_y0;
  wire h_u_cla24_and4789_y0;
  wire h_u_cla24_and4790_y0;
  wire h_u_cla24_and4791_y0;
  wire h_u_cla24_and4792_y0;
  wire h_u_cla24_and4793_y0;
  wire h_u_cla24_and4794_y0;
  wire h_u_cla24_and4795_y0;
  wire h_u_cla24_and4796_y0;
  wire h_u_cla24_and4797_y0;
  wire h_u_cla24_and4798_y0;
  wire h_u_cla24_and4799_y0;
  wire h_u_cla24_and4800_y0;
  wire h_u_cla24_and4801_y0;
  wire h_u_cla24_and4802_y0;
  wire h_u_cla24_and4803_y0;
  wire h_u_cla24_and4804_y0;
  wire h_u_cla24_and4805_y0;
  wire h_u_cla24_and4806_y0;
  wire h_u_cla24_and4807_y0;
  wire h_u_cla24_and4808_y0;
  wire h_u_cla24_and4809_y0;
  wire h_u_cla24_and4810_y0;
  wire h_u_cla24_and4811_y0;
  wire h_u_cla24_and4812_y0;
  wire h_u_cla24_and4813_y0;
  wire h_u_cla24_and4814_y0;
  wire h_u_cla24_and4815_y0;
  wire h_u_cla24_and4816_y0;
  wire h_u_cla24_and4817_y0;
  wire h_u_cla24_and4818_y0;
  wire h_u_cla24_and4819_y0;
  wire h_u_cla24_and4820_y0;
  wire h_u_cla24_and4821_y0;
  wire h_u_cla24_and4822_y0;
  wire h_u_cla24_and4823_y0;
  wire h_u_cla24_and4824_y0;
  wire h_u_cla24_and4825_y0;
  wire h_u_cla24_and4826_y0;
  wire h_u_cla24_and4827_y0;
  wire h_u_cla24_and4828_y0;
  wire h_u_cla24_and4829_y0;
  wire h_u_cla24_and4830_y0;
  wire h_u_cla24_and4831_y0;
  wire h_u_cla24_and4832_y0;
  wire h_u_cla24_and4833_y0;
  wire h_u_cla24_and4834_y0;
  wire h_u_cla24_and4835_y0;
  wire h_u_cla24_and4836_y0;
  wire h_u_cla24_and4837_y0;
  wire h_u_cla24_and4838_y0;
  wire h_u_cla24_and4839_y0;
  wire h_u_cla24_and4840_y0;
  wire h_u_cla24_and4841_y0;
  wire h_u_cla24_and4842_y0;
  wire h_u_cla24_and4843_y0;
  wire h_u_cla24_and4844_y0;
  wire h_u_cla24_and4845_y0;
  wire h_u_cla24_and4846_y0;
  wire h_u_cla24_and4847_y0;
  wire h_u_cla24_and4848_y0;
  wire h_u_cla24_and4849_y0;
  wire h_u_cla24_and4850_y0;
  wire h_u_cla24_and4851_y0;
  wire h_u_cla24_and4852_y0;
  wire h_u_cla24_and4853_y0;
  wire h_u_cla24_and4854_y0;
  wire h_u_cla24_and4855_y0;
  wire h_u_cla24_and4856_y0;
  wire h_u_cla24_and4857_y0;
  wire h_u_cla24_and4858_y0;
  wire h_u_cla24_and4859_y0;
  wire h_u_cla24_and4860_y0;
  wire h_u_cla24_and4861_y0;
  wire h_u_cla24_and4862_y0;
  wire h_u_cla24_and4863_y0;
  wire h_u_cla24_and4864_y0;
  wire h_u_cla24_and4865_y0;
  wire h_u_cla24_and4866_y0;
  wire h_u_cla24_and4867_y0;
  wire h_u_cla24_and4868_y0;
  wire h_u_cla24_and4869_y0;
  wire h_u_cla24_and4870_y0;
  wire h_u_cla24_and4871_y0;
  wire h_u_cla24_and4872_y0;
  wire h_u_cla24_and4873_y0;
  wire h_u_cla24_and4874_y0;
  wire h_u_cla24_and4875_y0;
  wire h_u_cla24_and4876_y0;
  wire h_u_cla24_and4877_y0;
  wire h_u_cla24_and4878_y0;
  wire h_u_cla24_and4879_y0;
  wire h_u_cla24_and4880_y0;
  wire h_u_cla24_and4881_y0;
  wire h_u_cla24_and4882_y0;
  wire h_u_cla24_and4883_y0;
  wire h_u_cla24_and4884_y0;
  wire h_u_cla24_and4885_y0;
  wire h_u_cla24_and4886_y0;
  wire h_u_cla24_and4887_y0;
  wire h_u_cla24_and4888_y0;
  wire h_u_cla24_and4889_y0;
  wire h_u_cla24_and4890_y0;
  wire h_u_cla24_and4891_y0;
  wire h_u_cla24_and4892_y0;
  wire h_u_cla24_and4893_y0;
  wire h_u_cla24_and4894_y0;
  wire h_u_cla24_and4895_y0;
  wire h_u_cla24_and4896_y0;
  wire h_u_cla24_and4897_y0;
  wire h_u_cla24_and4898_y0;
  wire h_u_cla24_and4899_y0;
  wire h_u_cla24_or276_y0;
  wire h_u_cla24_or277_y0;
  wire h_u_cla24_or278_y0;
  wire h_u_cla24_or279_y0;
  wire h_u_cla24_or280_y0;
  wire h_u_cla24_or281_y0;
  wire h_u_cla24_or282_y0;
  wire h_u_cla24_or283_y0;
  wire h_u_cla24_or284_y0;
  wire h_u_cla24_or285_y0;
  wire h_u_cla24_or286_y0;
  wire h_u_cla24_or287_y0;
  wire h_u_cla24_or288_y0;
  wire h_u_cla24_or289_y0;
  wire h_u_cla24_or290_y0;
  wire h_u_cla24_or291_y0;
  wire h_u_cla24_or292_y0;
  wire h_u_cla24_or293_y0;
  wire h_u_cla24_or294_y0;
  wire h_u_cla24_or295_y0;
  wire h_u_cla24_or296_y0;
  wire h_u_cla24_or297_y0;
  wire h_u_cla24_or298_y0;
  wire h_u_cla24_or299_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  constant_wire_value_0 constant_wire_value_0_constant_wire_0(a_0, b_0, constant_wire_0);
  pg_logic pg_logic_h_u_cla24_pg_logic0_y0(a_0, b_0, h_u_cla24_pg_logic0_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_pg_logic0_y2);
  xor_gate xor_gate_h_u_cla24_xor0_y0(h_u_cla24_pg_logic0_y2, constant_wire_0, h_u_cla24_xor0_y0);
  and_gate and_gate_h_u_cla24_and0_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and0_y0);
  or_gate or_gate_h_u_cla24_or0_y0(h_u_cla24_pg_logic0_y1, h_u_cla24_and0_y0, h_u_cla24_or0_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic1_y0(a_1, b_1, h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_pg_logic1_y2);
  xor_gate xor_gate_h_u_cla24_xor1_y0(h_u_cla24_pg_logic1_y2, h_u_cla24_or0_y0, h_u_cla24_xor1_y0);
  and_gate and_gate_h_u_cla24_and1_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and1_y0);
  and_gate and_gate_h_u_cla24_and2_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and2_y0);
  and_gate and_gate_h_u_cla24_and3_y0(h_u_cla24_and2_y0, h_u_cla24_and1_y0, h_u_cla24_and3_y0);
  and_gate and_gate_h_u_cla24_and4_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4_y0);
  or_gate or_gate_h_u_cla24_or1_y0(h_u_cla24_and4_y0, h_u_cla24_and3_y0, h_u_cla24_or1_y0);
  or_gate or_gate_h_u_cla24_or2_y0(h_u_cla24_pg_logic1_y1, h_u_cla24_or1_y0, h_u_cla24_or2_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic2_y0(a_2, b_2, h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_pg_logic2_y2);
  xor_gate xor_gate_h_u_cla24_xor2_y0(h_u_cla24_pg_logic2_y2, h_u_cla24_or2_y0, h_u_cla24_xor2_y0);
  and_gate and_gate_h_u_cla24_and5_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and5_y0);
  and_gate and_gate_h_u_cla24_and6_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and6_y0);
  and_gate and_gate_h_u_cla24_and7_y0(h_u_cla24_and6_y0, h_u_cla24_and5_y0, h_u_cla24_and7_y0);
  and_gate and_gate_h_u_cla24_and8_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and8_y0);
  and_gate and_gate_h_u_cla24_and9_y0(h_u_cla24_and8_y0, h_u_cla24_and7_y0, h_u_cla24_and9_y0);
  and_gate and_gate_h_u_cla24_and10_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and10_y0);
  and_gate and_gate_h_u_cla24_and11_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and11_y0);
  and_gate and_gate_h_u_cla24_and12_y0(h_u_cla24_and11_y0, h_u_cla24_and10_y0, h_u_cla24_and12_y0);
  and_gate and_gate_h_u_cla24_and13_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and13_y0);
  or_gate or_gate_h_u_cla24_or3_y0(h_u_cla24_and13_y0, h_u_cla24_and9_y0, h_u_cla24_or3_y0);
  or_gate or_gate_h_u_cla24_or4_y0(h_u_cla24_or3_y0, h_u_cla24_and12_y0, h_u_cla24_or4_y0);
  or_gate or_gate_h_u_cla24_or5_y0(h_u_cla24_pg_logic2_y1, h_u_cla24_or4_y0, h_u_cla24_or5_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic3_y0(a_3, b_3, h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_pg_logic3_y2);
  xor_gate xor_gate_h_u_cla24_xor3_y0(h_u_cla24_pg_logic3_y2, h_u_cla24_or5_y0, h_u_cla24_xor3_y0);
  and_gate and_gate_h_u_cla24_and14_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and14_y0);
  and_gate and_gate_h_u_cla24_and15_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and15_y0);
  and_gate and_gate_h_u_cla24_and16_y0(h_u_cla24_and15_y0, h_u_cla24_and14_y0, h_u_cla24_and16_y0);
  and_gate and_gate_h_u_cla24_and17_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and17_y0);
  and_gate and_gate_h_u_cla24_and18_y0(h_u_cla24_and17_y0, h_u_cla24_and16_y0, h_u_cla24_and18_y0);
  and_gate and_gate_h_u_cla24_and19_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and19_y0);
  and_gate and_gate_h_u_cla24_and20_y0(h_u_cla24_and19_y0, h_u_cla24_and18_y0, h_u_cla24_and20_y0);
  and_gate and_gate_h_u_cla24_and21_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and21_y0);
  and_gate and_gate_h_u_cla24_and22_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and22_y0);
  and_gate and_gate_h_u_cla24_and23_y0(h_u_cla24_and22_y0, h_u_cla24_and21_y0, h_u_cla24_and23_y0);
  and_gate and_gate_h_u_cla24_and24_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and24_y0);
  and_gate and_gate_h_u_cla24_and25_y0(h_u_cla24_and24_y0, h_u_cla24_and23_y0, h_u_cla24_and25_y0);
  and_gate and_gate_h_u_cla24_and26_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and26_y0);
  and_gate and_gate_h_u_cla24_and27_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and27_y0);
  and_gate and_gate_h_u_cla24_and28_y0(h_u_cla24_and27_y0, h_u_cla24_and26_y0, h_u_cla24_and28_y0);
  and_gate and_gate_h_u_cla24_and29_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and29_y0);
  or_gate or_gate_h_u_cla24_or6_y0(h_u_cla24_and29_y0, h_u_cla24_and20_y0, h_u_cla24_or6_y0);
  or_gate or_gate_h_u_cla24_or7_y0(h_u_cla24_or6_y0, h_u_cla24_and25_y0, h_u_cla24_or7_y0);
  or_gate or_gate_h_u_cla24_or8_y0(h_u_cla24_or7_y0, h_u_cla24_and28_y0, h_u_cla24_or8_y0);
  or_gate or_gate_h_u_cla24_or9_y0(h_u_cla24_pg_logic3_y1, h_u_cla24_or8_y0, h_u_cla24_or9_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic4_y0(a_4, b_4, h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_pg_logic4_y2);
  xor_gate xor_gate_h_u_cla24_xor4_y0(h_u_cla24_pg_logic4_y2, h_u_cla24_or9_y0, h_u_cla24_xor4_y0);
  and_gate and_gate_h_u_cla24_and30_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and30_y0);
  and_gate and_gate_h_u_cla24_and31_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and31_y0);
  and_gate and_gate_h_u_cla24_and32_y0(h_u_cla24_and31_y0, h_u_cla24_and30_y0, h_u_cla24_and32_y0);
  and_gate and_gate_h_u_cla24_and33_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and33_y0);
  and_gate and_gate_h_u_cla24_and34_y0(h_u_cla24_and33_y0, h_u_cla24_and32_y0, h_u_cla24_and34_y0);
  and_gate and_gate_h_u_cla24_and35_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and35_y0);
  and_gate and_gate_h_u_cla24_and36_y0(h_u_cla24_and35_y0, h_u_cla24_and34_y0, h_u_cla24_and36_y0);
  and_gate and_gate_h_u_cla24_and37_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and37_y0);
  and_gate and_gate_h_u_cla24_and38_y0(h_u_cla24_and37_y0, h_u_cla24_and36_y0, h_u_cla24_and38_y0);
  and_gate and_gate_h_u_cla24_and39_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and39_y0);
  and_gate and_gate_h_u_cla24_and40_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and40_y0);
  and_gate and_gate_h_u_cla24_and41_y0(h_u_cla24_and40_y0, h_u_cla24_and39_y0, h_u_cla24_and41_y0);
  and_gate and_gate_h_u_cla24_and42_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and42_y0);
  and_gate and_gate_h_u_cla24_and43_y0(h_u_cla24_and42_y0, h_u_cla24_and41_y0, h_u_cla24_and43_y0);
  and_gate and_gate_h_u_cla24_and44_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and44_y0);
  and_gate and_gate_h_u_cla24_and45_y0(h_u_cla24_and44_y0, h_u_cla24_and43_y0, h_u_cla24_and45_y0);
  and_gate and_gate_h_u_cla24_and46_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and46_y0);
  and_gate and_gate_h_u_cla24_and47_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and47_y0);
  and_gate and_gate_h_u_cla24_and48_y0(h_u_cla24_and47_y0, h_u_cla24_and46_y0, h_u_cla24_and48_y0);
  and_gate and_gate_h_u_cla24_and49_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and49_y0);
  and_gate and_gate_h_u_cla24_and50_y0(h_u_cla24_and49_y0, h_u_cla24_and48_y0, h_u_cla24_and50_y0);
  and_gate and_gate_h_u_cla24_and51_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and51_y0);
  and_gate and_gate_h_u_cla24_and52_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and52_y0);
  and_gate and_gate_h_u_cla24_and53_y0(h_u_cla24_and52_y0, h_u_cla24_and51_y0, h_u_cla24_and53_y0);
  and_gate and_gate_h_u_cla24_and54_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and54_y0);
  or_gate or_gate_h_u_cla24_or10_y0(h_u_cla24_and54_y0, h_u_cla24_and38_y0, h_u_cla24_or10_y0);
  or_gate or_gate_h_u_cla24_or11_y0(h_u_cla24_or10_y0, h_u_cla24_and45_y0, h_u_cla24_or11_y0);
  or_gate or_gate_h_u_cla24_or12_y0(h_u_cla24_or11_y0, h_u_cla24_and50_y0, h_u_cla24_or12_y0);
  or_gate or_gate_h_u_cla24_or13_y0(h_u_cla24_or12_y0, h_u_cla24_and53_y0, h_u_cla24_or13_y0);
  or_gate or_gate_h_u_cla24_or14_y0(h_u_cla24_pg_logic4_y1, h_u_cla24_or13_y0, h_u_cla24_or14_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic5_y0(a_5, b_5, h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_pg_logic5_y2);
  xor_gate xor_gate_h_u_cla24_xor5_y0(h_u_cla24_pg_logic5_y2, h_u_cla24_or14_y0, h_u_cla24_xor5_y0);
  and_gate and_gate_h_u_cla24_and55_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and55_y0);
  and_gate and_gate_h_u_cla24_and56_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and56_y0);
  and_gate and_gate_h_u_cla24_and57_y0(h_u_cla24_and56_y0, h_u_cla24_and55_y0, h_u_cla24_and57_y0);
  and_gate and_gate_h_u_cla24_and58_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and58_y0);
  and_gate and_gate_h_u_cla24_and59_y0(h_u_cla24_and58_y0, h_u_cla24_and57_y0, h_u_cla24_and59_y0);
  and_gate and_gate_h_u_cla24_and60_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and60_y0);
  and_gate and_gate_h_u_cla24_and61_y0(h_u_cla24_and60_y0, h_u_cla24_and59_y0, h_u_cla24_and61_y0);
  and_gate and_gate_h_u_cla24_and62_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and62_y0);
  and_gate and_gate_h_u_cla24_and63_y0(h_u_cla24_and62_y0, h_u_cla24_and61_y0, h_u_cla24_and63_y0);
  and_gate and_gate_h_u_cla24_and64_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and64_y0);
  and_gate and_gate_h_u_cla24_and65_y0(h_u_cla24_and64_y0, h_u_cla24_and63_y0, h_u_cla24_and65_y0);
  and_gate and_gate_h_u_cla24_and66_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and66_y0);
  and_gate and_gate_h_u_cla24_and67_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and67_y0);
  and_gate and_gate_h_u_cla24_and68_y0(h_u_cla24_and67_y0, h_u_cla24_and66_y0, h_u_cla24_and68_y0);
  and_gate and_gate_h_u_cla24_and69_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and69_y0);
  and_gate and_gate_h_u_cla24_and70_y0(h_u_cla24_and69_y0, h_u_cla24_and68_y0, h_u_cla24_and70_y0);
  and_gate and_gate_h_u_cla24_and71_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and71_y0);
  and_gate and_gate_h_u_cla24_and72_y0(h_u_cla24_and71_y0, h_u_cla24_and70_y0, h_u_cla24_and72_y0);
  and_gate and_gate_h_u_cla24_and73_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and73_y0);
  and_gate and_gate_h_u_cla24_and74_y0(h_u_cla24_and73_y0, h_u_cla24_and72_y0, h_u_cla24_and74_y0);
  and_gate and_gate_h_u_cla24_and75_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and75_y0);
  and_gate and_gate_h_u_cla24_and76_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and76_y0);
  and_gate and_gate_h_u_cla24_and77_y0(h_u_cla24_and76_y0, h_u_cla24_and75_y0, h_u_cla24_and77_y0);
  and_gate and_gate_h_u_cla24_and78_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and78_y0);
  and_gate and_gate_h_u_cla24_and79_y0(h_u_cla24_and78_y0, h_u_cla24_and77_y0, h_u_cla24_and79_y0);
  and_gate and_gate_h_u_cla24_and80_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and80_y0);
  and_gate and_gate_h_u_cla24_and81_y0(h_u_cla24_and80_y0, h_u_cla24_and79_y0, h_u_cla24_and81_y0);
  and_gate and_gate_h_u_cla24_and82_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and82_y0);
  and_gate and_gate_h_u_cla24_and83_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and83_y0);
  and_gate and_gate_h_u_cla24_and84_y0(h_u_cla24_and83_y0, h_u_cla24_and82_y0, h_u_cla24_and84_y0);
  and_gate and_gate_h_u_cla24_and85_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and85_y0);
  and_gate and_gate_h_u_cla24_and86_y0(h_u_cla24_and85_y0, h_u_cla24_and84_y0, h_u_cla24_and86_y0);
  and_gate and_gate_h_u_cla24_and87_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and87_y0);
  and_gate and_gate_h_u_cla24_and88_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and88_y0);
  and_gate and_gate_h_u_cla24_and89_y0(h_u_cla24_and88_y0, h_u_cla24_and87_y0, h_u_cla24_and89_y0);
  and_gate and_gate_h_u_cla24_and90_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and90_y0);
  or_gate or_gate_h_u_cla24_or15_y0(h_u_cla24_and90_y0, h_u_cla24_and65_y0, h_u_cla24_or15_y0);
  or_gate or_gate_h_u_cla24_or16_y0(h_u_cla24_or15_y0, h_u_cla24_and74_y0, h_u_cla24_or16_y0);
  or_gate or_gate_h_u_cla24_or17_y0(h_u_cla24_or16_y0, h_u_cla24_and81_y0, h_u_cla24_or17_y0);
  or_gate or_gate_h_u_cla24_or18_y0(h_u_cla24_or17_y0, h_u_cla24_and86_y0, h_u_cla24_or18_y0);
  or_gate or_gate_h_u_cla24_or19_y0(h_u_cla24_or18_y0, h_u_cla24_and89_y0, h_u_cla24_or19_y0);
  or_gate or_gate_h_u_cla24_or20_y0(h_u_cla24_pg_logic5_y1, h_u_cla24_or19_y0, h_u_cla24_or20_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic6_y0(a_6, b_6, h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_pg_logic6_y2);
  xor_gate xor_gate_h_u_cla24_xor6_y0(h_u_cla24_pg_logic6_y2, h_u_cla24_or20_y0, h_u_cla24_xor6_y0);
  and_gate and_gate_h_u_cla24_and91_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and91_y0);
  and_gate and_gate_h_u_cla24_and92_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and92_y0);
  and_gate and_gate_h_u_cla24_and93_y0(h_u_cla24_and92_y0, h_u_cla24_and91_y0, h_u_cla24_and93_y0);
  and_gate and_gate_h_u_cla24_and94_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and94_y0);
  and_gate and_gate_h_u_cla24_and95_y0(h_u_cla24_and94_y0, h_u_cla24_and93_y0, h_u_cla24_and95_y0);
  and_gate and_gate_h_u_cla24_and96_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and96_y0);
  and_gate and_gate_h_u_cla24_and97_y0(h_u_cla24_and96_y0, h_u_cla24_and95_y0, h_u_cla24_and97_y0);
  and_gate and_gate_h_u_cla24_and98_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and98_y0);
  and_gate and_gate_h_u_cla24_and99_y0(h_u_cla24_and98_y0, h_u_cla24_and97_y0, h_u_cla24_and99_y0);
  and_gate and_gate_h_u_cla24_and100_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and100_y0);
  and_gate and_gate_h_u_cla24_and101_y0(h_u_cla24_and100_y0, h_u_cla24_and99_y0, h_u_cla24_and101_y0);
  and_gate and_gate_h_u_cla24_and102_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and102_y0);
  and_gate and_gate_h_u_cla24_and103_y0(h_u_cla24_and102_y0, h_u_cla24_and101_y0, h_u_cla24_and103_y0);
  and_gate and_gate_h_u_cla24_and104_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and104_y0);
  and_gate and_gate_h_u_cla24_and105_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and105_y0);
  and_gate and_gate_h_u_cla24_and106_y0(h_u_cla24_and105_y0, h_u_cla24_and104_y0, h_u_cla24_and106_y0);
  and_gate and_gate_h_u_cla24_and107_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and107_y0);
  and_gate and_gate_h_u_cla24_and108_y0(h_u_cla24_and107_y0, h_u_cla24_and106_y0, h_u_cla24_and108_y0);
  and_gate and_gate_h_u_cla24_and109_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and109_y0);
  and_gate and_gate_h_u_cla24_and110_y0(h_u_cla24_and109_y0, h_u_cla24_and108_y0, h_u_cla24_and110_y0);
  and_gate and_gate_h_u_cla24_and111_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and111_y0);
  and_gate and_gate_h_u_cla24_and112_y0(h_u_cla24_and111_y0, h_u_cla24_and110_y0, h_u_cla24_and112_y0);
  and_gate and_gate_h_u_cla24_and113_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and113_y0);
  and_gate and_gate_h_u_cla24_and114_y0(h_u_cla24_and113_y0, h_u_cla24_and112_y0, h_u_cla24_and114_y0);
  and_gate and_gate_h_u_cla24_and115_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and115_y0);
  and_gate and_gate_h_u_cla24_and116_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and116_y0);
  and_gate and_gate_h_u_cla24_and117_y0(h_u_cla24_and116_y0, h_u_cla24_and115_y0, h_u_cla24_and117_y0);
  and_gate and_gate_h_u_cla24_and118_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and118_y0);
  and_gate and_gate_h_u_cla24_and119_y0(h_u_cla24_and118_y0, h_u_cla24_and117_y0, h_u_cla24_and119_y0);
  and_gate and_gate_h_u_cla24_and120_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and120_y0);
  and_gate and_gate_h_u_cla24_and121_y0(h_u_cla24_and120_y0, h_u_cla24_and119_y0, h_u_cla24_and121_y0);
  and_gate and_gate_h_u_cla24_and122_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and122_y0);
  and_gate and_gate_h_u_cla24_and123_y0(h_u_cla24_and122_y0, h_u_cla24_and121_y0, h_u_cla24_and123_y0);
  and_gate and_gate_h_u_cla24_and124_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and124_y0);
  and_gate and_gate_h_u_cla24_and125_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and125_y0);
  and_gate and_gate_h_u_cla24_and126_y0(h_u_cla24_and125_y0, h_u_cla24_and124_y0, h_u_cla24_and126_y0);
  and_gate and_gate_h_u_cla24_and127_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and127_y0);
  and_gate and_gate_h_u_cla24_and128_y0(h_u_cla24_and127_y0, h_u_cla24_and126_y0, h_u_cla24_and128_y0);
  and_gate and_gate_h_u_cla24_and129_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and129_y0);
  and_gate and_gate_h_u_cla24_and130_y0(h_u_cla24_and129_y0, h_u_cla24_and128_y0, h_u_cla24_and130_y0);
  and_gate and_gate_h_u_cla24_and131_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and131_y0);
  and_gate and_gate_h_u_cla24_and132_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and132_y0);
  and_gate and_gate_h_u_cla24_and133_y0(h_u_cla24_and132_y0, h_u_cla24_and131_y0, h_u_cla24_and133_y0);
  and_gate and_gate_h_u_cla24_and134_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and134_y0);
  and_gate and_gate_h_u_cla24_and135_y0(h_u_cla24_and134_y0, h_u_cla24_and133_y0, h_u_cla24_and135_y0);
  and_gate and_gate_h_u_cla24_and136_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and136_y0);
  and_gate and_gate_h_u_cla24_and137_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and137_y0);
  and_gate and_gate_h_u_cla24_and138_y0(h_u_cla24_and137_y0, h_u_cla24_and136_y0, h_u_cla24_and138_y0);
  and_gate and_gate_h_u_cla24_and139_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and139_y0);
  or_gate or_gate_h_u_cla24_or21_y0(h_u_cla24_and139_y0, h_u_cla24_and103_y0, h_u_cla24_or21_y0);
  or_gate or_gate_h_u_cla24_or22_y0(h_u_cla24_or21_y0, h_u_cla24_and114_y0, h_u_cla24_or22_y0);
  or_gate or_gate_h_u_cla24_or23_y0(h_u_cla24_or22_y0, h_u_cla24_and123_y0, h_u_cla24_or23_y0);
  or_gate or_gate_h_u_cla24_or24_y0(h_u_cla24_or23_y0, h_u_cla24_and130_y0, h_u_cla24_or24_y0);
  or_gate or_gate_h_u_cla24_or25_y0(h_u_cla24_or24_y0, h_u_cla24_and135_y0, h_u_cla24_or25_y0);
  or_gate or_gate_h_u_cla24_or26_y0(h_u_cla24_or25_y0, h_u_cla24_and138_y0, h_u_cla24_or26_y0);
  or_gate or_gate_h_u_cla24_or27_y0(h_u_cla24_pg_logic6_y1, h_u_cla24_or26_y0, h_u_cla24_or27_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic7_y0(a_7, b_7, h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_pg_logic7_y2);
  xor_gate xor_gate_h_u_cla24_xor7_y0(h_u_cla24_pg_logic7_y2, h_u_cla24_or27_y0, h_u_cla24_xor7_y0);
  and_gate and_gate_h_u_cla24_and140_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and140_y0);
  and_gate and_gate_h_u_cla24_and141_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and141_y0);
  and_gate and_gate_h_u_cla24_and142_y0(h_u_cla24_and141_y0, h_u_cla24_and140_y0, h_u_cla24_and142_y0);
  and_gate and_gate_h_u_cla24_and143_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and143_y0);
  and_gate and_gate_h_u_cla24_and144_y0(h_u_cla24_and143_y0, h_u_cla24_and142_y0, h_u_cla24_and144_y0);
  and_gate and_gate_h_u_cla24_and145_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and145_y0);
  and_gate and_gate_h_u_cla24_and146_y0(h_u_cla24_and145_y0, h_u_cla24_and144_y0, h_u_cla24_and146_y0);
  and_gate and_gate_h_u_cla24_and147_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and147_y0);
  and_gate and_gate_h_u_cla24_and148_y0(h_u_cla24_and147_y0, h_u_cla24_and146_y0, h_u_cla24_and148_y0);
  and_gate and_gate_h_u_cla24_and149_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and149_y0);
  and_gate and_gate_h_u_cla24_and150_y0(h_u_cla24_and149_y0, h_u_cla24_and148_y0, h_u_cla24_and150_y0);
  and_gate and_gate_h_u_cla24_and151_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and151_y0);
  and_gate and_gate_h_u_cla24_and152_y0(h_u_cla24_and151_y0, h_u_cla24_and150_y0, h_u_cla24_and152_y0);
  and_gate and_gate_h_u_cla24_and153_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and153_y0);
  and_gate and_gate_h_u_cla24_and154_y0(h_u_cla24_and153_y0, h_u_cla24_and152_y0, h_u_cla24_and154_y0);
  and_gate and_gate_h_u_cla24_and155_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and155_y0);
  and_gate and_gate_h_u_cla24_and156_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and156_y0);
  and_gate and_gate_h_u_cla24_and157_y0(h_u_cla24_and156_y0, h_u_cla24_and155_y0, h_u_cla24_and157_y0);
  and_gate and_gate_h_u_cla24_and158_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and158_y0);
  and_gate and_gate_h_u_cla24_and159_y0(h_u_cla24_and158_y0, h_u_cla24_and157_y0, h_u_cla24_and159_y0);
  and_gate and_gate_h_u_cla24_and160_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and160_y0);
  and_gate and_gate_h_u_cla24_and161_y0(h_u_cla24_and160_y0, h_u_cla24_and159_y0, h_u_cla24_and161_y0);
  and_gate and_gate_h_u_cla24_and162_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and162_y0);
  and_gate and_gate_h_u_cla24_and163_y0(h_u_cla24_and162_y0, h_u_cla24_and161_y0, h_u_cla24_and163_y0);
  and_gate and_gate_h_u_cla24_and164_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and164_y0);
  and_gate and_gate_h_u_cla24_and165_y0(h_u_cla24_and164_y0, h_u_cla24_and163_y0, h_u_cla24_and165_y0);
  and_gate and_gate_h_u_cla24_and166_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and166_y0);
  and_gate and_gate_h_u_cla24_and167_y0(h_u_cla24_and166_y0, h_u_cla24_and165_y0, h_u_cla24_and167_y0);
  and_gate and_gate_h_u_cla24_and168_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and168_y0);
  and_gate and_gate_h_u_cla24_and169_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and169_y0);
  and_gate and_gate_h_u_cla24_and170_y0(h_u_cla24_and169_y0, h_u_cla24_and168_y0, h_u_cla24_and170_y0);
  and_gate and_gate_h_u_cla24_and171_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and171_y0);
  and_gate and_gate_h_u_cla24_and172_y0(h_u_cla24_and171_y0, h_u_cla24_and170_y0, h_u_cla24_and172_y0);
  and_gate and_gate_h_u_cla24_and173_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and173_y0);
  and_gate and_gate_h_u_cla24_and174_y0(h_u_cla24_and173_y0, h_u_cla24_and172_y0, h_u_cla24_and174_y0);
  and_gate and_gate_h_u_cla24_and175_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and175_y0);
  and_gate and_gate_h_u_cla24_and176_y0(h_u_cla24_and175_y0, h_u_cla24_and174_y0, h_u_cla24_and176_y0);
  and_gate and_gate_h_u_cla24_and177_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and177_y0);
  and_gate and_gate_h_u_cla24_and178_y0(h_u_cla24_and177_y0, h_u_cla24_and176_y0, h_u_cla24_and178_y0);
  and_gate and_gate_h_u_cla24_and179_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and179_y0);
  and_gate and_gate_h_u_cla24_and180_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and180_y0);
  and_gate and_gate_h_u_cla24_and181_y0(h_u_cla24_and180_y0, h_u_cla24_and179_y0, h_u_cla24_and181_y0);
  and_gate and_gate_h_u_cla24_and182_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and182_y0);
  and_gate and_gate_h_u_cla24_and183_y0(h_u_cla24_and182_y0, h_u_cla24_and181_y0, h_u_cla24_and183_y0);
  and_gate and_gate_h_u_cla24_and184_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and184_y0);
  and_gate and_gate_h_u_cla24_and185_y0(h_u_cla24_and184_y0, h_u_cla24_and183_y0, h_u_cla24_and185_y0);
  and_gate and_gate_h_u_cla24_and186_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and186_y0);
  and_gate and_gate_h_u_cla24_and187_y0(h_u_cla24_and186_y0, h_u_cla24_and185_y0, h_u_cla24_and187_y0);
  and_gate and_gate_h_u_cla24_and188_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and188_y0);
  and_gate and_gate_h_u_cla24_and189_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and189_y0);
  and_gate and_gate_h_u_cla24_and190_y0(h_u_cla24_and189_y0, h_u_cla24_and188_y0, h_u_cla24_and190_y0);
  and_gate and_gate_h_u_cla24_and191_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and191_y0);
  and_gate and_gate_h_u_cla24_and192_y0(h_u_cla24_and191_y0, h_u_cla24_and190_y0, h_u_cla24_and192_y0);
  and_gate and_gate_h_u_cla24_and193_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and193_y0);
  and_gate and_gate_h_u_cla24_and194_y0(h_u_cla24_and193_y0, h_u_cla24_and192_y0, h_u_cla24_and194_y0);
  and_gate and_gate_h_u_cla24_and195_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and195_y0);
  and_gate and_gate_h_u_cla24_and196_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and196_y0);
  and_gate and_gate_h_u_cla24_and197_y0(h_u_cla24_and196_y0, h_u_cla24_and195_y0, h_u_cla24_and197_y0);
  and_gate and_gate_h_u_cla24_and198_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and198_y0);
  and_gate and_gate_h_u_cla24_and199_y0(h_u_cla24_and198_y0, h_u_cla24_and197_y0, h_u_cla24_and199_y0);
  and_gate and_gate_h_u_cla24_and200_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and200_y0);
  and_gate and_gate_h_u_cla24_and201_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and201_y0);
  and_gate and_gate_h_u_cla24_and202_y0(h_u_cla24_and201_y0, h_u_cla24_and200_y0, h_u_cla24_and202_y0);
  and_gate and_gate_h_u_cla24_and203_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and203_y0);
  or_gate or_gate_h_u_cla24_or28_y0(h_u_cla24_and203_y0, h_u_cla24_and154_y0, h_u_cla24_or28_y0);
  or_gate or_gate_h_u_cla24_or29_y0(h_u_cla24_or28_y0, h_u_cla24_and167_y0, h_u_cla24_or29_y0);
  or_gate or_gate_h_u_cla24_or30_y0(h_u_cla24_or29_y0, h_u_cla24_and178_y0, h_u_cla24_or30_y0);
  or_gate or_gate_h_u_cla24_or31_y0(h_u_cla24_or30_y0, h_u_cla24_and187_y0, h_u_cla24_or31_y0);
  or_gate or_gate_h_u_cla24_or32_y0(h_u_cla24_or31_y0, h_u_cla24_and194_y0, h_u_cla24_or32_y0);
  or_gate or_gate_h_u_cla24_or33_y0(h_u_cla24_or32_y0, h_u_cla24_and199_y0, h_u_cla24_or33_y0);
  or_gate or_gate_h_u_cla24_or34_y0(h_u_cla24_or33_y0, h_u_cla24_and202_y0, h_u_cla24_or34_y0);
  or_gate or_gate_h_u_cla24_or35_y0(h_u_cla24_pg_logic7_y1, h_u_cla24_or34_y0, h_u_cla24_or35_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic8_y0(a_8, b_8, h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_pg_logic8_y2);
  xor_gate xor_gate_h_u_cla24_xor8_y0(h_u_cla24_pg_logic8_y2, h_u_cla24_or35_y0, h_u_cla24_xor8_y0);
  and_gate and_gate_h_u_cla24_and204_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and204_y0);
  and_gate and_gate_h_u_cla24_and205_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and205_y0);
  and_gate and_gate_h_u_cla24_and206_y0(h_u_cla24_and205_y0, h_u_cla24_and204_y0, h_u_cla24_and206_y0);
  and_gate and_gate_h_u_cla24_and207_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and207_y0);
  and_gate and_gate_h_u_cla24_and208_y0(h_u_cla24_and207_y0, h_u_cla24_and206_y0, h_u_cla24_and208_y0);
  and_gate and_gate_h_u_cla24_and209_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and209_y0);
  and_gate and_gate_h_u_cla24_and210_y0(h_u_cla24_and209_y0, h_u_cla24_and208_y0, h_u_cla24_and210_y0);
  and_gate and_gate_h_u_cla24_and211_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and211_y0);
  and_gate and_gate_h_u_cla24_and212_y0(h_u_cla24_and211_y0, h_u_cla24_and210_y0, h_u_cla24_and212_y0);
  and_gate and_gate_h_u_cla24_and213_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and213_y0);
  and_gate and_gate_h_u_cla24_and214_y0(h_u_cla24_and213_y0, h_u_cla24_and212_y0, h_u_cla24_and214_y0);
  and_gate and_gate_h_u_cla24_and215_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and215_y0);
  and_gate and_gate_h_u_cla24_and216_y0(h_u_cla24_and215_y0, h_u_cla24_and214_y0, h_u_cla24_and216_y0);
  and_gate and_gate_h_u_cla24_and217_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and217_y0);
  and_gate and_gate_h_u_cla24_and218_y0(h_u_cla24_and217_y0, h_u_cla24_and216_y0, h_u_cla24_and218_y0);
  and_gate and_gate_h_u_cla24_and219_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and219_y0);
  and_gate and_gate_h_u_cla24_and220_y0(h_u_cla24_and219_y0, h_u_cla24_and218_y0, h_u_cla24_and220_y0);
  and_gate and_gate_h_u_cla24_and221_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and221_y0);
  and_gate and_gate_h_u_cla24_and222_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and222_y0);
  and_gate and_gate_h_u_cla24_and223_y0(h_u_cla24_and222_y0, h_u_cla24_and221_y0, h_u_cla24_and223_y0);
  and_gate and_gate_h_u_cla24_and224_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and224_y0);
  and_gate and_gate_h_u_cla24_and225_y0(h_u_cla24_and224_y0, h_u_cla24_and223_y0, h_u_cla24_and225_y0);
  and_gate and_gate_h_u_cla24_and226_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and226_y0);
  and_gate and_gate_h_u_cla24_and227_y0(h_u_cla24_and226_y0, h_u_cla24_and225_y0, h_u_cla24_and227_y0);
  and_gate and_gate_h_u_cla24_and228_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and228_y0);
  and_gate and_gate_h_u_cla24_and229_y0(h_u_cla24_and228_y0, h_u_cla24_and227_y0, h_u_cla24_and229_y0);
  and_gate and_gate_h_u_cla24_and230_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and230_y0);
  and_gate and_gate_h_u_cla24_and231_y0(h_u_cla24_and230_y0, h_u_cla24_and229_y0, h_u_cla24_and231_y0);
  and_gate and_gate_h_u_cla24_and232_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and232_y0);
  and_gate and_gate_h_u_cla24_and233_y0(h_u_cla24_and232_y0, h_u_cla24_and231_y0, h_u_cla24_and233_y0);
  and_gate and_gate_h_u_cla24_and234_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and234_y0);
  and_gate and_gate_h_u_cla24_and235_y0(h_u_cla24_and234_y0, h_u_cla24_and233_y0, h_u_cla24_and235_y0);
  and_gate and_gate_h_u_cla24_and236_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and236_y0);
  and_gate and_gate_h_u_cla24_and237_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and237_y0);
  and_gate and_gate_h_u_cla24_and238_y0(h_u_cla24_and237_y0, h_u_cla24_and236_y0, h_u_cla24_and238_y0);
  and_gate and_gate_h_u_cla24_and239_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and239_y0);
  and_gate and_gate_h_u_cla24_and240_y0(h_u_cla24_and239_y0, h_u_cla24_and238_y0, h_u_cla24_and240_y0);
  and_gate and_gate_h_u_cla24_and241_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and241_y0);
  and_gate and_gate_h_u_cla24_and242_y0(h_u_cla24_and241_y0, h_u_cla24_and240_y0, h_u_cla24_and242_y0);
  and_gate and_gate_h_u_cla24_and243_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and243_y0);
  and_gate and_gate_h_u_cla24_and244_y0(h_u_cla24_and243_y0, h_u_cla24_and242_y0, h_u_cla24_and244_y0);
  and_gate and_gate_h_u_cla24_and245_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and245_y0);
  and_gate and_gate_h_u_cla24_and246_y0(h_u_cla24_and245_y0, h_u_cla24_and244_y0, h_u_cla24_and246_y0);
  and_gate and_gate_h_u_cla24_and247_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and247_y0);
  and_gate and_gate_h_u_cla24_and248_y0(h_u_cla24_and247_y0, h_u_cla24_and246_y0, h_u_cla24_and248_y0);
  and_gate and_gate_h_u_cla24_and249_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and249_y0);
  and_gate and_gate_h_u_cla24_and250_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and250_y0);
  and_gate and_gate_h_u_cla24_and251_y0(h_u_cla24_and250_y0, h_u_cla24_and249_y0, h_u_cla24_and251_y0);
  and_gate and_gate_h_u_cla24_and252_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and252_y0);
  and_gate and_gate_h_u_cla24_and253_y0(h_u_cla24_and252_y0, h_u_cla24_and251_y0, h_u_cla24_and253_y0);
  and_gate and_gate_h_u_cla24_and254_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and254_y0);
  and_gate and_gate_h_u_cla24_and255_y0(h_u_cla24_and254_y0, h_u_cla24_and253_y0, h_u_cla24_and255_y0);
  and_gate and_gate_h_u_cla24_and256_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and256_y0);
  and_gate and_gate_h_u_cla24_and257_y0(h_u_cla24_and256_y0, h_u_cla24_and255_y0, h_u_cla24_and257_y0);
  and_gate and_gate_h_u_cla24_and258_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and258_y0);
  and_gate and_gate_h_u_cla24_and259_y0(h_u_cla24_and258_y0, h_u_cla24_and257_y0, h_u_cla24_and259_y0);
  and_gate and_gate_h_u_cla24_and260_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and260_y0);
  and_gate and_gate_h_u_cla24_and261_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and261_y0);
  and_gate and_gate_h_u_cla24_and262_y0(h_u_cla24_and261_y0, h_u_cla24_and260_y0, h_u_cla24_and262_y0);
  and_gate and_gate_h_u_cla24_and263_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and263_y0);
  and_gate and_gate_h_u_cla24_and264_y0(h_u_cla24_and263_y0, h_u_cla24_and262_y0, h_u_cla24_and264_y0);
  and_gate and_gate_h_u_cla24_and265_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and265_y0);
  and_gate and_gate_h_u_cla24_and266_y0(h_u_cla24_and265_y0, h_u_cla24_and264_y0, h_u_cla24_and266_y0);
  and_gate and_gate_h_u_cla24_and267_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and267_y0);
  and_gate and_gate_h_u_cla24_and268_y0(h_u_cla24_and267_y0, h_u_cla24_and266_y0, h_u_cla24_and268_y0);
  and_gate and_gate_h_u_cla24_and269_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and269_y0);
  and_gate and_gate_h_u_cla24_and270_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and270_y0);
  and_gate and_gate_h_u_cla24_and271_y0(h_u_cla24_and270_y0, h_u_cla24_and269_y0, h_u_cla24_and271_y0);
  and_gate and_gate_h_u_cla24_and272_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and272_y0);
  and_gate and_gate_h_u_cla24_and273_y0(h_u_cla24_and272_y0, h_u_cla24_and271_y0, h_u_cla24_and273_y0);
  and_gate and_gate_h_u_cla24_and274_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and274_y0);
  and_gate and_gate_h_u_cla24_and275_y0(h_u_cla24_and274_y0, h_u_cla24_and273_y0, h_u_cla24_and275_y0);
  and_gate and_gate_h_u_cla24_and276_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and276_y0);
  and_gate and_gate_h_u_cla24_and277_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and277_y0);
  and_gate and_gate_h_u_cla24_and278_y0(h_u_cla24_and277_y0, h_u_cla24_and276_y0, h_u_cla24_and278_y0);
  and_gate and_gate_h_u_cla24_and279_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and279_y0);
  and_gate and_gate_h_u_cla24_and280_y0(h_u_cla24_and279_y0, h_u_cla24_and278_y0, h_u_cla24_and280_y0);
  and_gate and_gate_h_u_cla24_and281_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and281_y0);
  and_gate and_gate_h_u_cla24_and282_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and282_y0);
  and_gate and_gate_h_u_cla24_and283_y0(h_u_cla24_and282_y0, h_u_cla24_and281_y0, h_u_cla24_and283_y0);
  and_gate and_gate_h_u_cla24_and284_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and284_y0);
  or_gate or_gate_h_u_cla24_or36_y0(h_u_cla24_and284_y0, h_u_cla24_and220_y0, h_u_cla24_or36_y0);
  or_gate or_gate_h_u_cla24_or37_y0(h_u_cla24_or36_y0, h_u_cla24_and235_y0, h_u_cla24_or37_y0);
  or_gate or_gate_h_u_cla24_or38_y0(h_u_cla24_or37_y0, h_u_cla24_and248_y0, h_u_cla24_or38_y0);
  or_gate or_gate_h_u_cla24_or39_y0(h_u_cla24_or38_y0, h_u_cla24_and259_y0, h_u_cla24_or39_y0);
  or_gate or_gate_h_u_cla24_or40_y0(h_u_cla24_or39_y0, h_u_cla24_and268_y0, h_u_cla24_or40_y0);
  or_gate or_gate_h_u_cla24_or41_y0(h_u_cla24_or40_y0, h_u_cla24_and275_y0, h_u_cla24_or41_y0);
  or_gate or_gate_h_u_cla24_or42_y0(h_u_cla24_or41_y0, h_u_cla24_and280_y0, h_u_cla24_or42_y0);
  or_gate or_gate_h_u_cla24_or43_y0(h_u_cla24_or42_y0, h_u_cla24_and283_y0, h_u_cla24_or43_y0);
  or_gate or_gate_h_u_cla24_or44_y0(h_u_cla24_pg_logic8_y1, h_u_cla24_or43_y0, h_u_cla24_or44_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic9_y0(a_9, b_9, h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_pg_logic9_y2);
  xor_gate xor_gate_h_u_cla24_xor9_y0(h_u_cla24_pg_logic9_y2, h_u_cla24_or44_y0, h_u_cla24_xor9_y0);
  and_gate and_gate_h_u_cla24_and285_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and285_y0);
  and_gate and_gate_h_u_cla24_and286_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and286_y0);
  and_gate and_gate_h_u_cla24_and287_y0(h_u_cla24_and286_y0, h_u_cla24_and285_y0, h_u_cla24_and287_y0);
  and_gate and_gate_h_u_cla24_and288_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and288_y0);
  and_gate and_gate_h_u_cla24_and289_y0(h_u_cla24_and288_y0, h_u_cla24_and287_y0, h_u_cla24_and289_y0);
  and_gate and_gate_h_u_cla24_and290_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and290_y0);
  and_gate and_gate_h_u_cla24_and291_y0(h_u_cla24_and290_y0, h_u_cla24_and289_y0, h_u_cla24_and291_y0);
  and_gate and_gate_h_u_cla24_and292_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and292_y0);
  and_gate and_gate_h_u_cla24_and293_y0(h_u_cla24_and292_y0, h_u_cla24_and291_y0, h_u_cla24_and293_y0);
  and_gate and_gate_h_u_cla24_and294_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and294_y0);
  and_gate and_gate_h_u_cla24_and295_y0(h_u_cla24_and294_y0, h_u_cla24_and293_y0, h_u_cla24_and295_y0);
  and_gate and_gate_h_u_cla24_and296_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and296_y0);
  and_gate and_gate_h_u_cla24_and297_y0(h_u_cla24_and296_y0, h_u_cla24_and295_y0, h_u_cla24_and297_y0);
  and_gate and_gate_h_u_cla24_and298_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and298_y0);
  and_gate and_gate_h_u_cla24_and299_y0(h_u_cla24_and298_y0, h_u_cla24_and297_y0, h_u_cla24_and299_y0);
  and_gate and_gate_h_u_cla24_and300_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and300_y0);
  and_gate and_gate_h_u_cla24_and301_y0(h_u_cla24_and300_y0, h_u_cla24_and299_y0, h_u_cla24_and301_y0);
  and_gate and_gate_h_u_cla24_and302_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and302_y0);
  and_gate and_gate_h_u_cla24_and303_y0(h_u_cla24_and302_y0, h_u_cla24_and301_y0, h_u_cla24_and303_y0);
  and_gate and_gate_h_u_cla24_and304_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and304_y0);
  and_gate and_gate_h_u_cla24_and305_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and305_y0);
  and_gate and_gate_h_u_cla24_and306_y0(h_u_cla24_and305_y0, h_u_cla24_and304_y0, h_u_cla24_and306_y0);
  and_gate and_gate_h_u_cla24_and307_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and307_y0);
  and_gate and_gate_h_u_cla24_and308_y0(h_u_cla24_and307_y0, h_u_cla24_and306_y0, h_u_cla24_and308_y0);
  and_gate and_gate_h_u_cla24_and309_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and309_y0);
  and_gate and_gate_h_u_cla24_and310_y0(h_u_cla24_and309_y0, h_u_cla24_and308_y0, h_u_cla24_and310_y0);
  and_gate and_gate_h_u_cla24_and311_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and311_y0);
  and_gate and_gate_h_u_cla24_and312_y0(h_u_cla24_and311_y0, h_u_cla24_and310_y0, h_u_cla24_and312_y0);
  and_gate and_gate_h_u_cla24_and313_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and313_y0);
  and_gate and_gate_h_u_cla24_and314_y0(h_u_cla24_and313_y0, h_u_cla24_and312_y0, h_u_cla24_and314_y0);
  and_gate and_gate_h_u_cla24_and315_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and315_y0);
  and_gate and_gate_h_u_cla24_and316_y0(h_u_cla24_and315_y0, h_u_cla24_and314_y0, h_u_cla24_and316_y0);
  and_gate and_gate_h_u_cla24_and317_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and317_y0);
  and_gate and_gate_h_u_cla24_and318_y0(h_u_cla24_and317_y0, h_u_cla24_and316_y0, h_u_cla24_and318_y0);
  and_gate and_gate_h_u_cla24_and319_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and319_y0);
  and_gate and_gate_h_u_cla24_and320_y0(h_u_cla24_and319_y0, h_u_cla24_and318_y0, h_u_cla24_and320_y0);
  and_gate and_gate_h_u_cla24_and321_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and321_y0);
  and_gate and_gate_h_u_cla24_and322_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and322_y0);
  and_gate and_gate_h_u_cla24_and323_y0(h_u_cla24_and322_y0, h_u_cla24_and321_y0, h_u_cla24_and323_y0);
  and_gate and_gate_h_u_cla24_and324_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and324_y0);
  and_gate and_gate_h_u_cla24_and325_y0(h_u_cla24_and324_y0, h_u_cla24_and323_y0, h_u_cla24_and325_y0);
  and_gate and_gate_h_u_cla24_and326_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and326_y0);
  and_gate and_gate_h_u_cla24_and327_y0(h_u_cla24_and326_y0, h_u_cla24_and325_y0, h_u_cla24_and327_y0);
  and_gate and_gate_h_u_cla24_and328_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and328_y0);
  and_gate and_gate_h_u_cla24_and329_y0(h_u_cla24_and328_y0, h_u_cla24_and327_y0, h_u_cla24_and329_y0);
  and_gate and_gate_h_u_cla24_and330_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and330_y0);
  and_gate and_gate_h_u_cla24_and331_y0(h_u_cla24_and330_y0, h_u_cla24_and329_y0, h_u_cla24_and331_y0);
  and_gate and_gate_h_u_cla24_and332_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and332_y0);
  and_gate and_gate_h_u_cla24_and333_y0(h_u_cla24_and332_y0, h_u_cla24_and331_y0, h_u_cla24_and333_y0);
  and_gate and_gate_h_u_cla24_and334_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and334_y0);
  and_gate and_gate_h_u_cla24_and335_y0(h_u_cla24_and334_y0, h_u_cla24_and333_y0, h_u_cla24_and335_y0);
  and_gate and_gate_h_u_cla24_and336_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and336_y0);
  and_gate and_gate_h_u_cla24_and337_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and337_y0);
  and_gate and_gate_h_u_cla24_and338_y0(h_u_cla24_and337_y0, h_u_cla24_and336_y0, h_u_cla24_and338_y0);
  and_gate and_gate_h_u_cla24_and339_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and339_y0);
  and_gate and_gate_h_u_cla24_and340_y0(h_u_cla24_and339_y0, h_u_cla24_and338_y0, h_u_cla24_and340_y0);
  and_gate and_gate_h_u_cla24_and341_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and341_y0);
  and_gate and_gate_h_u_cla24_and342_y0(h_u_cla24_and341_y0, h_u_cla24_and340_y0, h_u_cla24_and342_y0);
  and_gate and_gate_h_u_cla24_and343_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and343_y0);
  and_gate and_gate_h_u_cla24_and344_y0(h_u_cla24_and343_y0, h_u_cla24_and342_y0, h_u_cla24_and344_y0);
  and_gate and_gate_h_u_cla24_and345_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and345_y0);
  and_gate and_gate_h_u_cla24_and346_y0(h_u_cla24_and345_y0, h_u_cla24_and344_y0, h_u_cla24_and346_y0);
  and_gate and_gate_h_u_cla24_and347_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and347_y0);
  and_gate and_gate_h_u_cla24_and348_y0(h_u_cla24_and347_y0, h_u_cla24_and346_y0, h_u_cla24_and348_y0);
  and_gate and_gate_h_u_cla24_and349_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and349_y0);
  and_gate and_gate_h_u_cla24_and350_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and350_y0);
  and_gate and_gate_h_u_cla24_and351_y0(h_u_cla24_and350_y0, h_u_cla24_and349_y0, h_u_cla24_and351_y0);
  and_gate and_gate_h_u_cla24_and352_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and352_y0);
  and_gate and_gate_h_u_cla24_and353_y0(h_u_cla24_and352_y0, h_u_cla24_and351_y0, h_u_cla24_and353_y0);
  and_gate and_gate_h_u_cla24_and354_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and354_y0);
  and_gate and_gate_h_u_cla24_and355_y0(h_u_cla24_and354_y0, h_u_cla24_and353_y0, h_u_cla24_and355_y0);
  and_gate and_gate_h_u_cla24_and356_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and356_y0);
  and_gate and_gate_h_u_cla24_and357_y0(h_u_cla24_and356_y0, h_u_cla24_and355_y0, h_u_cla24_and357_y0);
  and_gate and_gate_h_u_cla24_and358_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and358_y0);
  and_gate and_gate_h_u_cla24_and359_y0(h_u_cla24_and358_y0, h_u_cla24_and357_y0, h_u_cla24_and359_y0);
  and_gate and_gate_h_u_cla24_and360_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and360_y0);
  and_gate and_gate_h_u_cla24_and361_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and361_y0);
  and_gate and_gate_h_u_cla24_and362_y0(h_u_cla24_and361_y0, h_u_cla24_and360_y0, h_u_cla24_and362_y0);
  and_gate and_gate_h_u_cla24_and363_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and363_y0);
  and_gate and_gate_h_u_cla24_and364_y0(h_u_cla24_and363_y0, h_u_cla24_and362_y0, h_u_cla24_and364_y0);
  and_gate and_gate_h_u_cla24_and365_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and365_y0);
  and_gate and_gate_h_u_cla24_and366_y0(h_u_cla24_and365_y0, h_u_cla24_and364_y0, h_u_cla24_and366_y0);
  and_gate and_gate_h_u_cla24_and367_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and367_y0);
  and_gate and_gate_h_u_cla24_and368_y0(h_u_cla24_and367_y0, h_u_cla24_and366_y0, h_u_cla24_and368_y0);
  and_gate and_gate_h_u_cla24_and369_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and369_y0);
  and_gate and_gate_h_u_cla24_and370_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and370_y0);
  and_gate and_gate_h_u_cla24_and371_y0(h_u_cla24_and370_y0, h_u_cla24_and369_y0, h_u_cla24_and371_y0);
  and_gate and_gate_h_u_cla24_and372_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and372_y0);
  and_gate and_gate_h_u_cla24_and373_y0(h_u_cla24_and372_y0, h_u_cla24_and371_y0, h_u_cla24_and373_y0);
  and_gate and_gate_h_u_cla24_and374_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and374_y0);
  and_gate and_gate_h_u_cla24_and375_y0(h_u_cla24_and374_y0, h_u_cla24_and373_y0, h_u_cla24_and375_y0);
  and_gate and_gate_h_u_cla24_and376_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and376_y0);
  and_gate and_gate_h_u_cla24_and377_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and377_y0);
  and_gate and_gate_h_u_cla24_and378_y0(h_u_cla24_and377_y0, h_u_cla24_and376_y0, h_u_cla24_and378_y0);
  and_gate and_gate_h_u_cla24_and379_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and379_y0);
  and_gate and_gate_h_u_cla24_and380_y0(h_u_cla24_and379_y0, h_u_cla24_and378_y0, h_u_cla24_and380_y0);
  and_gate and_gate_h_u_cla24_and381_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and381_y0);
  and_gate and_gate_h_u_cla24_and382_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and382_y0);
  and_gate and_gate_h_u_cla24_and383_y0(h_u_cla24_and382_y0, h_u_cla24_and381_y0, h_u_cla24_and383_y0);
  and_gate and_gate_h_u_cla24_and384_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and384_y0);
  or_gate or_gate_h_u_cla24_or45_y0(h_u_cla24_and384_y0, h_u_cla24_and303_y0, h_u_cla24_or45_y0);
  or_gate or_gate_h_u_cla24_or46_y0(h_u_cla24_or45_y0, h_u_cla24_and320_y0, h_u_cla24_or46_y0);
  or_gate or_gate_h_u_cla24_or47_y0(h_u_cla24_or46_y0, h_u_cla24_and335_y0, h_u_cla24_or47_y0);
  or_gate or_gate_h_u_cla24_or48_y0(h_u_cla24_or47_y0, h_u_cla24_and348_y0, h_u_cla24_or48_y0);
  or_gate or_gate_h_u_cla24_or49_y0(h_u_cla24_or48_y0, h_u_cla24_and359_y0, h_u_cla24_or49_y0);
  or_gate or_gate_h_u_cla24_or50_y0(h_u_cla24_or49_y0, h_u_cla24_and368_y0, h_u_cla24_or50_y0);
  or_gate or_gate_h_u_cla24_or51_y0(h_u_cla24_or50_y0, h_u_cla24_and375_y0, h_u_cla24_or51_y0);
  or_gate or_gate_h_u_cla24_or52_y0(h_u_cla24_or51_y0, h_u_cla24_and380_y0, h_u_cla24_or52_y0);
  or_gate or_gate_h_u_cla24_or53_y0(h_u_cla24_or52_y0, h_u_cla24_and383_y0, h_u_cla24_or53_y0);
  or_gate or_gate_h_u_cla24_or54_y0(h_u_cla24_pg_logic9_y1, h_u_cla24_or53_y0, h_u_cla24_or54_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic10_y0(a_10, b_10, h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_pg_logic10_y2);
  xor_gate xor_gate_h_u_cla24_xor10_y0(h_u_cla24_pg_logic10_y2, h_u_cla24_or54_y0, h_u_cla24_xor10_y0);
  and_gate and_gate_h_u_cla24_and385_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and385_y0);
  and_gate and_gate_h_u_cla24_and386_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and386_y0);
  and_gate and_gate_h_u_cla24_and387_y0(h_u_cla24_and386_y0, h_u_cla24_and385_y0, h_u_cla24_and387_y0);
  and_gate and_gate_h_u_cla24_and388_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and388_y0);
  and_gate and_gate_h_u_cla24_and389_y0(h_u_cla24_and388_y0, h_u_cla24_and387_y0, h_u_cla24_and389_y0);
  and_gate and_gate_h_u_cla24_and390_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and390_y0);
  and_gate and_gate_h_u_cla24_and391_y0(h_u_cla24_and390_y0, h_u_cla24_and389_y0, h_u_cla24_and391_y0);
  and_gate and_gate_h_u_cla24_and392_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and392_y0);
  and_gate and_gate_h_u_cla24_and393_y0(h_u_cla24_and392_y0, h_u_cla24_and391_y0, h_u_cla24_and393_y0);
  and_gate and_gate_h_u_cla24_and394_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and394_y0);
  and_gate and_gate_h_u_cla24_and395_y0(h_u_cla24_and394_y0, h_u_cla24_and393_y0, h_u_cla24_and395_y0);
  and_gate and_gate_h_u_cla24_and396_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and396_y0);
  and_gate and_gate_h_u_cla24_and397_y0(h_u_cla24_and396_y0, h_u_cla24_and395_y0, h_u_cla24_and397_y0);
  and_gate and_gate_h_u_cla24_and398_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and398_y0);
  and_gate and_gate_h_u_cla24_and399_y0(h_u_cla24_and398_y0, h_u_cla24_and397_y0, h_u_cla24_and399_y0);
  and_gate and_gate_h_u_cla24_and400_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and400_y0);
  and_gate and_gate_h_u_cla24_and401_y0(h_u_cla24_and400_y0, h_u_cla24_and399_y0, h_u_cla24_and401_y0);
  and_gate and_gate_h_u_cla24_and402_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and402_y0);
  and_gate and_gate_h_u_cla24_and403_y0(h_u_cla24_and402_y0, h_u_cla24_and401_y0, h_u_cla24_and403_y0);
  and_gate and_gate_h_u_cla24_and404_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and404_y0);
  and_gate and_gate_h_u_cla24_and405_y0(h_u_cla24_and404_y0, h_u_cla24_and403_y0, h_u_cla24_and405_y0);
  and_gate and_gate_h_u_cla24_and406_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and406_y0);
  and_gate and_gate_h_u_cla24_and407_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and407_y0);
  and_gate and_gate_h_u_cla24_and408_y0(h_u_cla24_and407_y0, h_u_cla24_and406_y0, h_u_cla24_and408_y0);
  and_gate and_gate_h_u_cla24_and409_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and409_y0);
  and_gate and_gate_h_u_cla24_and410_y0(h_u_cla24_and409_y0, h_u_cla24_and408_y0, h_u_cla24_and410_y0);
  and_gate and_gate_h_u_cla24_and411_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and411_y0);
  and_gate and_gate_h_u_cla24_and412_y0(h_u_cla24_and411_y0, h_u_cla24_and410_y0, h_u_cla24_and412_y0);
  and_gate and_gate_h_u_cla24_and413_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and413_y0);
  and_gate and_gate_h_u_cla24_and414_y0(h_u_cla24_and413_y0, h_u_cla24_and412_y0, h_u_cla24_and414_y0);
  and_gate and_gate_h_u_cla24_and415_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and415_y0);
  and_gate and_gate_h_u_cla24_and416_y0(h_u_cla24_and415_y0, h_u_cla24_and414_y0, h_u_cla24_and416_y0);
  and_gate and_gate_h_u_cla24_and417_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and417_y0);
  and_gate and_gate_h_u_cla24_and418_y0(h_u_cla24_and417_y0, h_u_cla24_and416_y0, h_u_cla24_and418_y0);
  and_gate and_gate_h_u_cla24_and419_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and419_y0);
  and_gate and_gate_h_u_cla24_and420_y0(h_u_cla24_and419_y0, h_u_cla24_and418_y0, h_u_cla24_and420_y0);
  and_gate and_gate_h_u_cla24_and421_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and421_y0);
  and_gate and_gate_h_u_cla24_and422_y0(h_u_cla24_and421_y0, h_u_cla24_and420_y0, h_u_cla24_and422_y0);
  and_gate and_gate_h_u_cla24_and423_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and423_y0);
  and_gate and_gate_h_u_cla24_and424_y0(h_u_cla24_and423_y0, h_u_cla24_and422_y0, h_u_cla24_and424_y0);
  and_gate and_gate_h_u_cla24_and425_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and425_y0);
  and_gate and_gate_h_u_cla24_and426_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and426_y0);
  and_gate and_gate_h_u_cla24_and427_y0(h_u_cla24_and426_y0, h_u_cla24_and425_y0, h_u_cla24_and427_y0);
  and_gate and_gate_h_u_cla24_and428_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and428_y0);
  and_gate and_gate_h_u_cla24_and429_y0(h_u_cla24_and428_y0, h_u_cla24_and427_y0, h_u_cla24_and429_y0);
  and_gate and_gate_h_u_cla24_and430_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and430_y0);
  and_gate and_gate_h_u_cla24_and431_y0(h_u_cla24_and430_y0, h_u_cla24_and429_y0, h_u_cla24_and431_y0);
  and_gate and_gate_h_u_cla24_and432_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and432_y0);
  and_gate and_gate_h_u_cla24_and433_y0(h_u_cla24_and432_y0, h_u_cla24_and431_y0, h_u_cla24_and433_y0);
  and_gate and_gate_h_u_cla24_and434_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and434_y0);
  and_gate and_gate_h_u_cla24_and435_y0(h_u_cla24_and434_y0, h_u_cla24_and433_y0, h_u_cla24_and435_y0);
  and_gate and_gate_h_u_cla24_and436_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and436_y0);
  and_gate and_gate_h_u_cla24_and437_y0(h_u_cla24_and436_y0, h_u_cla24_and435_y0, h_u_cla24_and437_y0);
  and_gate and_gate_h_u_cla24_and438_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and438_y0);
  and_gate and_gate_h_u_cla24_and439_y0(h_u_cla24_and438_y0, h_u_cla24_and437_y0, h_u_cla24_and439_y0);
  and_gate and_gate_h_u_cla24_and440_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and440_y0);
  and_gate and_gate_h_u_cla24_and441_y0(h_u_cla24_and440_y0, h_u_cla24_and439_y0, h_u_cla24_and441_y0);
  and_gate and_gate_h_u_cla24_and442_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and442_y0);
  and_gate and_gate_h_u_cla24_and443_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and443_y0);
  and_gate and_gate_h_u_cla24_and444_y0(h_u_cla24_and443_y0, h_u_cla24_and442_y0, h_u_cla24_and444_y0);
  and_gate and_gate_h_u_cla24_and445_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and445_y0);
  and_gate and_gate_h_u_cla24_and446_y0(h_u_cla24_and445_y0, h_u_cla24_and444_y0, h_u_cla24_and446_y0);
  and_gate and_gate_h_u_cla24_and447_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and447_y0);
  and_gate and_gate_h_u_cla24_and448_y0(h_u_cla24_and447_y0, h_u_cla24_and446_y0, h_u_cla24_and448_y0);
  and_gate and_gate_h_u_cla24_and449_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and449_y0);
  and_gate and_gate_h_u_cla24_and450_y0(h_u_cla24_and449_y0, h_u_cla24_and448_y0, h_u_cla24_and450_y0);
  and_gate and_gate_h_u_cla24_and451_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and451_y0);
  and_gate and_gate_h_u_cla24_and452_y0(h_u_cla24_and451_y0, h_u_cla24_and450_y0, h_u_cla24_and452_y0);
  and_gate and_gate_h_u_cla24_and453_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and453_y0);
  and_gate and_gate_h_u_cla24_and454_y0(h_u_cla24_and453_y0, h_u_cla24_and452_y0, h_u_cla24_and454_y0);
  and_gate and_gate_h_u_cla24_and455_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and455_y0);
  and_gate and_gate_h_u_cla24_and456_y0(h_u_cla24_and455_y0, h_u_cla24_and454_y0, h_u_cla24_and456_y0);
  and_gate and_gate_h_u_cla24_and457_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and457_y0);
  and_gate and_gate_h_u_cla24_and458_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and458_y0);
  and_gate and_gate_h_u_cla24_and459_y0(h_u_cla24_and458_y0, h_u_cla24_and457_y0, h_u_cla24_and459_y0);
  and_gate and_gate_h_u_cla24_and460_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and460_y0);
  and_gate and_gate_h_u_cla24_and461_y0(h_u_cla24_and460_y0, h_u_cla24_and459_y0, h_u_cla24_and461_y0);
  and_gate and_gate_h_u_cla24_and462_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and462_y0);
  and_gate and_gate_h_u_cla24_and463_y0(h_u_cla24_and462_y0, h_u_cla24_and461_y0, h_u_cla24_and463_y0);
  and_gate and_gate_h_u_cla24_and464_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and464_y0);
  and_gate and_gate_h_u_cla24_and465_y0(h_u_cla24_and464_y0, h_u_cla24_and463_y0, h_u_cla24_and465_y0);
  and_gate and_gate_h_u_cla24_and466_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and466_y0);
  and_gate and_gate_h_u_cla24_and467_y0(h_u_cla24_and466_y0, h_u_cla24_and465_y0, h_u_cla24_and467_y0);
  and_gate and_gate_h_u_cla24_and468_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and468_y0);
  and_gate and_gate_h_u_cla24_and469_y0(h_u_cla24_and468_y0, h_u_cla24_and467_y0, h_u_cla24_and469_y0);
  and_gate and_gate_h_u_cla24_and470_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and470_y0);
  and_gate and_gate_h_u_cla24_and471_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and471_y0);
  and_gate and_gate_h_u_cla24_and472_y0(h_u_cla24_and471_y0, h_u_cla24_and470_y0, h_u_cla24_and472_y0);
  and_gate and_gate_h_u_cla24_and473_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and473_y0);
  and_gate and_gate_h_u_cla24_and474_y0(h_u_cla24_and473_y0, h_u_cla24_and472_y0, h_u_cla24_and474_y0);
  and_gate and_gate_h_u_cla24_and475_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and475_y0);
  and_gate and_gate_h_u_cla24_and476_y0(h_u_cla24_and475_y0, h_u_cla24_and474_y0, h_u_cla24_and476_y0);
  and_gate and_gate_h_u_cla24_and477_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and477_y0);
  and_gate and_gate_h_u_cla24_and478_y0(h_u_cla24_and477_y0, h_u_cla24_and476_y0, h_u_cla24_and478_y0);
  and_gate and_gate_h_u_cla24_and479_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and479_y0);
  and_gate and_gate_h_u_cla24_and480_y0(h_u_cla24_and479_y0, h_u_cla24_and478_y0, h_u_cla24_and480_y0);
  and_gate and_gate_h_u_cla24_and481_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and481_y0);
  and_gate and_gate_h_u_cla24_and482_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and482_y0);
  and_gate and_gate_h_u_cla24_and483_y0(h_u_cla24_and482_y0, h_u_cla24_and481_y0, h_u_cla24_and483_y0);
  and_gate and_gate_h_u_cla24_and484_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and484_y0);
  and_gate and_gate_h_u_cla24_and485_y0(h_u_cla24_and484_y0, h_u_cla24_and483_y0, h_u_cla24_and485_y0);
  and_gate and_gate_h_u_cla24_and486_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and486_y0);
  and_gate and_gate_h_u_cla24_and487_y0(h_u_cla24_and486_y0, h_u_cla24_and485_y0, h_u_cla24_and487_y0);
  and_gate and_gate_h_u_cla24_and488_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and488_y0);
  and_gate and_gate_h_u_cla24_and489_y0(h_u_cla24_and488_y0, h_u_cla24_and487_y0, h_u_cla24_and489_y0);
  and_gate and_gate_h_u_cla24_and490_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and490_y0);
  and_gate and_gate_h_u_cla24_and491_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and491_y0);
  and_gate and_gate_h_u_cla24_and492_y0(h_u_cla24_and491_y0, h_u_cla24_and490_y0, h_u_cla24_and492_y0);
  and_gate and_gate_h_u_cla24_and493_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and493_y0);
  and_gate and_gate_h_u_cla24_and494_y0(h_u_cla24_and493_y0, h_u_cla24_and492_y0, h_u_cla24_and494_y0);
  and_gate and_gate_h_u_cla24_and495_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and495_y0);
  and_gate and_gate_h_u_cla24_and496_y0(h_u_cla24_and495_y0, h_u_cla24_and494_y0, h_u_cla24_and496_y0);
  and_gate and_gate_h_u_cla24_and497_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and497_y0);
  and_gate and_gate_h_u_cla24_and498_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and498_y0);
  and_gate and_gate_h_u_cla24_and499_y0(h_u_cla24_and498_y0, h_u_cla24_and497_y0, h_u_cla24_and499_y0);
  and_gate and_gate_h_u_cla24_and500_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and500_y0);
  and_gate and_gate_h_u_cla24_and501_y0(h_u_cla24_and500_y0, h_u_cla24_and499_y0, h_u_cla24_and501_y0);
  and_gate and_gate_h_u_cla24_and502_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and502_y0);
  and_gate and_gate_h_u_cla24_and503_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and503_y0);
  and_gate and_gate_h_u_cla24_and504_y0(h_u_cla24_and503_y0, h_u_cla24_and502_y0, h_u_cla24_and504_y0);
  and_gate and_gate_h_u_cla24_and505_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and505_y0);
  or_gate or_gate_h_u_cla24_or55_y0(h_u_cla24_and505_y0, h_u_cla24_and405_y0, h_u_cla24_or55_y0);
  or_gate or_gate_h_u_cla24_or56_y0(h_u_cla24_or55_y0, h_u_cla24_and424_y0, h_u_cla24_or56_y0);
  or_gate or_gate_h_u_cla24_or57_y0(h_u_cla24_or56_y0, h_u_cla24_and441_y0, h_u_cla24_or57_y0);
  or_gate or_gate_h_u_cla24_or58_y0(h_u_cla24_or57_y0, h_u_cla24_and456_y0, h_u_cla24_or58_y0);
  or_gate or_gate_h_u_cla24_or59_y0(h_u_cla24_or58_y0, h_u_cla24_and469_y0, h_u_cla24_or59_y0);
  or_gate or_gate_h_u_cla24_or60_y0(h_u_cla24_or59_y0, h_u_cla24_and480_y0, h_u_cla24_or60_y0);
  or_gate or_gate_h_u_cla24_or61_y0(h_u_cla24_or60_y0, h_u_cla24_and489_y0, h_u_cla24_or61_y0);
  or_gate or_gate_h_u_cla24_or62_y0(h_u_cla24_or61_y0, h_u_cla24_and496_y0, h_u_cla24_or62_y0);
  or_gate or_gate_h_u_cla24_or63_y0(h_u_cla24_or62_y0, h_u_cla24_and501_y0, h_u_cla24_or63_y0);
  or_gate or_gate_h_u_cla24_or64_y0(h_u_cla24_or63_y0, h_u_cla24_and504_y0, h_u_cla24_or64_y0);
  or_gate or_gate_h_u_cla24_or65_y0(h_u_cla24_pg_logic10_y1, h_u_cla24_or64_y0, h_u_cla24_or65_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic11_y0(a_11, b_11, h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_pg_logic11_y2);
  xor_gate xor_gate_h_u_cla24_xor11_y0(h_u_cla24_pg_logic11_y2, h_u_cla24_or65_y0, h_u_cla24_xor11_y0);
  and_gate and_gate_h_u_cla24_and506_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and506_y0);
  and_gate and_gate_h_u_cla24_and507_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and507_y0);
  and_gate and_gate_h_u_cla24_and508_y0(h_u_cla24_and507_y0, h_u_cla24_and506_y0, h_u_cla24_and508_y0);
  and_gate and_gate_h_u_cla24_and509_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and509_y0);
  and_gate and_gate_h_u_cla24_and510_y0(h_u_cla24_and509_y0, h_u_cla24_and508_y0, h_u_cla24_and510_y0);
  and_gate and_gate_h_u_cla24_and511_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and511_y0);
  and_gate and_gate_h_u_cla24_and512_y0(h_u_cla24_and511_y0, h_u_cla24_and510_y0, h_u_cla24_and512_y0);
  and_gate and_gate_h_u_cla24_and513_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and513_y0);
  and_gate and_gate_h_u_cla24_and514_y0(h_u_cla24_and513_y0, h_u_cla24_and512_y0, h_u_cla24_and514_y0);
  and_gate and_gate_h_u_cla24_and515_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and515_y0);
  and_gate and_gate_h_u_cla24_and516_y0(h_u_cla24_and515_y0, h_u_cla24_and514_y0, h_u_cla24_and516_y0);
  and_gate and_gate_h_u_cla24_and517_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and517_y0);
  and_gate and_gate_h_u_cla24_and518_y0(h_u_cla24_and517_y0, h_u_cla24_and516_y0, h_u_cla24_and518_y0);
  and_gate and_gate_h_u_cla24_and519_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and519_y0);
  and_gate and_gate_h_u_cla24_and520_y0(h_u_cla24_and519_y0, h_u_cla24_and518_y0, h_u_cla24_and520_y0);
  and_gate and_gate_h_u_cla24_and521_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and521_y0);
  and_gate and_gate_h_u_cla24_and522_y0(h_u_cla24_and521_y0, h_u_cla24_and520_y0, h_u_cla24_and522_y0);
  and_gate and_gate_h_u_cla24_and523_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and523_y0);
  and_gate and_gate_h_u_cla24_and524_y0(h_u_cla24_and523_y0, h_u_cla24_and522_y0, h_u_cla24_and524_y0);
  and_gate and_gate_h_u_cla24_and525_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and525_y0);
  and_gate and_gate_h_u_cla24_and526_y0(h_u_cla24_and525_y0, h_u_cla24_and524_y0, h_u_cla24_and526_y0);
  and_gate and_gate_h_u_cla24_and527_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and527_y0);
  and_gate and_gate_h_u_cla24_and528_y0(h_u_cla24_and527_y0, h_u_cla24_and526_y0, h_u_cla24_and528_y0);
  and_gate and_gate_h_u_cla24_and529_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and529_y0);
  and_gate and_gate_h_u_cla24_and530_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and530_y0);
  and_gate and_gate_h_u_cla24_and531_y0(h_u_cla24_and530_y0, h_u_cla24_and529_y0, h_u_cla24_and531_y0);
  and_gate and_gate_h_u_cla24_and532_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and532_y0);
  and_gate and_gate_h_u_cla24_and533_y0(h_u_cla24_and532_y0, h_u_cla24_and531_y0, h_u_cla24_and533_y0);
  and_gate and_gate_h_u_cla24_and534_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and534_y0);
  and_gate and_gate_h_u_cla24_and535_y0(h_u_cla24_and534_y0, h_u_cla24_and533_y0, h_u_cla24_and535_y0);
  and_gate and_gate_h_u_cla24_and536_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and536_y0);
  and_gate and_gate_h_u_cla24_and537_y0(h_u_cla24_and536_y0, h_u_cla24_and535_y0, h_u_cla24_and537_y0);
  and_gate and_gate_h_u_cla24_and538_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and538_y0);
  and_gate and_gate_h_u_cla24_and539_y0(h_u_cla24_and538_y0, h_u_cla24_and537_y0, h_u_cla24_and539_y0);
  and_gate and_gate_h_u_cla24_and540_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and540_y0);
  and_gate and_gate_h_u_cla24_and541_y0(h_u_cla24_and540_y0, h_u_cla24_and539_y0, h_u_cla24_and541_y0);
  and_gate and_gate_h_u_cla24_and542_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and542_y0);
  and_gate and_gate_h_u_cla24_and543_y0(h_u_cla24_and542_y0, h_u_cla24_and541_y0, h_u_cla24_and543_y0);
  and_gate and_gate_h_u_cla24_and544_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and544_y0);
  and_gate and_gate_h_u_cla24_and545_y0(h_u_cla24_and544_y0, h_u_cla24_and543_y0, h_u_cla24_and545_y0);
  and_gate and_gate_h_u_cla24_and546_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and546_y0);
  and_gate and_gate_h_u_cla24_and547_y0(h_u_cla24_and546_y0, h_u_cla24_and545_y0, h_u_cla24_and547_y0);
  and_gate and_gate_h_u_cla24_and548_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and548_y0);
  and_gate and_gate_h_u_cla24_and549_y0(h_u_cla24_and548_y0, h_u_cla24_and547_y0, h_u_cla24_and549_y0);
  and_gate and_gate_h_u_cla24_and550_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and550_y0);
  and_gate and_gate_h_u_cla24_and551_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and551_y0);
  and_gate and_gate_h_u_cla24_and552_y0(h_u_cla24_and551_y0, h_u_cla24_and550_y0, h_u_cla24_and552_y0);
  and_gate and_gate_h_u_cla24_and553_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and553_y0);
  and_gate and_gate_h_u_cla24_and554_y0(h_u_cla24_and553_y0, h_u_cla24_and552_y0, h_u_cla24_and554_y0);
  and_gate and_gate_h_u_cla24_and555_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and555_y0);
  and_gate and_gate_h_u_cla24_and556_y0(h_u_cla24_and555_y0, h_u_cla24_and554_y0, h_u_cla24_and556_y0);
  and_gate and_gate_h_u_cla24_and557_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and557_y0);
  and_gate and_gate_h_u_cla24_and558_y0(h_u_cla24_and557_y0, h_u_cla24_and556_y0, h_u_cla24_and558_y0);
  and_gate and_gate_h_u_cla24_and559_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and559_y0);
  and_gate and_gate_h_u_cla24_and560_y0(h_u_cla24_and559_y0, h_u_cla24_and558_y0, h_u_cla24_and560_y0);
  and_gate and_gate_h_u_cla24_and561_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and561_y0);
  and_gate and_gate_h_u_cla24_and562_y0(h_u_cla24_and561_y0, h_u_cla24_and560_y0, h_u_cla24_and562_y0);
  and_gate and_gate_h_u_cla24_and563_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and563_y0);
  and_gate and_gate_h_u_cla24_and564_y0(h_u_cla24_and563_y0, h_u_cla24_and562_y0, h_u_cla24_and564_y0);
  and_gate and_gate_h_u_cla24_and565_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and565_y0);
  and_gate and_gate_h_u_cla24_and566_y0(h_u_cla24_and565_y0, h_u_cla24_and564_y0, h_u_cla24_and566_y0);
  and_gate and_gate_h_u_cla24_and567_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and567_y0);
  and_gate and_gate_h_u_cla24_and568_y0(h_u_cla24_and567_y0, h_u_cla24_and566_y0, h_u_cla24_and568_y0);
  and_gate and_gate_h_u_cla24_and569_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and569_y0);
  and_gate and_gate_h_u_cla24_and570_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and570_y0);
  and_gate and_gate_h_u_cla24_and571_y0(h_u_cla24_and570_y0, h_u_cla24_and569_y0, h_u_cla24_and571_y0);
  and_gate and_gate_h_u_cla24_and572_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and572_y0);
  and_gate and_gate_h_u_cla24_and573_y0(h_u_cla24_and572_y0, h_u_cla24_and571_y0, h_u_cla24_and573_y0);
  and_gate and_gate_h_u_cla24_and574_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and574_y0);
  and_gate and_gate_h_u_cla24_and575_y0(h_u_cla24_and574_y0, h_u_cla24_and573_y0, h_u_cla24_and575_y0);
  and_gate and_gate_h_u_cla24_and576_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and576_y0);
  and_gate and_gate_h_u_cla24_and577_y0(h_u_cla24_and576_y0, h_u_cla24_and575_y0, h_u_cla24_and577_y0);
  and_gate and_gate_h_u_cla24_and578_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and578_y0);
  and_gate and_gate_h_u_cla24_and579_y0(h_u_cla24_and578_y0, h_u_cla24_and577_y0, h_u_cla24_and579_y0);
  and_gate and_gate_h_u_cla24_and580_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and580_y0);
  and_gate and_gate_h_u_cla24_and581_y0(h_u_cla24_and580_y0, h_u_cla24_and579_y0, h_u_cla24_and581_y0);
  and_gate and_gate_h_u_cla24_and582_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and582_y0);
  and_gate and_gate_h_u_cla24_and583_y0(h_u_cla24_and582_y0, h_u_cla24_and581_y0, h_u_cla24_and583_y0);
  and_gate and_gate_h_u_cla24_and584_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and584_y0);
  and_gate and_gate_h_u_cla24_and585_y0(h_u_cla24_and584_y0, h_u_cla24_and583_y0, h_u_cla24_and585_y0);
  and_gate and_gate_h_u_cla24_and586_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and586_y0);
  and_gate and_gate_h_u_cla24_and587_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and587_y0);
  and_gate and_gate_h_u_cla24_and588_y0(h_u_cla24_and587_y0, h_u_cla24_and586_y0, h_u_cla24_and588_y0);
  and_gate and_gate_h_u_cla24_and589_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and589_y0);
  and_gate and_gate_h_u_cla24_and590_y0(h_u_cla24_and589_y0, h_u_cla24_and588_y0, h_u_cla24_and590_y0);
  and_gate and_gate_h_u_cla24_and591_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and591_y0);
  and_gate and_gate_h_u_cla24_and592_y0(h_u_cla24_and591_y0, h_u_cla24_and590_y0, h_u_cla24_and592_y0);
  and_gate and_gate_h_u_cla24_and593_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and593_y0);
  and_gate and_gate_h_u_cla24_and594_y0(h_u_cla24_and593_y0, h_u_cla24_and592_y0, h_u_cla24_and594_y0);
  and_gate and_gate_h_u_cla24_and595_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and595_y0);
  and_gate and_gate_h_u_cla24_and596_y0(h_u_cla24_and595_y0, h_u_cla24_and594_y0, h_u_cla24_and596_y0);
  and_gate and_gate_h_u_cla24_and597_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and597_y0);
  and_gate and_gate_h_u_cla24_and598_y0(h_u_cla24_and597_y0, h_u_cla24_and596_y0, h_u_cla24_and598_y0);
  and_gate and_gate_h_u_cla24_and599_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and599_y0);
  and_gate and_gate_h_u_cla24_and600_y0(h_u_cla24_and599_y0, h_u_cla24_and598_y0, h_u_cla24_and600_y0);
  and_gate and_gate_h_u_cla24_and601_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and601_y0);
  and_gate and_gate_h_u_cla24_and602_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and602_y0);
  and_gate and_gate_h_u_cla24_and603_y0(h_u_cla24_and602_y0, h_u_cla24_and601_y0, h_u_cla24_and603_y0);
  and_gate and_gate_h_u_cla24_and604_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and604_y0);
  and_gate and_gate_h_u_cla24_and605_y0(h_u_cla24_and604_y0, h_u_cla24_and603_y0, h_u_cla24_and605_y0);
  and_gate and_gate_h_u_cla24_and606_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and606_y0);
  and_gate and_gate_h_u_cla24_and607_y0(h_u_cla24_and606_y0, h_u_cla24_and605_y0, h_u_cla24_and607_y0);
  and_gate and_gate_h_u_cla24_and608_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and608_y0);
  and_gate and_gate_h_u_cla24_and609_y0(h_u_cla24_and608_y0, h_u_cla24_and607_y0, h_u_cla24_and609_y0);
  and_gate and_gate_h_u_cla24_and610_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and610_y0);
  and_gate and_gate_h_u_cla24_and611_y0(h_u_cla24_and610_y0, h_u_cla24_and609_y0, h_u_cla24_and611_y0);
  and_gate and_gate_h_u_cla24_and612_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and612_y0);
  and_gate and_gate_h_u_cla24_and613_y0(h_u_cla24_and612_y0, h_u_cla24_and611_y0, h_u_cla24_and613_y0);
  and_gate and_gate_h_u_cla24_and614_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and614_y0);
  and_gate and_gate_h_u_cla24_and615_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and615_y0);
  and_gate and_gate_h_u_cla24_and616_y0(h_u_cla24_and615_y0, h_u_cla24_and614_y0, h_u_cla24_and616_y0);
  and_gate and_gate_h_u_cla24_and617_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and617_y0);
  and_gate and_gate_h_u_cla24_and618_y0(h_u_cla24_and617_y0, h_u_cla24_and616_y0, h_u_cla24_and618_y0);
  and_gate and_gate_h_u_cla24_and619_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and619_y0);
  and_gate and_gate_h_u_cla24_and620_y0(h_u_cla24_and619_y0, h_u_cla24_and618_y0, h_u_cla24_and620_y0);
  and_gate and_gate_h_u_cla24_and621_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and621_y0);
  and_gate and_gate_h_u_cla24_and622_y0(h_u_cla24_and621_y0, h_u_cla24_and620_y0, h_u_cla24_and622_y0);
  and_gate and_gate_h_u_cla24_and623_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and623_y0);
  and_gate and_gate_h_u_cla24_and624_y0(h_u_cla24_and623_y0, h_u_cla24_and622_y0, h_u_cla24_and624_y0);
  and_gate and_gate_h_u_cla24_and625_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and625_y0);
  and_gate and_gate_h_u_cla24_and626_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and626_y0);
  and_gate and_gate_h_u_cla24_and627_y0(h_u_cla24_and626_y0, h_u_cla24_and625_y0, h_u_cla24_and627_y0);
  and_gate and_gate_h_u_cla24_and628_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and628_y0);
  and_gate and_gate_h_u_cla24_and629_y0(h_u_cla24_and628_y0, h_u_cla24_and627_y0, h_u_cla24_and629_y0);
  and_gate and_gate_h_u_cla24_and630_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and630_y0);
  and_gate and_gate_h_u_cla24_and631_y0(h_u_cla24_and630_y0, h_u_cla24_and629_y0, h_u_cla24_and631_y0);
  and_gate and_gate_h_u_cla24_and632_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and632_y0);
  and_gate and_gate_h_u_cla24_and633_y0(h_u_cla24_and632_y0, h_u_cla24_and631_y0, h_u_cla24_and633_y0);
  and_gate and_gate_h_u_cla24_and634_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and634_y0);
  and_gate and_gate_h_u_cla24_and635_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and635_y0);
  and_gate and_gate_h_u_cla24_and636_y0(h_u_cla24_and635_y0, h_u_cla24_and634_y0, h_u_cla24_and636_y0);
  and_gate and_gate_h_u_cla24_and637_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and637_y0);
  and_gate and_gate_h_u_cla24_and638_y0(h_u_cla24_and637_y0, h_u_cla24_and636_y0, h_u_cla24_and638_y0);
  and_gate and_gate_h_u_cla24_and639_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and639_y0);
  and_gate and_gate_h_u_cla24_and640_y0(h_u_cla24_and639_y0, h_u_cla24_and638_y0, h_u_cla24_and640_y0);
  and_gate and_gate_h_u_cla24_and641_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and641_y0);
  and_gate and_gate_h_u_cla24_and642_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and642_y0);
  and_gate and_gate_h_u_cla24_and643_y0(h_u_cla24_and642_y0, h_u_cla24_and641_y0, h_u_cla24_and643_y0);
  and_gate and_gate_h_u_cla24_and644_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and644_y0);
  and_gate and_gate_h_u_cla24_and645_y0(h_u_cla24_and644_y0, h_u_cla24_and643_y0, h_u_cla24_and645_y0);
  and_gate and_gate_h_u_cla24_and646_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and646_y0);
  and_gate and_gate_h_u_cla24_and647_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and647_y0);
  and_gate and_gate_h_u_cla24_and648_y0(h_u_cla24_and647_y0, h_u_cla24_and646_y0, h_u_cla24_and648_y0);
  and_gate and_gate_h_u_cla24_and649_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and649_y0);
  or_gate or_gate_h_u_cla24_or66_y0(h_u_cla24_and649_y0, h_u_cla24_and528_y0, h_u_cla24_or66_y0);
  or_gate or_gate_h_u_cla24_or67_y0(h_u_cla24_or66_y0, h_u_cla24_and549_y0, h_u_cla24_or67_y0);
  or_gate or_gate_h_u_cla24_or68_y0(h_u_cla24_or67_y0, h_u_cla24_and568_y0, h_u_cla24_or68_y0);
  or_gate or_gate_h_u_cla24_or69_y0(h_u_cla24_or68_y0, h_u_cla24_and585_y0, h_u_cla24_or69_y0);
  or_gate or_gate_h_u_cla24_or70_y0(h_u_cla24_or69_y0, h_u_cla24_and600_y0, h_u_cla24_or70_y0);
  or_gate or_gate_h_u_cla24_or71_y0(h_u_cla24_or70_y0, h_u_cla24_and613_y0, h_u_cla24_or71_y0);
  or_gate or_gate_h_u_cla24_or72_y0(h_u_cla24_or71_y0, h_u_cla24_and624_y0, h_u_cla24_or72_y0);
  or_gate or_gate_h_u_cla24_or73_y0(h_u_cla24_or72_y0, h_u_cla24_and633_y0, h_u_cla24_or73_y0);
  or_gate or_gate_h_u_cla24_or74_y0(h_u_cla24_or73_y0, h_u_cla24_and640_y0, h_u_cla24_or74_y0);
  or_gate or_gate_h_u_cla24_or75_y0(h_u_cla24_or74_y0, h_u_cla24_and645_y0, h_u_cla24_or75_y0);
  or_gate or_gate_h_u_cla24_or76_y0(h_u_cla24_or75_y0, h_u_cla24_and648_y0, h_u_cla24_or76_y0);
  or_gate or_gate_h_u_cla24_or77_y0(h_u_cla24_pg_logic11_y1, h_u_cla24_or76_y0, h_u_cla24_or77_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic12_y0(a_12, b_12, h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_pg_logic12_y2);
  xor_gate xor_gate_h_u_cla24_xor12_y0(h_u_cla24_pg_logic12_y2, h_u_cla24_or77_y0, h_u_cla24_xor12_y0);
  and_gate and_gate_h_u_cla24_and650_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and650_y0);
  and_gate and_gate_h_u_cla24_and651_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and651_y0);
  and_gate and_gate_h_u_cla24_and652_y0(h_u_cla24_and651_y0, h_u_cla24_and650_y0, h_u_cla24_and652_y0);
  and_gate and_gate_h_u_cla24_and653_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and653_y0);
  and_gate and_gate_h_u_cla24_and654_y0(h_u_cla24_and653_y0, h_u_cla24_and652_y0, h_u_cla24_and654_y0);
  and_gate and_gate_h_u_cla24_and655_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and655_y0);
  and_gate and_gate_h_u_cla24_and656_y0(h_u_cla24_and655_y0, h_u_cla24_and654_y0, h_u_cla24_and656_y0);
  and_gate and_gate_h_u_cla24_and657_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and657_y0);
  and_gate and_gate_h_u_cla24_and658_y0(h_u_cla24_and657_y0, h_u_cla24_and656_y0, h_u_cla24_and658_y0);
  and_gate and_gate_h_u_cla24_and659_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and659_y0);
  and_gate and_gate_h_u_cla24_and660_y0(h_u_cla24_and659_y0, h_u_cla24_and658_y0, h_u_cla24_and660_y0);
  and_gate and_gate_h_u_cla24_and661_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and661_y0);
  and_gate and_gate_h_u_cla24_and662_y0(h_u_cla24_and661_y0, h_u_cla24_and660_y0, h_u_cla24_and662_y0);
  and_gate and_gate_h_u_cla24_and663_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and663_y0);
  and_gate and_gate_h_u_cla24_and664_y0(h_u_cla24_and663_y0, h_u_cla24_and662_y0, h_u_cla24_and664_y0);
  and_gate and_gate_h_u_cla24_and665_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and665_y0);
  and_gate and_gate_h_u_cla24_and666_y0(h_u_cla24_and665_y0, h_u_cla24_and664_y0, h_u_cla24_and666_y0);
  and_gate and_gate_h_u_cla24_and667_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and667_y0);
  and_gate and_gate_h_u_cla24_and668_y0(h_u_cla24_and667_y0, h_u_cla24_and666_y0, h_u_cla24_and668_y0);
  and_gate and_gate_h_u_cla24_and669_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and669_y0);
  and_gate and_gate_h_u_cla24_and670_y0(h_u_cla24_and669_y0, h_u_cla24_and668_y0, h_u_cla24_and670_y0);
  and_gate and_gate_h_u_cla24_and671_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and671_y0);
  and_gate and_gate_h_u_cla24_and672_y0(h_u_cla24_and671_y0, h_u_cla24_and670_y0, h_u_cla24_and672_y0);
  and_gate and_gate_h_u_cla24_and673_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and673_y0);
  and_gate and_gate_h_u_cla24_and674_y0(h_u_cla24_and673_y0, h_u_cla24_and672_y0, h_u_cla24_and674_y0);
  and_gate and_gate_h_u_cla24_and675_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and675_y0);
  and_gate and_gate_h_u_cla24_and676_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and676_y0);
  and_gate and_gate_h_u_cla24_and677_y0(h_u_cla24_and676_y0, h_u_cla24_and675_y0, h_u_cla24_and677_y0);
  and_gate and_gate_h_u_cla24_and678_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and678_y0);
  and_gate and_gate_h_u_cla24_and679_y0(h_u_cla24_and678_y0, h_u_cla24_and677_y0, h_u_cla24_and679_y0);
  and_gate and_gate_h_u_cla24_and680_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and680_y0);
  and_gate and_gate_h_u_cla24_and681_y0(h_u_cla24_and680_y0, h_u_cla24_and679_y0, h_u_cla24_and681_y0);
  and_gate and_gate_h_u_cla24_and682_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and682_y0);
  and_gate and_gate_h_u_cla24_and683_y0(h_u_cla24_and682_y0, h_u_cla24_and681_y0, h_u_cla24_and683_y0);
  and_gate and_gate_h_u_cla24_and684_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and684_y0);
  and_gate and_gate_h_u_cla24_and685_y0(h_u_cla24_and684_y0, h_u_cla24_and683_y0, h_u_cla24_and685_y0);
  and_gate and_gate_h_u_cla24_and686_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and686_y0);
  and_gate and_gate_h_u_cla24_and687_y0(h_u_cla24_and686_y0, h_u_cla24_and685_y0, h_u_cla24_and687_y0);
  and_gate and_gate_h_u_cla24_and688_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and688_y0);
  and_gate and_gate_h_u_cla24_and689_y0(h_u_cla24_and688_y0, h_u_cla24_and687_y0, h_u_cla24_and689_y0);
  and_gate and_gate_h_u_cla24_and690_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and690_y0);
  and_gate and_gate_h_u_cla24_and691_y0(h_u_cla24_and690_y0, h_u_cla24_and689_y0, h_u_cla24_and691_y0);
  and_gate and_gate_h_u_cla24_and692_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and692_y0);
  and_gate and_gate_h_u_cla24_and693_y0(h_u_cla24_and692_y0, h_u_cla24_and691_y0, h_u_cla24_and693_y0);
  and_gate and_gate_h_u_cla24_and694_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and694_y0);
  and_gate and_gate_h_u_cla24_and695_y0(h_u_cla24_and694_y0, h_u_cla24_and693_y0, h_u_cla24_and695_y0);
  and_gate and_gate_h_u_cla24_and696_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and696_y0);
  and_gate and_gate_h_u_cla24_and697_y0(h_u_cla24_and696_y0, h_u_cla24_and695_y0, h_u_cla24_and697_y0);
  and_gate and_gate_h_u_cla24_and698_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and698_y0);
  and_gate and_gate_h_u_cla24_and699_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and699_y0);
  and_gate and_gate_h_u_cla24_and700_y0(h_u_cla24_and699_y0, h_u_cla24_and698_y0, h_u_cla24_and700_y0);
  and_gate and_gate_h_u_cla24_and701_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and701_y0);
  and_gate and_gate_h_u_cla24_and702_y0(h_u_cla24_and701_y0, h_u_cla24_and700_y0, h_u_cla24_and702_y0);
  and_gate and_gate_h_u_cla24_and703_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and703_y0);
  and_gate and_gate_h_u_cla24_and704_y0(h_u_cla24_and703_y0, h_u_cla24_and702_y0, h_u_cla24_and704_y0);
  and_gate and_gate_h_u_cla24_and705_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and705_y0);
  and_gate and_gate_h_u_cla24_and706_y0(h_u_cla24_and705_y0, h_u_cla24_and704_y0, h_u_cla24_and706_y0);
  and_gate and_gate_h_u_cla24_and707_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and707_y0);
  and_gate and_gate_h_u_cla24_and708_y0(h_u_cla24_and707_y0, h_u_cla24_and706_y0, h_u_cla24_and708_y0);
  and_gate and_gate_h_u_cla24_and709_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and709_y0);
  and_gate and_gate_h_u_cla24_and710_y0(h_u_cla24_and709_y0, h_u_cla24_and708_y0, h_u_cla24_and710_y0);
  and_gate and_gate_h_u_cla24_and711_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and711_y0);
  and_gate and_gate_h_u_cla24_and712_y0(h_u_cla24_and711_y0, h_u_cla24_and710_y0, h_u_cla24_and712_y0);
  and_gate and_gate_h_u_cla24_and713_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and713_y0);
  and_gate and_gate_h_u_cla24_and714_y0(h_u_cla24_and713_y0, h_u_cla24_and712_y0, h_u_cla24_and714_y0);
  and_gate and_gate_h_u_cla24_and715_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and715_y0);
  and_gate and_gate_h_u_cla24_and716_y0(h_u_cla24_and715_y0, h_u_cla24_and714_y0, h_u_cla24_and716_y0);
  and_gate and_gate_h_u_cla24_and717_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and717_y0);
  and_gate and_gate_h_u_cla24_and718_y0(h_u_cla24_and717_y0, h_u_cla24_and716_y0, h_u_cla24_and718_y0);
  and_gate and_gate_h_u_cla24_and719_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and719_y0);
  and_gate and_gate_h_u_cla24_and720_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and720_y0);
  and_gate and_gate_h_u_cla24_and721_y0(h_u_cla24_and720_y0, h_u_cla24_and719_y0, h_u_cla24_and721_y0);
  and_gate and_gate_h_u_cla24_and722_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and722_y0);
  and_gate and_gate_h_u_cla24_and723_y0(h_u_cla24_and722_y0, h_u_cla24_and721_y0, h_u_cla24_and723_y0);
  and_gate and_gate_h_u_cla24_and724_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and724_y0);
  and_gate and_gate_h_u_cla24_and725_y0(h_u_cla24_and724_y0, h_u_cla24_and723_y0, h_u_cla24_and725_y0);
  and_gate and_gate_h_u_cla24_and726_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and726_y0);
  and_gate and_gate_h_u_cla24_and727_y0(h_u_cla24_and726_y0, h_u_cla24_and725_y0, h_u_cla24_and727_y0);
  and_gate and_gate_h_u_cla24_and728_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and728_y0);
  and_gate and_gate_h_u_cla24_and729_y0(h_u_cla24_and728_y0, h_u_cla24_and727_y0, h_u_cla24_and729_y0);
  and_gate and_gate_h_u_cla24_and730_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and730_y0);
  and_gate and_gate_h_u_cla24_and731_y0(h_u_cla24_and730_y0, h_u_cla24_and729_y0, h_u_cla24_and731_y0);
  and_gate and_gate_h_u_cla24_and732_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and732_y0);
  and_gate and_gate_h_u_cla24_and733_y0(h_u_cla24_and732_y0, h_u_cla24_and731_y0, h_u_cla24_and733_y0);
  and_gate and_gate_h_u_cla24_and734_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and734_y0);
  and_gate and_gate_h_u_cla24_and735_y0(h_u_cla24_and734_y0, h_u_cla24_and733_y0, h_u_cla24_and735_y0);
  and_gate and_gate_h_u_cla24_and736_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and736_y0);
  and_gate and_gate_h_u_cla24_and737_y0(h_u_cla24_and736_y0, h_u_cla24_and735_y0, h_u_cla24_and737_y0);
  and_gate and_gate_h_u_cla24_and738_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and738_y0);
  and_gate and_gate_h_u_cla24_and739_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and739_y0);
  and_gate and_gate_h_u_cla24_and740_y0(h_u_cla24_and739_y0, h_u_cla24_and738_y0, h_u_cla24_and740_y0);
  and_gate and_gate_h_u_cla24_and741_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and741_y0);
  and_gate and_gate_h_u_cla24_and742_y0(h_u_cla24_and741_y0, h_u_cla24_and740_y0, h_u_cla24_and742_y0);
  and_gate and_gate_h_u_cla24_and743_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and743_y0);
  and_gate and_gate_h_u_cla24_and744_y0(h_u_cla24_and743_y0, h_u_cla24_and742_y0, h_u_cla24_and744_y0);
  and_gate and_gate_h_u_cla24_and745_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and745_y0);
  and_gate and_gate_h_u_cla24_and746_y0(h_u_cla24_and745_y0, h_u_cla24_and744_y0, h_u_cla24_and746_y0);
  and_gate and_gate_h_u_cla24_and747_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and747_y0);
  and_gate and_gate_h_u_cla24_and748_y0(h_u_cla24_and747_y0, h_u_cla24_and746_y0, h_u_cla24_and748_y0);
  and_gate and_gate_h_u_cla24_and749_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and749_y0);
  and_gate and_gate_h_u_cla24_and750_y0(h_u_cla24_and749_y0, h_u_cla24_and748_y0, h_u_cla24_and750_y0);
  and_gate and_gate_h_u_cla24_and751_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and751_y0);
  and_gate and_gate_h_u_cla24_and752_y0(h_u_cla24_and751_y0, h_u_cla24_and750_y0, h_u_cla24_and752_y0);
  and_gate and_gate_h_u_cla24_and753_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and753_y0);
  and_gate and_gate_h_u_cla24_and754_y0(h_u_cla24_and753_y0, h_u_cla24_and752_y0, h_u_cla24_and754_y0);
  and_gate and_gate_h_u_cla24_and755_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and755_y0);
  and_gate and_gate_h_u_cla24_and756_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and756_y0);
  and_gate and_gate_h_u_cla24_and757_y0(h_u_cla24_and756_y0, h_u_cla24_and755_y0, h_u_cla24_and757_y0);
  and_gate and_gate_h_u_cla24_and758_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and758_y0);
  and_gate and_gate_h_u_cla24_and759_y0(h_u_cla24_and758_y0, h_u_cla24_and757_y0, h_u_cla24_and759_y0);
  and_gate and_gate_h_u_cla24_and760_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and760_y0);
  and_gate and_gate_h_u_cla24_and761_y0(h_u_cla24_and760_y0, h_u_cla24_and759_y0, h_u_cla24_and761_y0);
  and_gate and_gate_h_u_cla24_and762_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and762_y0);
  and_gate and_gate_h_u_cla24_and763_y0(h_u_cla24_and762_y0, h_u_cla24_and761_y0, h_u_cla24_and763_y0);
  and_gate and_gate_h_u_cla24_and764_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and764_y0);
  and_gate and_gate_h_u_cla24_and765_y0(h_u_cla24_and764_y0, h_u_cla24_and763_y0, h_u_cla24_and765_y0);
  and_gate and_gate_h_u_cla24_and766_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and766_y0);
  and_gate and_gate_h_u_cla24_and767_y0(h_u_cla24_and766_y0, h_u_cla24_and765_y0, h_u_cla24_and767_y0);
  and_gate and_gate_h_u_cla24_and768_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and768_y0);
  and_gate and_gate_h_u_cla24_and769_y0(h_u_cla24_and768_y0, h_u_cla24_and767_y0, h_u_cla24_and769_y0);
  and_gate and_gate_h_u_cla24_and770_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and770_y0);
  and_gate and_gate_h_u_cla24_and771_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and771_y0);
  and_gate and_gate_h_u_cla24_and772_y0(h_u_cla24_and771_y0, h_u_cla24_and770_y0, h_u_cla24_and772_y0);
  and_gate and_gate_h_u_cla24_and773_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and773_y0);
  and_gate and_gate_h_u_cla24_and774_y0(h_u_cla24_and773_y0, h_u_cla24_and772_y0, h_u_cla24_and774_y0);
  and_gate and_gate_h_u_cla24_and775_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and775_y0);
  and_gate and_gate_h_u_cla24_and776_y0(h_u_cla24_and775_y0, h_u_cla24_and774_y0, h_u_cla24_and776_y0);
  and_gate and_gate_h_u_cla24_and777_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and777_y0);
  and_gate and_gate_h_u_cla24_and778_y0(h_u_cla24_and777_y0, h_u_cla24_and776_y0, h_u_cla24_and778_y0);
  and_gate and_gate_h_u_cla24_and779_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and779_y0);
  and_gate and_gate_h_u_cla24_and780_y0(h_u_cla24_and779_y0, h_u_cla24_and778_y0, h_u_cla24_and780_y0);
  and_gate and_gate_h_u_cla24_and781_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and781_y0);
  and_gate and_gate_h_u_cla24_and782_y0(h_u_cla24_and781_y0, h_u_cla24_and780_y0, h_u_cla24_and782_y0);
  and_gate and_gate_h_u_cla24_and783_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and783_y0);
  and_gate and_gate_h_u_cla24_and784_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and784_y0);
  and_gate and_gate_h_u_cla24_and785_y0(h_u_cla24_and784_y0, h_u_cla24_and783_y0, h_u_cla24_and785_y0);
  and_gate and_gate_h_u_cla24_and786_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and786_y0);
  and_gate and_gate_h_u_cla24_and787_y0(h_u_cla24_and786_y0, h_u_cla24_and785_y0, h_u_cla24_and787_y0);
  and_gate and_gate_h_u_cla24_and788_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and788_y0);
  and_gate and_gate_h_u_cla24_and789_y0(h_u_cla24_and788_y0, h_u_cla24_and787_y0, h_u_cla24_and789_y0);
  and_gate and_gate_h_u_cla24_and790_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and790_y0);
  and_gate and_gate_h_u_cla24_and791_y0(h_u_cla24_and790_y0, h_u_cla24_and789_y0, h_u_cla24_and791_y0);
  and_gate and_gate_h_u_cla24_and792_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and792_y0);
  and_gate and_gate_h_u_cla24_and793_y0(h_u_cla24_and792_y0, h_u_cla24_and791_y0, h_u_cla24_and793_y0);
  and_gate and_gate_h_u_cla24_and794_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and794_y0);
  and_gate and_gate_h_u_cla24_and795_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and795_y0);
  and_gate and_gate_h_u_cla24_and796_y0(h_u_cla24_and795_y0, h_u_cla24_and794_y0, h_u_cla24_and796_y0);
  and_gate and_gate_h_u_cla24_and797_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and797_y0);
  and_gate and_gate_h_u_cla24_and798_y0(h_u_cla24_and797_y0, h_u_cla24_and796_y0, h_u_cla24_and798_y0);
  and_gate and_gate_h_u_cla24_and799_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and799_y0);
  and_gate and_gate_h_u_cla24_and800_y0(h_u_cla24_and799_y0, h_u_cla24_and798_y0, h_u_cla24_and800_y0);
  and_gate and_gate_h_u_cla24_and801_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and801_y0);
  and_gate and_gate_h_u_cla24_and802_y0(h_u_cla24_and801_y0, h_u_cla24_and800_y0, h_u_cla24_and802_y0);
  and_gate and_gate_h_u_cla24_and803_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and803_y0);
  and_gate and_gate_h_u_cla24_and804_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and804_y0);
  and_gate and_gate_h_u_cla24_and805_y0(h_u_cla24_and804_y0, h_u_cla24_and803_y0, h_u_cla24_and805_y0);
  and_gate and_gate_h_u_cla24_and806_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and806_y0);
  and_gate and_gate_h_u_cla24_and807_y0(h_u_cla24_and806_y0, h_u_cla24_and805_y0, h_u_cla24_and807_y0);
  and_gate and_gate_h_u_cla24_and808_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and808_y0);
  and_gate and_gate_h_u_cla24_and809_y0(h_u_cla24_and808_y0, h_u_cla24_and807_y0, h_u_cla24_and809_y0);
  and_gate and_gate_h_u_cla24_and810_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and810_y0);
  and_gate and_gate_h_u_cla24_and811_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and811_y0);
  and_gate and_gate_h_u_cla24_and812_y0(h_u_cla24_and811_y0, h_u_cla24_and810_y0, h_u_cla24_and812_y0);
  and_gate and_gate_h_u_cla24_and813_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and813_y0);
  and_gate and_gate_h_u_cla24_and814_y0(h_u_cla24_and813_y0, h_u_cla24_and812_y0, h_u_cla24_and814_y0);
  and_gate and_gate_h_u_cla24_and815_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and815_y0);
  and_gate and_gate_h_u_cla24_and816_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and816_y0);
  and_gate and_gate_h_u_cla24_and817_y0(h_u_cla24_and816_y0, h_u_cla24_and815_y0, h_u_cla24_and817_y0);
  and_gate and_gate_h_u_cla24_and818_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and818_y0);
  or_gate or_gate_h_u_cla24_or78_y0(h_u_cla24_and818_y0, h_u_cla24_and674_y0, h_u_cla24_or78_y0);
  or_gate or_gate_h_u_cla24_or79_y0(h_u_cla24_or78_y0, h_u_cla24_and697_y0, h_u_cla24_or79_y0);
  or_gate or_gate_h_u_cla24_or80_y0(h_u_cla24_or79_y0, h_u_cla24_and718_y0, h_u_cla24_or80_y0);
  or_gate or_gate_h_u_cla24_or81_y0(h_u_cla24_or80_y0, h_u_cla24_and737_y0, h_u_cla24_or81_y0);
  or_gate or_gate_h_u_cla24_or82_y0(h_u_cla24_or81_y0, h_u_cla24_and754_y0, h_u_cla24_or82_y0);
  or_gate or_gate_h_u_cla24_or83_y0(h_u_cla24_or82_y0, h_u_cla24_and769_y0, h_u_cla24_or83_y0);
  or_gate or_gate_h_u_cla24_or84_y0(h_u_cla24_or83_y0, h_u_cla24_and782_y0, h_u_cla24_or84_y0);
  or_gate or_gate_h_u_cla24_or85_y0(h_u_cla24_or84_y0, h_u_cla24_and793_y0, h_u_cla24_or85_y0);
  or_gate or_gate_h_u_cla24_or86_y0(h_u_cla24_or85_y0, h_u_cla24_and802_y0, h_u_cla24_or86_y0);
  or_gate or_gate_h_u_cla24_or87_y0(h_u_cla24_or86_y0, h_u_cla24_and809_y0, h_u_cla24_or87_y0);
  or_gate or_gate_h_u_cla24_or88_y0(h_u_cla24_or87_y0, h_u_cla24_and814_y0, h_u_cla24_or88_y0);
  or_gate or_gate_h_u_cla24_or89_y0(h_u_cla24_or88_y0, h_u_cla24_and817_y0, h_u_cla24_or89_y0);
  or_gate or_gate_h_u_cla24_or90_y0(h_u_cla24_pg_logic12_y1, h_u_cla24_or89_y0, h_u_cla24_or90_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic13_y0(a_13, b_13, h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_pg_logic13_y2);
  xor_gate xor_gate_h_u_cla24_xor13_y0(h_u_cla24_pg_logic13_y2, h_u_cla24_or90_y0, h_u_cla24_xor13_y0);
  and_gate and_gate_h_u_cla24_and819_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and819_y0);
  and_gate and_gate_h_u_cla24_and820_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and820_y0);
  and_gate and_gate_h_u_cla24_and821_y0(h_u_cla24_and820_y0, h_u_cla24_and819_y0, h_u_cla24_and821_y0);
  and_gate and_gate_h_u_cla24_and822_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and822_y0);
  and_gate and_gate_h_u_cla24_and823_y0(h_u_cla24_and822_y0, h_u_cla24_and821_y0, h_u_cla24_and823_y0);
  and_gate and_gate_h_u_cla24_and824_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and824_y0);
  and_gate and_gate_h_u_cla24_and825_y0(h_u_cla24_and824_y0, h_u_cla24_and823_y0, h_u_cla24_and825_y0);
  and_gate and_gate_h_u_cla24_and826_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and826_y0);
  and_gate and_gate_h_u_cla24_and827_y0(h_u_cla24_and826_y0, h_u_cla24_and825_y0, h_u_cla24_and827_y0);
  and_gate and_gate_h_u_cla24_and828_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and828_y0);
  and_gate and_gate_h_u_cla24_and829_y0(h_u_cla24_and828_y0, h_u_cla24_and827_y0, h_u_cla24_and829_y0);
  and_gate and_gate_h_u_cla24_and830_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and830_y0);
  and_gate and_gate_h_u_cla24_and831_y0(h_u_cla24_and830_y0, h_u_cla24_and829_y0, h_u_cla24_and831_y0);
  and_gate and_gate_h_u_cla24_and832_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and832_y0);
  and_gate and_gate_h_u_cla24_and833_y0(h_u_cla24_and832_y0, h_u_cla24_and831_y0, h_u_cla24_and833_y0);
  and_gate and_gate_h_u_cla24_and834_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and834_y0);
  and_gate and_gate_h_u_cla24_and835_y0(h_u_cla24_and834_y0, h_u_cla24_and833_y0, h_u_cla24_and835_y0);
  and_gate and_gate_h_u_cla24_and836_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and836_y0);
  and_gate and_gate_h_u_cla24_and837_y0(h_u_cla24_and836_y0, h_u_cla24_and835_y0, h_u_cla24_and837_y0);
  and_gate and_gate_h_u_cla24_and838_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and838_y0);
  and_gate and_gate_h_u_cla24_and839_y0(h_u_cla24_and838_y0, h_u_cla24_and837_y0, h_u_cla24_and839_y0);
  and_gate and_gate_h_u_cla24_and840_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and840_y0);
  and_gate and_gate_h_u_cla24_and841_y0(h_u_cla24_and840_y0, h_u_cla24_and839_y0, h_u_cla24_and841_y0);
  and_gate and_gate_h_u_cla24_and842_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and842_y0);
  and_gate and_gate_h_u_cla24_and843_y0(h_u_cla24_and842_y0, h_u_cla24_and841_y0, h_u_cla24_and843_y0);
  and_gate and_gate_h_u_cla24_and844_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and844_y0);
  and_gate and_gate_h_u_cla24_and845_y0(h_u_cla24_and844_y0, h_u_cla24_and843_y0, h_u_cla24_and845_y0);
  and_gate and_gate_h_u_cla24_and846_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and846_y0);
  and_gate and_gate_h_u_cla24_and847_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and847_y0);
  and_gate and_gate_h_u_cla24_and848_y0(h_u_cla24_and847_y0, h_u_cla24_and846_y0, h_u_cla24_and848_y0);
  and_gate and_gate_h_u_cla24_and849_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and849_y0);
  and_gate and_gate_h_u_cla24_and850_y0(h_u_cla24_and849_y0, h_u_cla24_and848_y0, h_u_cla24_and850_y0);
  and_gate and_gate_h_u_cla24_and851_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and851_y0);
  and_gate and_gate_h_u_cla24_and852_y0(h_u_cla24_and851_y0, h_u_cla24_and850_y0, h_u_cla24_and852_y0);
  and_gate and_gate_h_u_cla24_and853_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and853_y0);
  and_gate and_gate_h_u_cla24_and854_y0(h_u_cla24_and853_y0, h_u_cla24_and852_y0, h_u_cla24_and854_y0);
  and_gate and_gate_h_u_cla24_and855_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and855_y0);
  and_gate and_gate_h_u_cla24_and856_y0(h_u_cla24_and855_y0, h_u_cla24_and854_y0, h_u_cla24_and856_y0);
  and_gate and_gate_h_u_cla24_and857_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and857_y0);
  and_gate and_gate_h_u_cla24_and858_y0(h_u_cla24_and857_y0, h_u_cla24_and856_y0, h_u_cla24_and858_y0);
  and_gate and_gate_h_u_cla24_and859_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and859_y0);
  and_gate and_gate_h_u_cla24_and860_y0(h_u_cla24_and859_y0, h_u_cla24_and858_y0, h_u_cla24_and860_y0);
  and_gate and_gate_h_u_cla24_and861_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and861_y0);
  and_gate and_gate_h_u_cla24_and862_y0(h_u_cla24_and861_y0, h_u_cla24_and860_y0, h_u_cla24_and862_y0);
  and_gate and_gate_h_u_cla24_and863_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and863_y0);
  and_gate and_gate_h_u_cla24_and864_y0(h_u_cla24_and863_y0, h_u_cla24_and862_y0, h_u_cla24_and864_y0);
  and_gate and_gate_h_u_cla24_and865_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and865_y0);
  and_gate and_gate_h_u_cla24_and866_y0(h_u_cla24_and865_y0, h_u_cla24_and864_y0, h_u_cla24_and866_y0);
  and_gate and_gate_h_u_cla24_and867_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and867_y0);
  and_gate and_gate_h_u_cla24_and868_y0(h_u_cla24_and867_y0, h_u_cla24_and866_y0, h_u_cla24_and868_y0);
  and_gate and_gate_h_u_cla24_and869_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and869_y0);
  and_gate and_gate_h_u_cla24_and870_y0(h_u_cla24_and869_y0, h_u_cla24_and868_y0, h_u_cla24_and870_y0);
  and_gate and_gate_h_u_cla24_and871_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and871_y0);
  and_gate and_gate_h_u_cla24_and872_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and872_y0);
  and_gate and_gate_h_u_cla24_and873_y0(h_u_cla24_and872_y0, h_u_cla24_and871_y0, h_u_cla24_and873_y0);
  and_gate and_gate_h_u_cla24_and874_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and874_y0);
  and_gate and_gate_h_u_cla24_and875_y0(h_u_cla24_and874_y0, h_u_cla24_and873_y0, h_u_cla24_and875_y0);
  and_gate and_gate_h_u_cla24_and876_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and876_y0);
  and_gate and_gate_h_u_cla24_and877_y0(h_u_cla24_and876_y0, h_u_cla24_and875_y0, h_u_cla24_and877_y0);
  and_gate and_gate_h_u_cla24_and878_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and878_y0);
  and_gate and_gate_h_u_cla24_and879_y0(h_u_cla24_and878_y0, h_u_cla24_and877_y0, h_u_cla24_and879_y0);
  and_gate and_gate_h_u_cla24_and880_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and880_y0);
  and_gate and_gate_h_u_cla24_and881_y0(h_u_cla24_and880_y0, h_u_cla24_and879_y0, h_u_cla24_and881_y0);
  and_gate and_gate_h_u_cla24_and882_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and882_y0);
  and_gate and_gate_h_u_cla24_and883_y0(h_u_cla24_and882_y0, h_u_cla24_and881_y0, h_u_cla24_and883_y0);
  and_gate and_gate_h_u_cla24_and884_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and884_y0);
  and_gate and_gate_h_u_cla24_and885_y0(h_u_cla24_and884_y0, h_u_cla24_and883_y0, h_u_cla24_and885_y0);
  and_gate and_gate_h_u_cla24_and886_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and886_y0);
  and_gate and_gate_h_u_cla24_and887_y0(h_u_cla24_and886_y0, h_u_cla24_and885_y0, h_u_cla24_and887_y0);
  and_gate and_gate_h_u_cla24_and888_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and888_y0);
  and_gate and_gate_h_u_cla24_and889_y0(h_u_cla24_and888_y0, h_u_cla24_and887_y0, h_u_cla24_and889_y0);
  and_gate and_gate_h_u_cla24_and890_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and890_y0);
  and_gate and_gate_h_u_cla24_and891_y0(h_u_cla24_and890_y0, h_u_cla24_and889_y0, h_u_cla24_and891_y0);
  and_gate and_gate_h_u_cla24_and892_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and892_y0);
  and_gate and_gate_h_u_cla24_and893_y0(h_u_cla24_and892_y0, h_u_cla24_and891_y0, h_u_cla24_and893_y0);
  and_gate and_gate_h_u_cla24_and894_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and894_y0);
  and_gate and_gate_h_u_cla24_and895_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and895_y0);
  and_gate and_gate_h_u_cla24_and896_y0(h_u_cla24_and895_y0, h_u_cla24_and894_y0, h_u_cla24_and896_y0);
  and_gate and_gate_h_u_cla24_and897_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and897_y0);
  and_gate and_gate_h_u_cla24_and898_y0(h_u_cla24_and897_y0, h_u_cla24_and896_y0, h_u_cla24_and898_y0);
  and_gate and_gate_h_u_cla24_and899_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and899_y0);
  and_gate and_gate_h_u_cla24_and900_y0(h_u_cla24_and899_y0, h_u_cla24_and898_y0, h_u_cla24_and900_y0);
  and_gate and_gate_h_u_cla24_and901_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and901_y0);
  and_gate and_gate_h_u_cla24_and902_y0(h_u_cla24_and901_y0, h_u_cla24_and900_y0, h_u_cla24_and902_y0);
  and_gate and_gate_h_u_cla24_and903_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and903_y0);
  and_gate and_gate_h_u_cla24_and904_y0(h_u_cla24_and903_y0, h_u_cla24_and902_y0, h_u_cla24_and904_y0);
  and_gate and_gate_h_u_cla24_and905_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and905_y0);
  and_gate and_gate_h_u_cla24_and906_y0(h_u_cla24_and905_y0, h_u_cla24_and904_y0, h_u_cla24_and906_y0);
  and_gate and_gate_h_u_cla24_and907_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and907_y0);
  and_gate and_gate_h_u_cla24_and908_y0(h_u_cla24_and907_y0, h_u_cla24_and906_y0, h_u_cla24_and908_y0);
  and_gate and_gate_h_u_cla24_and909_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and909_y0);
  and_gate and_gate_h_u_cla24_and910_y0(h_u_cla24_and909_y0, h_u_cla24_and908_y0, h_u_cla24_and910_y0);
  and_gate and_gate_h_u_cla24_and911_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and911_y0);
  and_gate and_gate_h_u_cla24_and912_y0(h_u_cla24_and911_y0, h_u_cla24_and910_y0, h_u_cla24_and912_y0);
  and_gate and_gate_h_u_cla24_and913_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and913_y0);
  and_gate and_gate_h_u_cla24_and914_y0(h_u_cla24_and913_y0, h_u_cla24_and912_y0, h_u_cla24_and914_y0);
  and_gate and_gate_h_u_cla24_and915_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and915_y0);
  and_gate and_gate_h_u_cla24_and916_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and916_y0);
  and_gate and_gate_h_u_cla24_and917_y0(h_u_cla24_and916_y0, h_u_cla24_and915_y0, h_u_cla24_and917_y0);
  and_gate and_gate_h_u_cla24_and918_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and918_y0);
  and_gate and_gate_h_u_cla24_and919_y0(h_u_cla24_and918_y0, h_u_cla24_and917_y0, h_u_cla24_and919_y0);
  and_gate and_gate_h_u_cla24_and920_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and920_y0);
  and_gate and_gate_h_u_cla24_and921_y0(h_u_cla24_and920_y0, h_u_cla24_and919_y0, h_u_cla24_and921_y0);
  and_gate and_gate_h_u_cla24_and922_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and922_y0);
  and_gate and_gate_h_u_cla24_and923_y0(h_u_cla24_and922_y0, h_u_cla24_and921_y0, h_u_cla24_and923_y0);
  and_gate and_gate_h_u_cla24_and924_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and924_y0);
  and_gate and_gate_h_u_cla24_and925_y0(h_u_cla24_and924_y0, h_u_cla24_and923_y0, h_u_cla24_and925_y0);
  and_gate and_gate_h_u_cla24_and926_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and926_y0);
  and_gate and_gate_h_u_cla24_and927_y0(h_u_cla24_and926_y0, h_u_cla24_and925_y0, h_u_cla24_and927_y0);
  and_gate and_gate_h_u_cla24_and928_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and928_y0);
  and_gate and_gate_h_u_cla24_and929_y0(h_u_cla24_and928_y0, h_u_cla24_and927_y0, h_u_cla24_and929_y0);
  and_gate and_gate_h_u_cla24_and930_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and930_y0);
  and_gate and_gate_h_u_cla24_and931_y0(h_u_cla24_and930_y0, h_u_cla24_and929_y0, h_u_cla24_and931_y0);
  and_gate and_gate_h_u_cla24_and932_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and932_y0);
  and_gate and_gate_h_u_cla24_and933_y0(h_u_cla24_and932_y0, h_u_cla24_and931_y0, h_u_cla24_and933_y0);
  and_gate and_gate_h_u_cla24_and934_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and934_y0);
  and_gate and_gate_h_u_cla24_and935_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and935_y0);
  and_gate and_gate_h_u_cla24_and936_y0(h_u_cla24_and935_y0, h_u_cla24_and934_y0, h_u_cla24_and936_y0);
  and_gate and_gate_h_u_cla24_and937_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and937_y0);
  and_gate and_gate_h_u_cla24_and938_y0(h_u_cla24_and937_y0, h_u_cla24_and936_y0, h_u_cla24_and938_y0);
  and_gate and_gate_h_u_cla24_and939_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and939_y0);
  and_gate and_gate_h_u_cla24_and940_y0(h_u_cla24_and939_y0, h_u_cla24_and938_y0, h_u_cla24_and940_y0);
  and_gate and_gate_h_u_cla24_and941_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and941_y0);
  and_gate and_gate_h_u_cla24_and942_y0(h_u_cla24_and941_y0, h_u_cla24_and940_y0, h_u_cla24_and942_y0);
  and_gate and_gate_h_u_cla24_and943_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and943_y0);
  and_gate and_gate_h_u_cla24_and944_y0(h_u_cla24_and943_y0, h_u_cla24_and942_y0, h_u_cla24_and944_y0);
  and_gate and_gate_h_u_cla24_and945_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and945_y0);
  and_gate and_gate_h_u_cla24_and946_y0(h_u_cla24_and945_y0, h_u_cla24_and944_y0, h_u_cla24_and946_y0);
  and_gate and_gate_h_u_cla24_and947_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and947_y0);
  and_gate and_gate_h_u_cla24_and948_y0(h_u_cla24_and947_y0, h_u_cla24_and946_y0, h_u_cla24_and948_y0);
  and_gate and_gate_h_u_cla24_and949_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and949_y0);
  and_gate and_gate_h_u_cla24_and950_y0(h_u_cla24_and949_y0, h_u_cla24_and948_y0, h_u_cla24_and950_y0);
  and_gate and_gate_h_u_cla24_and951_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and951_y0);
  and_gate and_gate_h_u_cla24_and952_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and952_y0);
  and_gate and_gate_h_u_cla24_and953_y0(h_u_cla24_and952_y0, h_u_cla24_and951_y0, h_u_cla24_and953_y0);
  and_gate and_gate_h_u_cla24_and954_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and954_y0);
  and_gate and_gate_h_u_cla24_and955_y0(h_u_cla24_and954_y0, h_u_cla24_and953_y0, h_u_cla24_and955_y0);
  and_gate and_gate_h_u_cla24_and956_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and956_y0);
  and_gate and_gate_h_u_cla24_and957_y0(h_u_cla24_and956_y0, h_u_cla24_and955_y0, h_u_cla24_and957_y0);
  and_gate and_gate_h_u_cla24_and958_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and958_y0);
  and_gate and_gate_h_u_cla24_and959_y0(h_u_cla24_and958_y0, h_u_cla24_and957_y0, h_u_cla24_and959_y0);
  and_gate and_gate_h_u_cla24_and960_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and960_y0);
  and_gate and_gate_h_u_cla24_and961_y0(h_u_cla24_and960_y0, h_u_cla24_and959_y0, h_u_cla24_and961_y0);
  and_gate and_gate_h_u_cla24_and962_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and962_y0);
  and_gate and_gate_h_u_cla24_and963_y0(h_u_cla24_and962_y0, h_u_cla24_and961_y0, h_u_cla24_and963_y0);
  and_gate and_gate_h_u_cla24_and964_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and964_y0);
  and_gate and_gate_h_u_cla24_and965_y0(h_u_cla24_and964_y0, h_u_cla24_and963_y0, h_u_cla24_and965_y0);
  and_gate and_gate_h_u_cla24_and966_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and966_y0);
  and_gate and_gate_h_u_cla24_and967_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and967_y0);
  and_gate and_gate_h_u_cla24_and968_y0(h_u_cla24_and967_y0, h_u_cla24_and966_y0, h_u_cla24_and968_y0);
  and_gate and_gate_h_u_cla24_and969_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and969_y0);
  and_gate and_gate_h_u_cla24_and970_y0(h_u_cla24_and969_y0, h_u_cla24_and968_y0, h_u_cla24_and970_y0);
  and_gate and_gate_h_u_cla24_and971_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and971_y0);
  and_gate and_gate_h_u_cla24_and972_y0(h_u_cla24_and971_y0, h_u_cla24_and970_y0, h_u_cla24_and972_y0);
  and_gate and_gate_h_u_cla24_and973_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and973_y0);
  and_gate and_gate_h_u_cla24_and974_y0(h_u_cla24_and973_y0, h_u_cla24_and972_y0, h_u_cla24_and974_y0);
  and_gate and_gate_h_u_cla24_and975_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and975_y0);
  and_gate and_gate_h_u_cla24_and976_y0(h_u_cla24_and975_y0, h_u_cla24_and974_y0, h_u_cla24_and976_y0);
  and_gate and_gate_h_u_cla24_and977_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and977_y0);
  and_gate and_gate_h_u_cla24_and978_y0(h_u_cla24_and977_y0, h_u_cla24_and976_y0, h_u_cla24_and978_y0);
  and_gate and_gate_h_u_cla24_and979_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and979_y0);
  and_gate and_gate_h_u_cla24_and980_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and980_y0);
  and_gate and_gate_h_u_cla24_and981_y0(h_u_cla24_and980_y0, h_u_cla24_and979_y0, h_u_cla24_and981_y0);
  and_gate and_gate_h_u_cla24_and982_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and982_y0);
  and_gate and_gate_h_u_cla24_and983_y0(h_u_cla24_and982_y0, h_u_cla24_and981_y0, h_u_cla24_and983_y0);
  and_gate and_gate_h_u_cla24_and984_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and984_y0);
  and_gate and_gate_h_u_cla24_and985_y0(h_u_cla24_and984_y0, h_u_cla24_and983_y0, h_u_cla24_and985_y0);
  and_gate and_gate_h_u_cla24_and986_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and986_y0);
  and_gate and_gate_h_u_cla24_and987_y0(h_u_cla24_and986_y0, h_u_cla24_and985_y0, h_u_cla24_and987_y0);
  and_gate and_gate_h_u_cla24_and988_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and988_y0);
  and_gate and_gate_h_u_cla24_and989_y0(h_u_cla24_and988_y0, h_u_cla24_and987_y0, h_u_cla24_and989_y0);
  and_gate and_gate_h_u_cla24_and990_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and990_y0);
  and_gate and_gate_h_u_cla24_and991_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and991_y0);
  and_gate and_gate_h_u_cla24_and992_y0(h_u_cla24_and991_y0, h_u_cla24_and990_y0, h_u_cla24_and992_y0);
  and_gate and_gate_h_u_cla24_and993_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and993_y0);
  and_gate and_gate_h_u_cla24_and994_y0(h_u_cla24_and993_y0, h_u_cla24_and992_y0, h_u_cla24_and994_y0);
  and_gate and_gate_h_u_cla24_and995_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and995_y0);
  and_gate and_gate_h_u_cla24_and996_y0(h_u_cla24_and995_y0, h_u_cla24_and994_y0, h_u_cla24_and996_y0);
  and_gate and_gate_h_u_cla24_and997_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and997_y0);
  and_gate and_gate_h_u_cla24_and998_y0(h_u_cla24_and997_y0, h_u_cla24_and996_y0, h_u_cla24_and998_y0);
  and_gate and_gate_h_u_cla24_and999_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and999_y0);
  and_gate and_gate_h_u_cla24_and1000_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1000_y0);
  and_gate and_gate_h_u_cla24_and1001_y0(h_u_cla24_and1000_y0, h_u_cla24_and999_y0, h_u_cla24_and1001_y0);
  and_gate and_gate_h_u_cla24_and1002_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1002_y0);
  and_gate and_gate_h_u_cla24_and1003_y0(h_u_cla24_and1002_y0, h_u_cla24_and1001_y0, h_u_cla24_and1003_y0);
  and_gate and_gate_h_u_cla24_and1004_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1004_y0);
  and_gate and_gate_h_u_cla24_and1005_y0(h_u_cla24_and1004_y0, h_u_cla24_and1003_y0, h_u_cla24_and1005_y0);
  and_gate and_gate_h_u_cla24_and1006_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1006_y0);
  and_gate and_gate_h_u_cla24_and1007_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1007_y0);
  and_gate and_gate_h_u_cla24_and1008_y0(h_u_cla24_and1007_y0, h_u_cla24_and1006_y0, h_u_cla24_and1008_y0);
  and_gate and_gate_h_u_cla24_and1009_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1009_y0);
  and_gate and_gate_h_u_cla24_and1010_y0(h_u_cla24_and1009_y0, h_u_cla24_and1008_y0, h_u_cla24_and1010_y0);
  and_gate and_gate_h_u_cla24_and1011_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1011_y0);
  and_gate and_gate_h_u_cla24_and1012_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1012_y0);
  and_gate and_gate_h_u_cla24_and1013_y0(h_u_cla24_and1012_y0, h_u_cla24_and1011_y0, h_u_cla24_and1013_y0);
  and_gate and_gate_h_u_cla24_and1014_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1014_y0);
  or_gate or_gate_h_u_cla24_or91_y0(h_u_cla24_and1014_y0, h_u_cla24_and845_y0, h_u_cla24_or91_y0);
  or_gate or_gate_h_u_cla24_or92_y0(h_u_cla24_or91_y0, h_u_cla24_and870_y0, h_u_cla24_or92_y0);
  or_gate or_gate_h_u_cla24_or93_y0(h_u_cla24_or92_y0, h_u_cla24_and893_y0, h_u_cla24_or93_y0);
  or_gate or_gate_h_u_cla24_or94_y0(h_u_cla24_or93_y0, h_u_cla24_and914_y0, h_u_cla24_or94_y0);
  or_gate or_gate_h_u_cla24_or95_y0(h_u_cla24_or94_y0, h_u_cla24_and933_y0, h_u_cla24_or95_y0);
  or_gate or_gate_h_u_cla24_or96_y0(h_u_cla24_or95_y0, h_u_cla24_and950_y0, h_u_cla24_or96_y0);
  or_gate or_gate_h_u_cla24_or97_y0(h_u_cla24_or96_y0, h_u_cla24_and965_y0, h_u_cla24_or97_y0);
  or_gate or_gate_h_u_cla24_or98_y0(h_u_cla24_or97_y0, h_u_cla24_and978_y0, h_u_cla24_or98_y0);
  or_gate or_gate_h_u_cla24_or99_y0(h_u_cla24_or98_y0, h_u_cla24_and989_y0, h_u_cla24_or99_y0);
  or_gate or_gate_h_u_cla24_or100_y0(h_u_cla24_or99_y0, h_u_cla24_and998_y0, h_u_cla24_or100_y0);
  or_gate or_gate_h_u_cla24_or101_y0(h_u_cla24_or100_y0, h_u_cla24_and1005_y0, h_u_cla24_or101_y0);
  or_gate or_gate_h_u_cla24_or102_y0(h_u_cla24_or101_y0, h_u_cla24_and1010_y0, h_u_cla24_or102_y0);
  or_gate or_gate_h_u_cla24_or103_y0(h_u_cla24_or102_y0, h_u_cla24_and1013_y0, h_u_cla24_or103_y0);
  or_gate or_gate_h_u_cla24_or104_y0(h_u_cla24_pg_logic13_y1, h_u_cla24_or103_y0, h_u_cla24_or104_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic14_y0(a_14, b_14, h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_pg_logic14_y2);
  xor_gate xor_gate_h_u_cla24_xor14_y0(h_u_cla24_pg_logic14_y2, h_u_cla24_or104_y0, h_u_cla24_xor14_y0);
  and_gate and_gate_h_u_cla24_and1015_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and1015_y0);
  and_gate and_gate_h_u_cla24_and1016_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and1016_y0);
  and_gate and_gate_h_u_cla24_and1017_y0(h_u_cla24_and1016_y0, h_u_cla24_and1015_y0, h_u_cla24_and1017_y0);
  and_gate and_gate_h_u_cla24_and1018_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and1018_y0);
  and_gate and_gate_h_u_cla24_and1019_y0(h_u_cla24_and1018_y0, h_u_cla24_and1017_y0, h_u_cla24_and1019_y0);
  and_gate and_gate_h_u_cla24_and1020_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and1020_y0);
  and_gate and_gate_h_u_cla24_and1021_y0(h_u_cla24_and1020_y0, h_u_cla24_and1019_y0, h_u_cla24_and1021_y0);
  and_gate and_gate_h_u_cla24_and1022_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and1022_y0);
  and_gate and_gate_h_u_cla24_and1023_y0(h_u_cla24_and1022_y0, h_u_cla24_and1021_y0, h_u_cla24_and1023_y0);
  and_gate and_gate_h_u_cla24_and1024_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and1024_y0);
  and_gate and_gate_h_u_cla24_and1025_y0(h_u_cla24_and1024_y0, h_u_cla24_and1023_y0, h_u_cla24_and1025_y0);
  and_gate and_gate_h_u_cla24_and1026_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and1026_y0);
  and_gate and_gate_h_u_cla24_and1027_y0(h_u_cla24_and1026_y0, h_u_cla24_and1025_y0, h_u_cla24_and1027_y0);
  and_gate and_gate_h_u_cla24_and1028_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and1028_y0);
  and_gate and_gate_h_u_cla24_and1029_y0(h_u_cla24_and1028_y0, h_u_cla24_and1027_y0, h_u_cla24_and1029_y0);
  and_gate and_gate_h_u_cla24_and1030_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and1030_y0);
  and_gate and_gate_h_u_cla24_and1031_y0(h_u_cla24_and1030_y0, h_u_cla24_and1029_y0, h_u_cla24_and1031_y0);
  and_gate and_gate_h_u_cla24_and1032_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and1032_y0);
  and_gate and_gate_h_u_cla24_and1033_y0(h_u_cla24_and1032_y0, h_u_cla24_and1031_y0, h_u_cla24_and1033_y0);
  and_gate and_gate_h_u_cla24_and1034_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and1034_y0);
  and_gate and_gate_h_u_cla24_and1035_y0(h_u_cla24_and1034_y0, h_u_cla24_and1033_y0, h_u_cla24_and1035_y0);
  and_gate and_gate_h_u_cla24_and1036_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and1036_y0);
  and_gate and_gate_h_u_cla24_and1037_y0(h_u_cla24_and1036_y0, h_u_cla24_and1035_y0, h_u_cla24_and1037_y0);
  and_gate and_gate_h_u_cla24_and1038_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and1038_y0);
  and_gate and_gate_h_u_cla24_and1039_y0(h_u_cla24_and1038_y0, h_u_cla24_and1037_y0, h_u_cla24_and1039_y0);
  and_gate and_gate_h_u_cla24_and1040_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and1040_y0);
  and_gate and_gate_h_u_cla24_and1041_y0(h_u_cla24_and1040_y0, h_u_cla24_and1039_y0, h_u_cla24_and1041_y0);
  and_gate and_gate_h_u_cla24_and1042_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and1042_y0);
  and_gate and_gate_h_u_cla24_and1043_y0(h_u_cla24_and1042_y0, h_u_cla24_and1041_y0, h_u_cla24_and1043_y0);
  and_gate and_gate_h_u_cla24_and1044_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1044_y0);
  and_gate and_gate_h_u_cla24_and1045_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1045_y0);
  and_gate and_gate_h_u_cla24_and1046_y0(h_u_cla24_and1045_y0, h_u_cla24_and1044_y0, h_u_cla24_and1046_y0);
  and_gate and_gate_h_u_cla24_and1047_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1047_y0);
  and_gate and_gate_h_u_cla24_and1048_y0(h_u_cla24_and1047_y0, h_u_cla24_and1046_y0, h_u_cla24_and1048_y0);
  and_gate and_gate_h_u_cla24_and1049_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1049_y0);
  and_gate and_gate_h_u_cla24_and1050_y0(h_u_cla24_and1049_y0, h_u_cla24_and1048_y0, h_u_cla24_and1050_y0);
  and_gate and_gate_h_u_cla24_and1051_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1051_y0);
  and_gate and_gate_h_u_cla24_and1052_y0(h_u_cla24_and1051_y0, h_u_cla24_and1050_y0, h_u_cla24_and1052_y0);
  and_gate and_gate_h_u_cla24_and1053_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1053_y0);
  and_gate and_gate_h_u_cla24_and1054_y0(h_u_cla24_and1053_y0, h_u_cla24_and1052_y0, h_u_cla24_and1054_y0);
  and_gate and_gate_h_u_cla24_and1055_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1055_y0);
  and_gate and_gate_h_u_cla24_and1056_y0(h_u_cla24_and1055_y0, h_u_cla24_and1054_y0, h_u_cla24_and1056_y0);
  and_gate and_gate_h_u_cla24_and1057_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1057_y0);
  and_gate and_gate_h_u_cla24_and1058_y0(h_u_cla24_and1057_y0, h_u_cla24_and1056_y0, h_u_cla24_and1058_y0);
  and_gate and_gate_h_u_cla24_and1059_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1059_y0);
  and_gate and_gate_h_u_cla24_and1060_y0(h_u_cla24_and1059_y0, h_u_cla24_and1058_y0, h_u_cla24_and1060_y0);
  and_gate and_gate_h_u_cla24_and1061_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1061_y0);
  and_gate and_gate_h_u_cla24_and1062_y0(h_u_cla24_and1061_y0, h_u_cla24_and1060_y0, h_u_cla24_and1062_y0);
  and_gate and_gate_h_u_cla24_and1063_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1063_y0);
  and_gate and_gate_h_u_cla24_and1064_y0(h_u_cla24_and1063_y0, h_u_cla24_and1062_y0, h_u_cla24_and1064_y0);
  and_gate and_gate_h_u_cla24_and1065_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1065_y0);
  and_gate and_gate_h_u_cla24_and1066_y0(h_u_cla24_and1065_y0, h_u_cla24_and1064_y0, h_u_cla24_and1066_y0);
  and_gate and_gate_h_u_cla24_and1067_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1067_y0);
  and_gate and_gate_h_u_cla24_and1068_y0(h_u_cla24_and1067_y0, h_u_cla24_and1066_y0, h_u_cla24_and1068_y0);
  and_gate and_gate_h_u_cla24_and1069_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1069_y0);
  and_gate and_gate_h_u_cla24_and1070_y0(h_u_cla24_and1069_y0, h_u_cla24_and1068_y0, h_u_cla24_and1070_y0);
  and_gate and_gate_h_u_cla24_and1071_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1071_y0);
  and_gate and_gate_h_u_cla24_and1072_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1072_y0);
  and_gate and_gate_h_u_cla24_and1073_y0(h_u_cla24_and1072_y0, h_u_cla24_and1071_y0, h_u_cla24_and1073_y0);
  and_gate and_gate_h_u_cla24_and1074_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1074_y0);
  and_gate and_gate_h_u_cla24_and1075_y0(h_u_cla24_and1074_y0, h_u_cla24_and1073_y0, h_u_cla24_and1075_y0);
  and_gate and_gate_h_u_cla24_and1076_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1076_y0);
  and_gate and_gate_h_u_cla24_and1077_y0(h_u_cla24_and1076_y0, h_u_cla24_and1075_y0, h_u_cla24_and1077_y0);
  and_gate and_gate_h_u_cla24_and1078_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1078_y0);
  and_gate and_gate_h_u_cla24_and1079_y0(h_u_cla24_and1078_y0, h_u_cla24_and1077_y0, h_u_cla24_and1079_y0);
  and_gate and_gate_h_u_cla24_and1080_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1080_y0);
  and_gate and_gate_h_u_cla24_and1081_y0(h_u_cla24_and1080_y0, h_u_cla24_and1079_y0, h_u_cla24_and1081_y0);
  and_gate and_gate_h_u_cla24_and1082_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1082_y0);
  and_gate and_gate_h_u_cla24_and1083_y0(h_u_cla24_and1082_y0, h_u_cla24_and1081_y0, h_u_cla24_and1083_y0);
  and_gate and_gate_h_u_cla24_and1084_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1084_y0);
  and_gate and_gate_h_u_cla24_and1085_y0(h_u_cla24_and1084_y0, h_u_cla24_and1083_y0, h_u_cla24_and1085_y0);
  and_gate and_gate_h_u_cla24_and1086_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1086_y0);
  and_gate and_gate_h_u_cla24_and1087_y0(h_u_cla24_and1086_y0, h_u_cla24_and1085_y0, h_u_cla24_and1087_y0);
  and_gate and_gate_h_u_cla24_and1088_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1088_y0);
  and_gate and_gate_h_u_cla24_and1089_y0(h_u_cla24_and1088_y0, h_u_cla24_and1087_y0, h_u_cla24_and1089_y0);
  and_gate and_gate_h_u_cla24_and1090_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1090_y0);
  and_gate and_gate_h_u_cla24_and1091_y0(h_u_cla24_and1090_y0, h_u_cla24_and1089_y0, h_u_cla24_and1091_y0);
  and_gate and_gate_h_u_cla24_and1092_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1092_y0);
  and_gate and_gate_h_u_cla24_and1093_y0(h_u_cla24_and1092_y0, h_u_cla24_and1091_y0, h_u_cla24_and1093_y0);
  and_gate and_gate_h_u_cla24_and1094_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1094_y0);
  and_gate and_gate_h_u_cla24_and1095_y0(h_u_cla24_and1094_y0, h_u_cla24_and1093_y0, h_u_cla24_and1095_y0);
  and_gate and_gate_h_u_cla24_and1096_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1096_y0);
  and_gate and_gate_h_u_cla24_and1097_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1097_y0);
  and_gate and_gate_h_u_cla24_and1098_y0(h_u_cla24_and1097_y0, h_u_cla24_and1096_y0, h_u_cla24_and1098_y0);
  and_gate and_gate_h_u_cla24_and1099_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1099_y0);
  and_gate and_gate_h_u_cla24_and1100_y0(h_u_cla24_and1099_y0, h_u_cla24_and1098_y0, h_u_cla24_and1100_y0);
  and_gate and_gate_h_u_cla24_and1101_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1101_y0);
  and_gate and_gate_h_u_cla24_and1102_y0(h_u_cla24_and1101_y0, h_u_cla24_and1100_y0, h_u_cla24_and1102_y0);
  and_gate and_gate_h_u_cla24_and1103_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1103_y0);
  and_gate and_gate_h_u_cla24_and1104_y0(h_u_cla24_and1103_y0, h_u_cla24_and1102_y0, h_u_cla24_and1104_y0);
  and_gate and_gate_h_u_cla24_and1105_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1105_y0);
  and_gate and_gate_h_u_cla24_and1106_y0(h_u_cla24_and1105_y0, h_u_cla24_and1104_y0, h_u_cla24_and1106_y0);
  and_gate and_gate_h_u_cla24_and1107_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1107_y0);
  and_gate and_gate_h_u_cla24_and1108_y0(h_u_cla24_and1107_y0, h_u_cla24_and1106_y0, h_u_cla24_and1108_y0);
  and_gate and_gate_h_u_cla24_and1109_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1109_y0);
  and_gate and_gate_h_u_cla24_and1110_y0(h_u_cla24_and1109_y0, h_u_cla24_and1108_y0, h_u_cla24_and1110_y0);
  and_gate and_gate_h_u_cla24_and1111_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1111_y0);
  and_gate and_gate_h_u_cla24_and1112_y0(h_u_cla24_and1111_y0, h_u_cla24_and1110_y0, h_u_cla24_and1112_y0);
  and_gate and_gate_h_u_cla24_and1113_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1113_y0);
  and_gate and_gate_h_u_cla24_and1114_y0(h_u_cla24_and1113_y0, h_u_cla24_and1112_y0, h_u_cla24_and1114_y0);
  and_gate and_gate_h_u_cla24_and1115_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1115_y0);
  and_gate and_gate_h_u_cla24_and1116_y0(h_u_cla24_and1115_y0, h_u_cla24_and1114_y0, h_u_cla24_and1116_y0);
  and_gate and_gate_h_u_cla24_and1117_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1117_y0);
  and_gate and_gate_h_u_cla24_and1118_y0(h_u_cla24_and1117_y0, h_u_cla24_and1116_y0, h_u_cla24_and1118_y0);
  and_gate and_gate_h_u_cla24_and1119_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1119_y0);
  and_gate and_gate_h_u_cla24_and1120_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1120_y0);
  and_gate and_gate_h_u_cla24_and1121_y0(h_u_cla24_and1120_y0, h_u_cla24_and1119_y0, h_u_cla24_and1121_y0);
  and_gate and_gate_h_u_cla24_and1122_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1122_y0);
  and_gate and_gate_h_u_cla24_and1123_y0(h_u_cla24_and1122_y0, h_u_cla24_and1121_y0, h_u_cla24_and1123_y0);
  and_gate and_gate_h_u_cla24_and1124_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1124_y0);
  and_gate and_gate_h_u_cla24_and1125_y0(h_u_cla24_and1124_y0, h_u_cla24_and1123_y0, h_u_cla24_and1125_y0);
  and_gate and_gate_h_u_cla24_and1126_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1126_y0);
  and_gate and_gate_h_u_cla24_and1127_y0(h_u_cla24_and1126_y0, h_u_cla24_and1125_y0, h_u_cla24_and1127_y0);
  and_gate and_gate_h_u_cla24_and1128_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1128_y0);
  and_gate and_gate_h_u_cla24_and1129_y0(h_u_cla24_and1128_y0, h_u_cla24_and1127_y0, h_u_cla24_and1129_y0);
  and_gate and_gate_h_u_cla24_and1130_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1130_y0);
  and_gate and_gate_h_u_cla24_and1131_y0(h_u_cla24_and1130_y0, h_u_cla24_and1129_y0, h_u_cla24_and1131_y0);
  and_gate and_gate_h_u_cla24_and1132_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1132_y0);
  and_gate and_gate_h_u_cla24_and1133_y0(h_u_cla24_and1132_y0, h_u_cla24_and1131_y0, h_u_cla24_and1133_y0);
  and_gate and_gate_h_u_cla24_and1134_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1134_y0);
  and_gate and_gate_h_u_cla24_and1135_y0(h_u_cla24_and1134_y0, h_u_cla24_and1133_y0, h_u_cla24_and1135_y0);
  and_gate and_gate_h_u_cla24_and1136_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1136_y0);
  and_gate and_gate_h_u_cla24_and1137_y0(h_u_cla24_and1136_y0, h_u_cla24_and1135_y0, h_u_cla24_and1137_y0);
  and_gate and_gate_h_u_cla24_and1138_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1138_y0);
  and_gate and_gate_h_u_cla24_and1139_y0(h_u_cla24_and1138_y0, h_u_cla24_and1137_y0, h_u_cla24_and1139_y0);
  and_gate and_gate_h_u_cla24_and1140_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1140_y0);
  and_gate and_gate_h_u_cla24_and1141_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1141_y0);
  and_gate and_gate_h_u_cla24_and1142_y0(h_u_cla24_and1141_y0, h_u_cla24_and1140_y0, h_u_cla24_and1142_y0);
  and_gate and_gate_h_u_cla24_and1143_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1143_y0);
  and_gate and_gate_h_u_cla24_and1144_y0(h_u_cla24_and1143_y0, h_u_cla24_and1142_y0, h_u_cla24_and1144_y0);
  and_gate and_gate_h_u_cla24_and1145_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1145_y0);
  and_gate and_gate_h_u_cla24_and1146_y0(h_u_cla24_and1145_y0, h_u_cla24_and1144_y0, h_u_cla24_and1146_y0);
  and_gate and_gate_h_u_cla24_and1147_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1147_y0);
  and_gate and_gate_h_u_cla24_and1148_y0(h_u_cla24_and1147_y0, h_u_cla24_and1146_y0, h_u_cla24_and1148_y0);
  and_gate and_gate_h_u_cla24_and1149_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1149_y0);
  and_gate and_gate_h_u_cla24_and1150_y0(h_u_cla24_and1149_y0, h_u_cla24_and1148_y0, h_u_cla24_and1150_y0);
  and_gate and_gate_h_u_cla24_and1151_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1151_y0);
  and_gate and_gate_h_u_cla24_and1152_y0(h_u_cla24_and1151_y0, h_u_cla24_and1150_y0, h_u_cla24_and1152_y0);
  and_gate and_gate_h_u_cla24_and1153_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1153_y0);
  and_gate and_gate_h_u_cla24_and1154_y0(h_u_cla24_and1153_y0, h_u_cla24_and1152_y0, h_u_cla24_and1154_y0);
  and_gate and_gate_h_u_cla24_and1155_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1155_y0);
  and_gate and_gate_h_u_cla24_and1156_y0(h_u_cla24_and1155_y0, h_u_cla24_and1154_y0, h_u_cla24_and1156_y0);
  and_gate and_gate_h_u_cla24_and1157_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1157_y0);
  and_gate and_gate_h_u_cla24_and1158_y0(h_u_cla24_and1157_y0, h_u_cla24_and1156_y0, h_u_cla24_and1158_y0);
  and_gate and_gate_h_u_cla24_and1159_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1159_y0);
  and_gate and_gate_h_u_cla24_and1160_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1160_y0);
  and_gate and_gate_h_u_cla24_and1161_y0(h_u_cla24_and1160_y0, h_u_cla24_and1159_y0, h_u_cla24_and1161_y0);
  and_gate and_gate_h_u_cla24_and1162_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1162_y0);
  and_gate and_gate_h_u_cla24_and1163_y0(h_u_cla24_and1162_y0, h_u_cla24_and1161_y0, h_u_cla24_and1163_y0);
  and_gate and_gate_h_u_cla24_and1164_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1164_y0);
  and_gate and_gate_h_u_cla24_and1165_y0(h_u_cla24_and1164_y0, h_u_cla24_and1163_y0, h_u_cla24_and1165_y0);
  and_gate and_gate_h_u_cla24_and1166_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1166_y0);
  and_gate and_gate_h_u_cla24_and1167_y0(h_u_cla24_and1166_y0, h_u_cla24_and1165_y0, h_u_cla24_and1167_y0);
  and_gate and_gate_h_u_cla24_and1168_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1168_y0);
  and_gate and_gate_h_u_cla24_and1169_y0(h_u_cla24_and1168_y0, h_u_cla24_and1167_y0, h_u_cla24_and1169_y0);
  and_gate and_gate_h_u_cla24_and1170_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1170_y0);
  and_gate and_gate_h_u_cla24_and1171_y0(h_u_cla24_and1170_y0, h_u_cla24_and1169_y0, h_u_cla24_and1171_y0);
  and_gate and_gate_h_u_cla24_and1172_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1172_y0);
  and_gate and_gate_h_u_cla24_and1173_y0(h_u_cla24_and1172_y0, h_u_cla24_and1171_y0, h_u_cla24_and1173_y0);
  and_gate and_gate_h_u_cla24_and1174_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1174_y0);
  and_gate and_gate_h_u_cla24_and1175_y0(h_u_cla24_and1174_y0, h_u_cla24_and1173_y0, h_u_cla24_and1175_y0);
  and_gate and_gate_h_u_cla24_and1176_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1176_y0);
  and_gate and_gate_h_u_cla24_and1177_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1177_y0);
  and_gate and_gate_h_u_cla24_and1178_y0(h_u_cla24_and1177_y0, h_u_cla24_and1176_y0, h_u_cla24_and1178_y0);
  and_gate and_gate_h_u_cla24_and1179_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1179_y0);
  and_gate and_gate_h_u_cla24_and1180_y0(h_u_cla24_and1179_y0, h_u_cla24_and1178_y0, h_u_cla24_and1180_y0);
  and_gate and_gate_h_u_cla24_and1181_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1181_y0);
  and_gate and_gate_h_u_cla24_and1182_y0(h_u_cla24_and1181_y0, h_u_cla24_and1180_y0, h_u_cla24_and1182_y0);
  and_gate and_gate_h_u_cla24_and1183_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1183_y0);
  and_gate and_gate_h_u_cla24_and1184_y0(h_u_cla24_and1183_y0, h_u_cla24_and1182_y0, h_u_cla24_and1184_y0);
  and_gate and_gate_h_u_cla24_and1185_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1185_y0);
  and_gate and_gate_h_u_cla24_and1186_y0(h_u_cla24_and1185_y0, h_u_cla24_and1184_y0, h_u_cla24_and1186_y0);
  and_gate and_gate_h_u_cla24_and1187_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1187_y0);
  and_gate and_gate_h_u_cla24_and1188_y0(h_u_cla24_and1187_y0, h_u_cla24_and1186_y0, h_u_cla24_and1188_y0);
  and_gate and_gate_h_u_cla24_and1189_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1189_y0);
  and_gate and_gate_h_u_cla24_and1190_y0(h_u_cla24_and1189_y0, h_u_cla24_and1188_y0, h_u_cla24_and1190_y0);
  and_gate and_gate_h_u_cla24_and1191_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1191_y0);
  and_gate and_gate_h_u_cla24_and1192_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1192_y0);
  and_gate and_gate_h_u_cla24_and1193_y0(h_u_cla24_and1192_y0, h_u_cla24_and1191_y0, h_u_cla24_and1193_y0);
  and_gate and_gate_h_u_cla24_and1194_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1194_y0);
  and_gate and_gate_h_u_cla24_and1195_y0(h_u_cla24_and1194_y0, h_u_cla24_and1193_y0, h_u_cla24_and1195_y0);
  and_gate and_gate_h_u_cla24_and1196_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1196_y0);
  and_gate and_gate_h_u_cla24_and1197_y0(h_u_cla24_and1196_y0, h_u_cla24_and1195_y0, h_u_cla24_and1197_y0);
  and_gate and_gate_h_u_cla24_and1198_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1198_y0);
  and_gate and_gate_h_u_cla24_and1199_y0(h_u_cla24_and1198_y0, h_u_cla24_and1197_y0, h_u_cla24_and1199_y0);
  and_gate and_gate_h_u_cla24_and1200_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1200_y0);
  and_gate and_gate_h_u_cla24_and1201_y0(h_u_cla24_and1200_y0, h_u_cla24_and1199_y0, h_u_cla24_and1201_y0);
  and_gate and_gate_h_u_cla24_and1202_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1202_y0);
  and_gate and_gate_h_u_cla24_and1203_y0(h_u_cla24_and1202_y0, h_u_cla24_and1201_y0, h_u_cla24_and1203_y0);
  and_gate and_gate_h_u_cla24_and1204_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1204_y0);
  and_gate and_gate_h_u_cla24_and1205_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1205_y0);
  and_gate and_gate_h_u_cla24_and1206_y0(h_u_cla24_and1205_y0, h_u_cla24_and1204_y0, h_u_cla24_and1206_y0);
  and_gate and_gate_h_u_cla24_and1207_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1207_y0);
  and_gate and_gate_h_u_cla24_and1208_y0(h_u_cla24_and1207_y0, h_u_cla24_and1206_y0, h_u_cla24_and1208_y0);
  and_gate and_gate_h_u_cla24_and1209_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1209_y0);
  and_gate and_gate_h_u_cla24_and1210_y0(h_u_cla24_and1209_y0, h_u_cla24_and1208_y0, h_u_cla24_and1210_y0);
  and_gate and_gate_h_u_cla24_and1211_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1211_y0);
  and_gate and_gate_h_u_cla24_and1212_y0(h_u_cla24_and1211_y0, h_u_cla24_and1210_y0, h_u_cla24_and1212_y0);
  and_gate and_gate_h_u_cla24_and1213_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1213_y0);
  and_gate and_gate_h_u_cla24_and1214_y0(h_u_cla24_and1213_y0, h_u_cla24_and1212_y0, h_u_cla24_and1214_y0);
  and_gate and_gate_h_u_cla24_and1215_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1215_y0);
  and_gate and_gate_h_u_cla24_and1216_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1216_y0);
  and_gate and_gate_h_u_cla24_and1217_y0(h_u_cla24_and1216_y0, h_u_cla24_and1215_y0, h_u_cla24_and1217_y0);
  and_gate and_gate_h_u_cla24_and1218_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1218_y0);
  and_gate and_gate_h_u_cla24_and1219_y0(h_u_cla24_and1218_y0, h_u_cla24_and1217_y0, h_u_cla24_and1219_y0);
  and_gate and_gate_h_u_cla24_and1220_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1220_y0);
  and_gate and_gate_h_u_cla24_and1221_y0(h_u_cla24_and1220_y0, h_u_cla24_and1219_y0, h_u_cla24_and1221_y0);
  and_gate and_gate_h_u_cla24_and1222_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1222_y0);
  and_gate and_gate_h_u_cla24_and1223_y0(h_u_cla24_and1222_y0, h_u_cla24_and1221_y0, h_u_cla24_and1223_y0);
  and_gate and_gate_h_u_cla24_and1224_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1224_y0);
  and_gate and_gate_h_u_cla24_and1225_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1225_y0);
  and_gate and_gate_h_u_cla24_and1226_y0(h_u_cla24_and1225_y0, h_u_cla24_and1224_y0, h_u_cla24_and1226_y0);
  and_gate and_gate_h_u_cla24_and1227_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1227_y0);
  and_gate and_gate_h_u_cla24_and1228_y0(h_u_cla24_and1227_y0, h_u_cla24_and1226_y0, h_u_cla24_and1228_y0);
  and_gate and_gate_h_u_cla24_and1229_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1229_y0);
  and_gate and_gate_h_u_cla24_and1230_y0(h_u_cla24_and1229_y0, h_u_cla24_and1228_y0, h_u_cla24_and1230_y0);
  and_gate and_gate_h_u_cla24_and1231_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1231_y0);
  and_gate and_gate_h_u_cla24_and1232_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1232_y0);
  and_gate and_gate_h_u_cla24_and1233_y0(h_u_cla24_and1232_y0, h_u_cla24_and1231_y0, h_u_cla24_and1233_y0);
  and_gate and_gate_h_u_cla24_and1234_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1234_y0);
  and_gate and_gate_h_u_cla24_and1235_y0(h_u_cla24_and1234_y0, h_u_cla24_and1233_y0, h_u_cla24_and1235_y0);
  and_gate and_gate_h_u_cla24_and1236_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1236_y0);
  and_gate and_gate_h_u_cla24_and1237_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1237_y0);
  and_gate and_gate_h_u_cla24_and1238_y0(h_u_cla24_and1237_y0, h_u_cla24_and1236_y0, h_u_cla24_and1238_y0);
  and_gate and_gate_h_u_cla24_and1239_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and1239_y0);
  or_gate or_gate_h_u_cla24_or105_y0(h_u_cla24_and1239_y0, h_u_cla24_and1043_y0, h_u_cla24_or105_y0);
  or_gate or_gate_h_u_cla24_or106_y0(h_u_cla24_or105_y0, h_u_cla24_and1070_y0, h_u_cla24_or106_y0);
  or_gate or_gate_h_u_cla24_or107_y0(h_u_cla24_or106_y0, h_u_cla24_and1095_y0, h_u_cla24_or107_y0);
  or_gate or_gate_h_u_cla24_or108_y0(h_u_cla24_or107_y0, h_u_cla24_and1118_y0, h_u_cla24_or108_y0);
  or_gate or_gate_h_u_cla24_or109_y0(h_u_cla24_or108_y0, h_u_cla24_and1139_y0, h_u_cla24_or109_y0);
  or_gate or_gate_h_u_cla24_or110_y0(h_u_cla24_or109_y0, h_u_cla24_and1158_y0, h_u_cla24_or110_y0);
  or_gate or_gate_h_u_cla24_or111_y0(h_u_cla24_or110_y0, h_u_cla24_and1175_y0, h_u_cla24_or111_y0);
  or_gate or_gate_h_u_cla24_or112_y0(h_u_cla24_or111_y0, h_u_cla24_and1190_y0, h_u_cla24_or112_y0);
  or_gate or_gate_h_u_cla24_or113_y0(h_u_cla24_or112_y0, h_u_cla24_and1203_y0, h_u_cla24_or113_y0);
  or_gate or_gate_h_u_cla24_or114_y0(h_u_cla24_or113_y0, h_u_cla24_and1214_y0, h_u_cla24_or114_y0);
  or_gate or_gate_h_u_cla24_or115_y0(h_u_cla24_or114_y0, h_u_cla24_and1223_y0, h_u_cla24_or115_y0);
  or_gate or_gate_h_u_cla24_or116_y0(h_u_cla24_or115_y0, h_u_cla24_and1230_y0, h_u_cla24_or116_y0);
  or_gate or_gate_h_u_cla24_or117_y0(h_u_cla24_or116_y0, h_u_cla24_and1235_y0, h_u_cla24_or117_y0);
  or_gate or_gate_h_u_cla24_or118_y0(h_u_cla24_or117_y0, h_u_cla24_and1238_y0, h_u_cla24_or118_y0);
  or_gate or_gate_h_u_cla24_or119_y0(h_u_cla24_pg_logic14_y1, h_u_cla24_or118_y0, h_u_cla24_or119_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic15_y0(a_15, b_15, h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_pg_logic15_y2);
  xor_gate xor_gate_h_u_cla24_xor15_y0(h_u_cla24_pg_logic15_y2, h_u_cla24_or119_y0, h_u_cla24_xor15_y0);
  and_gate and_gate_h_u_cla24_and1240_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and1240_y0);
  and_gate and_gate_h_u_cla24_and1241_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and1241_y0);
  and_gate and_gate_h_u_cla24_and1242_y0(h_u_cla24_and1241_y0, h_u_cla24_and1240_y0, h_u_cla24_and1242_y0);
  and_gate and_gate_h_u_cla24_and1243_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and1243_y0);
  and_gate and_gate_h_u_cla24_and1244_y0(h_u_cla24_and1243_y0, h_u_cla24_and1242_y0, h_u_cla24_and1244_y0);
  and_gate and_gate_h_u_cla24_and1245_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and1245_y0);
  and_gate and_gate_h_u_cla24_and1246_y0(h_u_cla24_and1245_y0, h_u_cla24_and1244_y0, h_u_cla24_and1246_y0);
  and_gate and_gate_h_u_cla24_and1247_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and1247_y0);
  and_gate and_gate_h_u_cla24_and1248_y0(h_u_cla24_and1247_y0, h_u_cla24_and1246_y0, h_u_cla24_and1248_y0);
  and_gate and_gate_h_u_cla24_and1249_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and1249_y0);
  and_gate and_gate_h_u_cla24_and1250_y0(h_u_cla24_and1249_y0, h_u_cla24_and1248_y0, h_u_cla24_and1250_y0);
  and_gate and_gate_h_u_cla24_and1251_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and1251_y0);
  and_gate and_gate_h_u_cla24_and1252_y0(h_u_cla24_and1251_y0, h_u_cla24_and1250_y0, h_u_cla24_and1252_y0);
  and_gate and_gate_h_u_cla24_and1253_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and1253_y0);
  and_gate and_gate_h_u_cla24_and1254_y0(h_u_cla24_and1253_y0, h_u_cla24_and1252_y0, h_u_cla24_and1254_y0);
  and_gate and_gate_h_u_cla24_and1255_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and1255_y0);
  and_gate and_gate_h_u_cla24_and1256_y0(h_u_cla24_and1255_y0, h_u_cla24_and1254_y0, h_u_cla24_and1256_y0);
  and_gate and_gate_h_u_cla24_and1257_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and1257_y0);
  and_gate and_gate_h_u_cla24_and1258_y0(h_u_cla24_and1257_y0, h_u_cla24_and1256_y0, h_u_cla24_and1258_y0);
  and_gate and_gate_h_u_cla24_and1259_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and1259_y0);
  and_gate and_gate_h_u_cla24_and1260_y0(h_u_cla24_and1259_y0, h_u_cla24_and1258_y0, h_u_cla24_and1260_y0);
  and_gate and_gate_h_u_cla24_and1261_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and1261_y0);
  and_gate and_gate_h_u_cla24_and1262_y0(h_u_cla24_and1261_y0, h_u_cla24_and1260_y0, h_u_cla24_and1262_y0);
  and_gate and_gate_h_u_cla24_and1263_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and1263_y0);
  and_gate and_gate_h_u_cla24_and1264_y0(h_u_cla24_and1263_y0, h_u_cla24_and1262_y0, h_u_cla24_and1264_y0);
  and_gate and_gate_h_u_cla24_and1265_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and1265_y0);
  and_gate and_gate_h_u_cla24_and1266_y0(h_u_cla24_and1265_y0, h_u_cla24_and1264_y0, h_u_cla24_and1266_y0);
  and_gate and_gate_h_u_cla24_and1267_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and1267_y0);
  and_gate and_gate_h_u_cla24_and1268_y0(h_u_cla24_and1267_y0, h_u_cla24_and1266_y0, h_u_cla24_and1268_y0);
  and_gate and_gate_h_u_cla24_and1269_y0(h_u_cla24_pg_logic15_y0, constant_wire_0, h_u_cla24_and1269_y0);
  and_gate and_gate_h_u_cla24_and1270_y0(h_u_cla24_and1269_y0, h_u_cla24_and1268_y0, h_u_cla24_and1270_y0);
  and_gate and_gate_h_u_cla24_and1271_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1271_y0);
  and_gate and_gate_h_u_cla24_and1272_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1272_y0);
  and_gate and_gate_h_u_cla24_and1273_y0(h_u_cla24_and1272_y0, h_u_cla24_and1271_y0, h_u_cla24_and1273_y0);
  and_gate and_gate_h_u_cla24_and1274_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1274_y0);
  and_gate and_gate_h_u_cla24_and1275_y0(h_u_cla24_and1274_y0, h_u_cla24_and1273_y0, h_u_cla24_and1275_y0);
  and_gate and_gate_h_u_cla24_and1276_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1276_y0);
  and_gate and_gate_h_u_cla24_and1277_y0(h_u_cla24_and1276_y0, h_u_cla24_and1275_y0, h_u_cla24_and1277_y0);
  and_gate and_gate_h_u_cla24_and1278_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1278_y0);
  and_gate and_gate_h_u_cla24_and1279_y0(h_u_cla24_and1278_y0, h_u_cla24_and1277_y0, h_u_cla24_and1279_y0);
  and_gate and_gate_h_u_cla24_and1280_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1280_y0);
  and_gate and_gate_h_u_cla24_and1281_y0(h_u_cla24_and1280_y0, h_u_cla24_and1279_y0, h_u_cla24_and1281_y0);
  and_gate and_gate_h_u_cla24_and1282_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1282_y0);
  and_gate and_gate_h_u_cla24_and1283_y0(h_u_cla24_and1282_y0, h_u_cla24_and1281_y0, h_u_cla24_and1283_y0);
  and_gate and_gate_h_u_cla24_and1284_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1284_y0);
  and_gate and_gate_h_u_cla24_and1285_y0(h_u_cla24_and1284_y0, h_u_cla24_and1283_y0, h_u_cla24_and1285_y0);
  and_gate and_gate_h_u_cla24_and1286_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1286_y0);
  and_gate and_gate_h_u_cla24_and1287_y0(h_u_cla24_and1286_y0, h_u_cla24_and1285_y0, h_u_cla24_and1287_y0);
  and_gate and_gate_h_u_cla24_and1288_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1288_y0);
  and_gate and_gate_h_u_cla24_and1289_y0(h_u_cla24_and1288_y0, h_u_cla24_and1287_y0, h_u_cla24_and1289_y0);
  and_gate and_gate_h_u_cla24_and1290_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1290_y0);
  and_gate and_gate_h_u_cla24_and1291_y0(h_u_cla24_and1290_y0, h_u_cla24_and1289_y0, h_u_cla24_and1291_y0);
  and_gate and_gate_h_u_cla24_and1292_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1292_y0);
  and_gate and_gate_h_u_cla24_and1293_y0(h_u_cla24_and1292_y0, h_u_cla24_and1291_y0, h_u_cla24_and1293_y0);
  and_gate and_gate_h_u_cla24_and1294_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1294_y0);
  and_gate and_gate_h_u_cla24_and1295_y0(h_u_cla24_and1294_y0, h_u_cla24_and1293_y0, h_u_cla24_and1295_y0);
  and_gate and_gate_h_u_cla24_and1296_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1296_y0);
  and_gate and_gate_h_u_cla24_and1297_y0(h_u_cla24_and1296_y0, h_u_cla24_and1295_y0, h_u_cla24_and1297_y0);
  and_gate and_gate_h_u_cla24_and1298_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1298_y0);
  and_gate and_gate_h_u_cla24_and1299_y0(h_u_cla24_and1298_y0, h_u_cla24_and1297_y0, h_u_cla24_and1299_y0);
  and_gate and_gate_h_u_cla24_and1300_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1300_y0);
  and_gate and_gate_h_u_cla24_and1301_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1301_y0);
  and_gate and_gate_h_u_cla24_and1302_y0(h_u_cla24_and1301_y0, h_u_cla24_and1300_y0, h_u_cla24_and1302_y0);
  and_gate and_gate_h_u_cla24_and1303_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1303_y0);
  and_gate and_gate_h_u_cla24_and1304_y0(h_u_cla24_and1303_y0, h_u_cla24_and1302_y0, h_u_cla24_and1304_y0);
  and_gate and_gate_h_u_cla24_and1305_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1305_y0);
  and_gate and_gate_h_u_cla24_and1306_y0(h_u_cla24_and1305_y0, h_u_cla24_and1304_y0, h_u_cla24_and1306_y0);
  and_gate and_gate_h_u_cla24_and1307_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1307_y0);
  and_gate and_gate_h_u_cla24_and1308_y0(h_u_cla24_and1307_y0, h_u_cla24_and1306_y0, h_u_cla24_and1308_y0);
  and_gate and_gate_h_u_cla24_and1309_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1309_y0);
  and_gate and_gate_h_u_cla24_and1310_y0(h_u_cla24_and1309_y0, h_u_cla24_and1308_y0, h_u_cla24_and1310_y0);
  and_gate and_gate_h_u_cla24_and1311_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1311_y0);
  and_gate and_gate_h_u_cla24_and1312_y0(h_u_cla24_and1311_y0, h_u_cla24_and1310_y0, h_u_cla24_and1312_y0);
  and_gate and_gate_h_u_cla24_and1313_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1313_y0);
  and_gate and_gate_h_u_cla24_and1314_y0(h_u_cla24_and1313_y0, h_u_cla24_and1312_y0, h_u_cla24_and1314_y0);
  and_gate and_gate_h_u_cla24_and1315_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1315_y0);
  and_gate and_gate_h_u_cla24_and1316_y0(h_u_cla24_and1315_y0, h_u_cla24_and1314_y0, h_u_cla24_and1316_y0);
  and_gate and_gate_h_u_cla24_and1317_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1317_y0);
  and_gate and_gate_h_u_cla24_and1318_y0(h_u_cla24_and1317_y0, h_u_cla24_and1316_y0, h_u_cla24_and1318_y0);
  and_gate and_gate_h_u_cla24_and1319_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1319_y0);
  and_gate and_gate_h_u_cla24_and1320_y0(h_u_cla24_and1319_y0, h_u_cla24_and1318_y0, h_u_cla24_and1320_y0);
  and_gate and_gate_h_u_cla24_and1321_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1321_y0);
  and_gate and_gate_h_u_cla24_and1322_y0(h_u_cla24_and1321_y0, h_u_cla24_and1320_y0, h_u_cla24_and1322_y0);
  and_gate and_gate_h_u_cla24_and1323_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1323_y0);
  and_gate and_gate_h_u_cla24_and1324_y0(h_u_cla24_and1323_y0, h_u_cla24_and1322_y0, h_u_cla24_and1324_y0);
  and_gate and_gate_h_u_cla24_and1325_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1325_y0);
  and_gate and_gate_h_u_cla24_and1326_y0(h_u_cla24_and1325_y0, h_u_cla24_and1324_y0, h_u_cla24_and1326_y0);
  and_gate and_gate_h_u_cla24_and1327_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1327_y0);
  and_gate and_gate_h_u_cla24_and1328_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1328_y0);
  and_gate and_gate_h_u_cla24_and1329_y0(h_u_cla24_and1328_y0, h_u_cla24_and1327_y0, h_u_cla24_and1329_y0);
  and_gate and_gate_h_u_cla24_and1330_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1330_y0);
  and_gate and_gate_h_u_cla24_and1331_y0(h_u_cla24_and1330_y0, h_u_cla24_and1329_y0, h_u_cla24_and1331_y0);
  and_gate and_gate_h_u_cla24_and1332_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1332_y0);
  and_gate and_gate_h_u_cla24_and1333_y0(h_u_cla24_and1332_y0, h_u_cla24_and1331_y0, h_u_cla24_and1333_y0);
  and_gate and_gate_h_u_cla24_and1334_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1334_y0);
  and_gate and_gate_h_u_cla24_and1335_y0(h_u_cla24_and1334_y0, h_u_cla24_and1333_y0, h_u_cla24_and1335_y0);
  and_gate and_gate_h_u_cla24_and1336_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1336_y0);
  and_gate and_gate_h_u_cla24_and1337_y0(h_u_cla24_and1336_y0, h_u_cla24_and1335_y0, h_u_cla24_and1337_y0);
  and_gate and_gate_h_u_cla24_and1338_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1338_y0);
  and_gate and_gate_h_u_cla24_and1339_y0(h_u_cla24_and1338_y0, h_u_cla24_and1337_y0, h_u_cla24_and1339_y0);
  and_gate and_gate_h_u_cla24_and1340_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1340_y0);
  and_gate and_gate_h_u_cla24_and1341_y0(h_u_cla24_and1340_y0, h_u_cla24_and1339_y0, h_u_cla24_and1341_y0);
  and_gate and_gate_h_u_cla24_and1342_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1342_y0);
  and_gate and_gate_h_u_cla24_and1343_y0(h_u_cla24_and1342_y0, h_u_cla24_and1341_y0, h_u_cla24_and1343_y0);
  and_gate and_gate_h_u_cla24_and1344_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1344_y0);
  and_gate and_gate_h_u_cla24_and1345_y0(h_u_cla24_and1344_y0, h_u_cla24_and1343_y0, h_u_cla24_and1345_y0);
  and_gate and_gate_h_u_cla24_and1346_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1346_y0);
  and_gate and_gate_h_u_cla24_and1347_y0(h_u_cla24_and1346_y0, h_u_cla24_and1345_y0, h_u_cla24_and1347_y0);
  and_gate and_gate_h_u_cla24_and1348_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1348_y0);
  and_gate and_gate_h_u_cla24_and1349_y0(h_u_cla24_and1348_y0, h_u_cla24_and1347_y0, h_u_cla24_and1349_y0);
  and_gate and_gate_h_u_cla24_and1350_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1350_y0);
  and_gate and_gate_h_u_cla24_and1351_y0(h_u_cla24_and1350_y0, h_u_cla24_and1349_y0, h_u_cla24_and1351_y0);
  and_gate and_gate_h_u_cla24_and1352_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1352_y0);
  and_gate and_gate_h_u_cla24_and1353_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1353_y0);
  and_gate and_gate_h_u_cla24_and1354_y0(h_u_cla24_and1353_y0, h_u_cla24_and1352_y0, h_u_cla24_and1354_y0);
  and_gate and_gate_h_u_cla24_and1355_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1355_y0);
  and_gate and_gate_h_u_cla24_and1356_y0(h_u_cla24_and1355_y0, h_u_cla24_and1354_y0, h_u_cla24_and1356_y0);
  and_gate and_gate_h_u_cla24_and1357_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1357_y0);
  and_gate and_gate_h_u_cla24_and1358_y0(h_u_cla24_and1357_y0, h_u_cla24_and1356_y0, h_u_cla24_and1358_y0);
  and_gate and_gate_h_u_cla24_and1359_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1359_y0);
  and_gate and_gate_h_u_cla24_and1360_y0(h_u_cla24_and1359_y0, h_u_cla24_and1358_y0, h_u_cla24_and1360_y0);
  and_gate and_gate_h_u_cla24_and1361_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1361_y0);
  and_gate and_gate_h_u_cla24_and1362_y0(h_u_cla24_and1361_y0, h_u_cla24_and1360_y0, h_u_cla24_and1362_y0);
  and_gate and_gate_h_u_cla24_and1363_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1363_y0);
  and_gate and_gate_h_u_cla24_and1364_y0(h_u_cla24_and1363_y0, h_u_cla24_and1362_y0, h_u_cla24_and1364_y0);
  and_gate and_gate_h_u_cla24_and1365_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1365_y0);
  and_gate and_gate_h_u_cla24_and1366_y0(h_u_cla24_and1365_y0, h_u_cla24_and1364_y0, h_u_cla24_and1366_y0);
  and_gate and_gate_h_u_cla24_and1367_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1367_y0);
  and_gate and_gate_h_u_cla24_and1368_y0(h_u_cla24_and1367_y0, h_u_cla24_and1366_y0, h_u_cla24_and1368_y0);
  and_gate and_gate_h_u_cla24_and1369_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1369_y0);
  and_gate and_gate_h_u_cla24_and1370_y0(h_u_cla24_and1369_y0, h_u_cla24_and1368_y0, h_u_cla24_and1370_y0);
  and_gate and_gate_h_u_cla24_and1371_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1371_y0);
  and_gate and_gate_h_u_cla24_and1372_y0(h_u_cla24_and1371_y0, h_u_cla24_and1370_y0, h_u_cla24_and1372_y0);
  and_gate and_gate_h_u_cla24_and1373_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1373_y0);
  and_gate and_gate_h_u_cla24_and1374_y0(h_u_cla24_and1373_y0, h_u_cla24_and1372_y0, h_u_cla24_and1374_y0);
  and_gate and_gate_h_u_cla24_and1375_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1375_y0);
  and_gate and_gate_h_u_cla24_and1376_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1376_y0);
  and_gate and_gate_h_u_cla24_and1377_y0(h_u_cla24_and1376_y0, h_u_cla24_and1375_y0, h_u_cla24_and1377_y0);
  and_gate and_gate_h_u_cla24_and1378_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1378_y0);
  and_gate and_gate_h_u_cla24_and1379_y0(h_u_cla24_and1378_y0, h_u_cla24_and1377_y0, h_u_cla24_and1379_y0);
  and_gate and_gate_h_u_cla24_and1380_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1380_y0);
  and_gate and_gate_h_u_cla24_and1381_y0(h_u_cla24_and1380_y0, h_u_cla24_and1379_y0, h_u_cla24_and1381_y0);
  and_gate and_gate_h_u_cla24_and1382_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1382_y0);
  and_gate and_gate_h_u_cla24_and1383_y0(h_u_cla24_and1382_y0, h_u_cla24_and1381_y0, h_u_cla24_and1383_y0);
  and_gate and_gate_h_u_cla24_and1384_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1384_y0);
  and_gate and_gate_h_u_cla24_and1385_y0(h_u_cla24_and1384_y0, h_u_cla24_and1383_y0, h_u_cla24_and1385_y0);
  and_gate and_gate_h_u_cla24_and1386_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1386_y0);
  and_gate and_gate_h_u_cla24_and1387_y0(h_u_cla24_and1386_y0, h_u_cla24_and1385_y0, h_u_cla24_and1387_y0);
  and_gate and_gate_h_u_cla24_and1388_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1388_y0);
  and_gate and_gate_h_u_cla24_and1389_y0(h_u_cla24_and1388_y0, h_u_cla24_and1387_y0, h_u_cla24_and1389_y0);
  and_gate and_gate_h_u_cla24_and1390_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1390_y0);
  and_gate and_gate_h_u_cla24_and1391_y0(h_u_cla24_and1390_y0, h_u_cla24_and1389_y0, h_u_cla24_and1391_y0);
  and_gate and_gate_h_u_cla24_and1392_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1392_y0);
  and_gate and_gate_h_u_cla24_and1393_y0(h_u_cla24_and1392_y0, h_u_cla24_and1391_y0, h_u_cla24_and1393_y0);
  and_gate and_gate_h_u_cla24_and1394_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1394_y0);
  and_gate and_gate_h_u_cla24_and1395_y0(h_u_cla24_and1394_y0, h_u_cla24_and1393_y0, h_u_cla24_and1395_y0);
  and_gate and_gate_h_u_cla24_and1396_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1396_y0);
  and_gate and_gate_h_u_cla24_and1397_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1397_y0);
  and_gate and_gate_h_u_cla24_and1398_y0(h_u_cla24_and1397_y0, h_u_cla24_and1396_y0, h_u_cla24_and1398_y0);
  and_gate and_gate_h_u_cla24_and1399_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1399_y0);
  and_gate and_gate_h_u_cla24_and1400_y0(h_u_cla24_and1399_y0, h_u_cla24_and1398_y0, h_u_cla24_and1400_y0);
  and_gate and_gate_h_u_cla24_and1401_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1401_y0);
  and_gate and_gate_h_u_cla24_and1402_y0(h_u_cla24_and1401_y0, h_u_cla24_and1400_y0, h_u_cla24_and1402_y0);
  and_gate and_gate_h_u_cla24_and1403_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1403_y0);
  and_gate and_gate_h_u_cla24_and1404_y0(h_u_cla24_and1403_y0, h_u_cla24_and1402_y0, h_u_cla24_and1404_y0);
  and_gate and_gate_h_u_cla24_and1405_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1405_y0);
  and_gate and_gate_h_u_cla24_and1406_y0(h_u_cla24_and1405_y0, h_u_cla24_and1404_y0, h_u_cla24_and1406_y0);
  and_gate and_gate_h_u_cla24_and1407_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1407_y0);
  and_gate and_gate_h_u_cla24_and1408_y0(h_u_cla24_and1407_y0, h_u_cla24_and1406_y0, h_u_cla24_and1408_y0);
  and_gate and_gate_h_u_cla24_and1409_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1409_y0);
  and_gate and_gate_h_u_cla24_and1410_y0(h_u_cla24_and1409_y0, h_u_cla24_and1408_y0, h_u_cla24_and1410_y0);
  and_gate and_gate_h_u_cla24_and1411_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1411_y0);
  and_gate and_gate_h_u_cla24_and1412_y0(h_u_cla24_and1411_y0, h_u_cla24_and1410_y0, h_u_cla24_and1412_y0);
  and_gate and_gate_h_u_cla24_and1413_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1413_y0);
  and_gate and_gate_h_u_cla24_and1414_y0(h_u_cla24_and1413_y0, h_u_cla24_and1412_y0, h_u_cla24_and1414_y0);
  and_gate and_gate_h_u_cla24_and1415_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1415_y0);
  and_gate and_gate_h_u_cla24_and1416_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1416_y0);
  and_gate and_gate_h_u_cla24_and1417_y0(h_u_cla24_and1416_y0, h_u_cla24_and1415_y0, h_u_cla24_and1417_y0);
  and_gate and_gate_h_u_cla24_and1418_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1418_y0);
  and_gate and_gate_h_u_cla24_and1419_y0(h_u_cla24_and1418_y0, h_u_cla24_and1417_y0, h_u_cla24_and1419_y0);
  and_gate and_gate_h_u_cla24_and1420_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1420_y0);
  and_gate and_gate_h_u_cla24_and1421_y0(h_u_cla24_and1420_y0, h_u_cla24_and1419_y0, h_u_cla24_and1421_y0);
  and_gate and_gate_h_u_cla24_and1422_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1422_y0);
  and_gate and_gate_h_u_cla24_and1423_y0(h_u_cla24_and1422_y0, h_u_cla24_and1421_y0, h_u_cla24_and1423_y0);
  and_gate and_gate_h_u_cla24_and1424_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1424_y0);
  and_gate and_gate_h_u_cla24_and1425_y0(h_u_cla24_and1424_y0, h_u_cla24_and1423_y0, h_u_cla24_and1425_y0);
  and_gate and_gate_h_u_cla24_and1426_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1426_y0);
  and_gate and_gate_h_u_cla24_and1427_y0(h_u_cla24_and1426_y0, h_u_cla24_and1425_y0, h_u_cla24_and1427_y0);
  and_gate and_gate_h_u_cla24_and1428_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1428_y0);
  and_gate and_gate_h_u_cla24_and1429_y0(h_u_cla24_and1428_y0, h_u_cla24_and1427_y0, h_u_cla24_and1429_y0);
  and_gate and_gate_h_u_cla24_and1430_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1430_y0);
  and_gate and_gate_h_u_cla24_and1431_y0(h_u_cla24_and1430_y0, h_u_cla24_and1429_y0, h_u_cla24_and1431_y0);
  and_gate and_gate_h_u_cla24_and1432_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1432_y0);
  and_gate and_gate_h_u_cla24_and1433_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1433_y0);
  and_gate and_gate_h_u_cla24_and1434_y0(h_u_cla24_and1433_y0, h_u_cla24_and1432_y0, h_u_cla24_and1434_y0);
  and_gate and_gate_h_u_cla24_and1435_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1435_y0);
  and_gate and_gate_h_u_cla24_and1436_y0(h_u_cla24_and1435_y0, h_u_cla24_and1434_y0, h_u_cla24_and1436_y0);
  and_gate and_gate_h_u_cla24_and1437_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1437_y0);
  and_gate and_gate_h_u_cla24_and1438_y0(h_u_cla24_and1437_y0, h_u_cla24_and1436_y0, h_u_cla24_and1438_y0);
  and_gate and_gate_h_u_cla24_and1439_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1439_y0);
  and_gate and_gate_h_u_cla24_and1440_y0(h_u_cla24_and1439_y0, h_u_cla24_and1438_y0, h_u_cla24_and1440_y0);
  and_gate and_gate_h_u_cla24_and1441_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1441_y0);
  and_gate and_gate_h_u_cla24_and1442_y0(h_u_cla24_and1441_y0, h_u_cla24_and1440_y0, h_u_cla24_and1442_y0);
  and_gate and_gate_h_u_cla24_and1443_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1443_y0);
  and_gate and_gate_h_u_cla24_and1444_y0(h_u_cla24_and1443_y0, h_u_cla24_and1442_y0, h_u_cla24_and1444_y0);
  and_gate and_gate_h_u_cla24_and1445_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1445_y0);
  and_gate and_gate_h_u_cla24_and1446_y0(h_u_cla24_and1445_y0, h_u_cla24_and1444_y0, h_u_cla24_and1446_y0);
  and_gate and_gate_h_u_cla24_and1447_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1447_y0);
  and_gate and_gate_h_u_cla24_and1448_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1448_y0);
  and_gate and_gate_h_u_cla24_and1449_y0(h_u_cla24_and1448_y0, h_u_cla24_and1447_y0, h_u_cla24_and1449_y0);
  and_gate and_gate_h_u_cla24_and1450_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1450_y0);
  and_gate and_gate_h_u_cla24_and1451_y0(h_u_cla24_and1450_y0, h_u_cla24_and1449_y0, h_u_cla24_and1451_y0);
  and_gate and_gate_h_u_cla24_and1452_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1452_y0);
  and_gate and_gate_h_u_cla24_and1453_y0(h_u_cla24_and1452_y0, h_u_cla24_and1451_y0, h_u_cla24_and1453_y0);
  and_gate and_gate_h_u_cla24_and1454_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1454_y0);
  and_gate and_gate_h_u_cla24_and1455_y0(h_u_cla24_and1454_y0, h_u_cla24_and1453_y0, h_u_cla24_and1455_y0);
  and_gate and_gate_h_u_cla24_and1456_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1456_y0);
  and_gate and_gate_h_u_cla24_and1457_y0(h_u_cla24_and1456_y0, h_u_cla24_and1455_y0, h_u_cla24_and1457_y0);
  and_gate and_gate_h_u_cla24_and1458_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1458_y0);
  and_gate and_gate_h_u_cla24_and1459_y0(h_u_cla24_and1458_y0, h_u_cla24_and1457_y0, h_u_cla24_and1459_y0);
  and_gate and_gate_h_u_cla24_and1460_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1460_y0);
  and_gate and_gate_h_u_cla24_and1461_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1461_y0);
  and_gate and_gate_h_u_cla24_and1462_y0(h_u_cla24_and1461_y0, h_u_cla24_and1460_y0, h_u_cla24_and1462_y0);
  and_gate and_gate_h_u_cla24_and1463_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1463_y0);
  and_gate and_gate_h_u_cla24_and1464_y0(h_u_cla24_and1463_y0, h_u_cla24_and1462_y0, h_u_cla24_and1464_y0);
  and_gate and_gate_h_u_cla24_and1465_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1465_y0);
  and_gate and_gate_h_u_cla24_and1466_y0(h_u_cla24_and1465_y0, h_u_cla24_and1464_y0, h_u_cla24_and1466_y0);
  and_gate and_gate_h_u_cla24_and1467_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1467_y0);
  and_gate and_gate_h_u_cla24_and1468_y0(h_u_cla24_and1467_y0, h_u_cla24_and1466_y0, h_u_cla24_and1468_y0);
  and_gate and_gate_h_u_cla24_and1469_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1469_y0);
  and_gate and_gate_h_u_cla24_and1470_y0(h_u_cla24_and1469_y0, h_u_cla24_and1468_y0, h_u_cla24_and1470_y0);
  and_gate and_gate_h_u_cla24_and1471_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1471_y0);
  and_gate and_gate_h_u_cla24_and1472_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1472_y0);
  and_gate and_gate_h_u_cla24_and1473_y0(h_u_cla24_and1472_y0, h_u_cla24_and1471_y0, h_u_cla24_and1473_y0);
  and_gate and_gate_h_u_cla24_and1474_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1474_y0);
  and_gate and_gate_h_u_cla24_and1475_y0(h_u_cla24_and1474_y0, h_u_cla24_and1473_y0, h_u_cla24_and1475_y0);
  and_gate and_gate_h_u_cla24_and1476_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1476_y0);
  and_gate and_gate_h_u_cla24_and1477_y0(h_u_cla24_and1476_y0, h_u_cla24_and1475_y0, h_u_cla24_and1477_y0);
  and_gate and_gate_h_u_cla24_and1478_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1478_y0);
  and_gate and_gate_h_u_cla24_and1479_y0(h_u_cla24_and1478_y0, h_u_cla24_and1477_y0, h_u_cla24_and1479_y0);
  and_gate and_gate_h_u_cla24_and1480_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1480_y0);
  and_gate and_gate_h_u_cla24_and1481_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1481_y0);
  and_gate and_gate_h_u_cla24_and1482_y0(h_u_cla24_and1481_y0, h_u_cla24_and1480_y0, h_u_cla24_and1482_y0);
  and_gate and_gate_h_u_cla24_and1483_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1483_y0);
  and_gate and_gate_h_u_cla24_and1484_y0(h_u_cla24_and1483_y0, h_u_cla24_and1482_y0, h_u_cla24_and1484_y0);
  and_gate and_gate_h_u_cla24_and1485_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1485_y0);
  and_gate and_gate_h_u_cla24_and1486_y0(h_u_cla24_and1485_y0, h_u_cla24_and1484_y0, h_u_cla24_and1486_y0);
  and_gate and_gate_h_u_cla24_and1487_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1487_y0);
  and_gate and_gate_h_u_cla24_and1488_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1488_y0);
  and_gate and_gate_h_u_cla24_and1489_y0(h_u_cla24_and1488_y0, h_u_cla24_and1487_y0, h_u_cla24_and1489_y0);
  and_gate and_gate_h_u_cla24_and1490_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1490_y0);
  and_gate and_gate_h_u_cla24_and1491_y0(h_u_cla24_and1490_y0, h_u_cla24_and1489_y0, h_u_cla24_and1491_y0);
  and_gate and_gate_h_u_cla24_and1492_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and1492_y0);
  and_gate and_gate_h_u_cla24_and1493_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and1493_y0);
  and_gate and_gate_h_u_cla24_and1494_y0(h_u_cla24_and1493_y0, h_u_cla24_and1492_y0, h_u_cla24_and1494_y0);
  and_gate and_gate_h_u_cla24_and1495_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and1495_y0);
  or_gate or_gate_h_u_cla24_or120_y0(h_u_cla24_and1495_y0, h_u_cla24_and1270_y0, h_u_cla24_or120_y0);
  or_gate or_gate_h_u_cla24_or121_y0(h_u_cla24_or120_y0, h_u_cla24_and1299_y0, h_u_cla24_or121_y0);
  or_gate or_gate_h_u_cla24_or122_y0(h_u_cla24_or121_y0, h_u_cla24_and1326_y0, h_u_cla24_or122_y0);
  or_gate or_gate_h_u_cla24_or123_y0(h_u_cla24_or122_y0, h_u_cla24_and1351_y0, h_u_cla24_or123_y0);
  or_gate or_gate_h_u_cla24_or124_y0(h_u_cla24_or123_y0, h_u_cla24_and1374_y0, h_u_cla24_or124_y0);
  or_gate or_gate_h_u_cla24_or125_y0(h_u_cla24_or124_y0, h_u_cla24_and1395_y0, h_u_cla24_or125_y0);
  or_gate or_gate_h_u_cla24_or126_y0(h_u_cla24_or125_y0, h_u_cla24_and1414_y0, h_u_cla24_or126_y0);
  or_gate or_gate_h_u_cla24_or127_y0(h_u_cla24_or126_y0, h_u_cla24_and1431_y0, h_u_cla24_or127_y0);
  or_gate or_gate_h_u_cla24_or128_y0(h_u_cla24_or127_y0, h_u_cla24_and1446_y0, h_u_cla24_or128_y0);
  or_gate or_gate_h_u_cla24_or129_y0(h_u_cla24_or128_y0, h_u_cla24_and1459_y0, h_u_cla24_or129_y0);
  or_gate or_gate_h_u_cla24_or130_y0(h_u_cla24_or129_y0, h_u_cla24_and1470_y0, h_u_cla24_or130_y0);
  or_gate or_gate_h_u_cla24_or131_y0(h_u_cla24_or130_y0, h_u_cla24_and1479_y0, h_u_cla24_or131_y0);
  or_gate or_gate_h_u_cla24_or132_y0(h_u_cla24_or131_y0, h_u_cla24_and1486_y0, h_u_cla24_or132_y0);
  or_gate or_gate_h_u_cla24_or133_y0(h_u_cla24_or132_y0, h_u_cla24_and1491_y0, h_u_cla24_or133_y0);
  or_gate or_gate_h_u_cla24_or134_y0(h_u_cla24_or133_y0, h_u_cla24_and1494_y0, h_u_cla24_or134_y0);
  or_gate or_gate_h_u_cla24_or135_y0(h_u_cla24_pg_logic15_y1, h_u_cla24_or134_y0, h_u_cla24_or135_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic16_y0(a_16, b_16, h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_pg_logic16_y2);
  xor_gate xor_gate_h_u_cla24_xor16_y0(h_u_cla24_pg_logic16_y2, h_u_cla24_or135_y0, h_u_cla24_xor16_y0);
  and_gate and_gate_h_u_cla24_and1496_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and1496_y0);
  and_gate and_gate_h_u_cla24_and1497_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and1497_y0);
  and_gate and_gate_h_u_cla24_and1498_y0(h_u_cla24_and1497_y0, h_u_cla24_and1496_y0, h_u_cla24_and1498_y0);
  and_gate and_gate_h_u_cla24_and1499_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and1499_y0);
  and_gate and_gate_h_u_cla24_and1500_y0(h_u_cla24_and1499_y0, h_u_cla24_and1498_y0, h_u_cla24_and1500_y0);
  and_gate and_gate_h_u_cla24_and1501_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and1501_y0);
  and_gate and_gate_h_u_cla24_and1502_y0(h_u_cla24_and1501_y0, h_u_cla24_and1500_y0, h_u_cla24_and1502_y0);
  and_gate and_gate_h_u_cla24_and1503_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and1503_y0);
  and_gate and_gate_h_u_cla24_and1504_y0(h_u_cla24_and1503_y0, h_u_cla24_and1502_y0, h_u_cla24_and1504_y0);
  and_gate and_gate_h_u_cla24_and1505_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and1505_y0);
  and_gate and_gate_h_u_cla24_and1506_y0(h_u_cla24_and1505_y0, h_u_cla24_and1504_y0, h_u_cla24_and1506_y0);
  and_gate and_gate_h_u_cla24_and1507_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and1507_y0);
  and_gate and_gate_h_u_cla24_and1508_y0(h_u_cla24_and1507_y0, h_u_cla24_and1506_y0, h_u_cla24_and1508_y0);
  and_gate and_gate_h_u_cla24_and1509_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and1509_y0);
  and_gate and_gate_h_u_cla24_and1510_y0(h_u_cla24_and1509_y0, h_u_cla24_and1508_y0, h_u_cla24_and1510_y0);
  and_gate and_gate_h_u_cla24_and1511_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and1511_y0);
  and_gate and_gate_h_u_cla24_and1512_y0(h_u_cla24_and1511_y0, h_u_cla24_and1510_y0, h_u_cla24_and1512_y0);
  and_gate and_gate_h_u_cla24_and1513_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and1513_y0);
  and_gate and_gate_h_u_cla24_and1514_y0(h_u_cla24_and1513_y0, h_u_cla24_and1512_y0, h_u_cla24_and1514_y0);
  and_gate and_gate_h_u_cla24_and1515_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and1515_y0);
  and_gate and_gate_h_u_cla24_and1516_y0(h_u_cla24_and1515_y0, h_u_cla24_and1514_y0, h_u_cla24_and1516_y0);
  and_gate and_gate_h_u_cla24_and1517_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and1517_y0);
  and_gate and_gate_h_u_cla24_and1518_y0(h_u_cla24_and1517_y0, h_u_cla24_and1516_y0, h_u_cla24_and1518_y0);
  and_gate and_gate_h_u_cla24_and1519_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and1519_y0);
  and_gate and_gate_h_u_cla24_and1520_y0(h_u_cla24_and1519_y0, h_u_cla24_and1518_y0, h_u_cla24_and1520_y0);
  and_gate and_gate_h_u_cla24_and1521_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and1521_y0);
  and_gate and_gate_h_u_cla24_and1522_y0(h_u_cla24_and1521_y0, h_u_cla24_and1520_y0, h_u_cla24_and1522_y0);
  and_gate and_gate_h_u_cla24_and1523_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and1523_y0);
  and_gate and_gate_h_u_cla24_and1524_y0(h_u_cla24_and1523_y0, h_u_cla24_and1522_y0, h_u_cla24_and1524_y0);
  and_gate and_gate_h_u_cla24_and1525_y0(h_u_cla24_pg_logic15_y0, constant_wire_0, h_u_cla24_and1525_y0);
  and_gate and_gate_h_u_cla24_and1526_y0(h_u_cla24_and1525_y0, h_u_cla24_and1524_y0, h_u_cla24_and1526_y0);
  and_gate and_gate_h_u_cla24_and1527_y0(h_u_cla24_pg_logic16_y0, constant_wire_0, h_u_cla24_and1527_y0);
  and_gate and_gate_h_u_cla24_and1528_y0(h_u_cla24_and1527_y0, h_u_cla24_and1526_y0, h_u_cla24_and1528_y0);
  and_gate and_gate_h_u_cla24_and1529_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1529_y0);
  and_gate and_gate_h_u_cla24_and1530_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1530_y0);
  and_gate and_gate_h_u_cla24_and1531_y0(h_u_cla24_and1530_y0, h_u_cla24_and1529_y0, h_u_cla24_and1531_y0);
  and_gate and_gate_h_u_cla24_and1532_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1532_y0);
  and_gate and_gate_h_u_cla24_and1533_y0(h_u_cla24_and1532_y0, h_u_cla24_and1531_y0, h_u_cla24_and1533_y0);
  and_gate and_gate_h_u_cla24_and1534_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1534_y0);
  and_gate and_gate_h_u_cla24_and1535_y0(h_u_cla24_and1534_y0, h_u_cla24_and1533_y0, h_u_cla24_and1535_y0);
  and_gate and_gate_h_u_cla24_and1536_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1536_y0);
  and_gate and_gate_h_u_cla24_and1537_y0(h_u_cla24_and1536_y0, h_u_cla24_and1535_y0, h_u_cla24_and1537_y0);
  and_gate and_gate_h_u_cla24_and1538_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1538_y0);
  and_gate and_gate_h_u_cla24_and1539_y0(h_u_cla24_and1538_y0, h_u_cla24_and1537_y0, h_u_cla24_and1539_y0);
  and_gate and_gate_h_u_cla24_and1540_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1540_y0);
  and_gate and_gate_h_u_cla24_and1541_y0(h_u_cla24_and1540_y0, h_u_cla24_and1539_y0, h_u_cla24_and1541_y0);
  and_gate and_gate_h_u_cla24_and1542_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1542_y0);
  and_gate and_gate_h_u_cla24_and1543_y0(h_u_cla24_and1542_y0, h_u_cla24_and1541_y0, h_u_cla24_and1543_y0);
  and_gate and_gate_h_u_cla24_and1544_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1544_y0);
  and_gate and_gate_h_u_cla24_and1545_y0(h_u_cla24_and1544_y0, h_u_cla24_and1543_y0, h_u_cla24_and1545_y0);
  and_gate and_gate_h_u_cla24_and1546_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1546_y0);
  and_gate and_gate_h_u_cla24_and1547_y0(h_u_cla24_and1546_y0, h_u_cla24_and1545_y0, h_u_cla24_and1547_y0);
  and_gate and_gate_h_u_cla24_and1548_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1548_y0);
  and_gate and_gate_h_u_cla24_and1549_y0(h_u_cla24_and1548_y0, h_u_cla24_and1547_y0, h_u_cla24_and1549_y0);
  and_gate and_gate_h_u_cla24_and1550_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1550_y0);
  and_gate and_gate_h_u_cla24_and1551_y0(h_u_cla24_and1550_y0, h_u_cla24_and1549_y0, h_u_cla24_and1551_y0);
  and_gate and_gate_h_u_cla24_and1552_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1552_y0);
  and_gate and_gate_h_u_cla24_and1553_y0(h_u_cla24_and1552_y0, h_u_cla24_and1551_y0, h_u_cla24_and1553_y0);
  and_gate and_gate_h_u_cla24_and1554_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1554_y0);
  and_gate and_gate_h_u_cla24_and1555_y0(h_u_cla24_and1554_y0, h_u_cla24_and1553_y0, h_u_cla24_and1555_y0);
  and_gate and_gate_h_u_cla24_and1556_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1556_y0);
  and_gate and_gate_h_u_cla24_and1557_y0(h_u_cla24_and1556_y0, h_u_cla24_and1555_y0, h_u_cla24_and1557_y0);
  and_gate and_gate_h_u_cla24_and1558_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1558_y0);
  and_gate and_gate_h_u_cla24_and1559_y0(h_u_cla24_and1558_y0, h_u_cla24_and1557_y0, h_u_cla24_and1559_y0);
  and_gate and_gate_h_u_cla24_and1560_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1560_y0);
  and_gate and_gate_h_u_cla24_and1561_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1561_y0);
  and_gate and_gate_h_u_cla24_and1562_y0(h_u_cla24_and1561_y0, h_u_cla24_and1560_y0, h_u_cla24_and1562_y0);
  and_gate and_gate_h_u_cla24_and1563_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1563_y0);
  and_gate and_gate_h_u_cla24_and1564_y0(h_u_cla24_and1563_y0, h_u_cla24_and1562_y0, h_u_cla24_and1564_y0);
  and_gate and_gate_h_u_cla24_and1565_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1565_y0);
  and_gate and_gate_h_u_cla24_and1566_y0(h_u_cla24_and1565_y0, h_u_cla24_and1564_y0, h_u_cla24_and1566_y0);
  and_gate and_gate_h_u_cla24_and1567_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1567_y0);
  and_gate and_gate_h_u_cla24_and1568_y0(h_u_cla24_and1567_y0, h_u_cla24_and1566_y0, h_u_cla24_and1568_y0);
  and_gate and_gate_h_u_cla24_and1569_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1569_y0);
  and_gate and_gate_h_u_cla24_and1570_y0(h_u_cla24_and1569_y0, h_u_cla24_and1568_y0, h_u_cla24_and1570_y0);
  and_gate and_gate_h_u_cla24_and1571_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1571_y0);
  and_gate and_gate_h_u_cla24_and1572_y0(h_u_cla24_and1571_y0, h_u_cla24_and1570_y0, h_u_cla24_and1572_y0);
  and_gate and_gate_h_u_cla24_and1573_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1573_y0);
  and_gate and_gate_h_u_cla24_and1574_y0(h_u_cla24_and1573_y0, h_u_cla24_and1572_y0, h_u_cla24_and1574_y0);
  and_gate and_gate_h_u_cla24_and1575_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1575_y0);
  and_gate and_gate_h_u_cla24_and1576_y0(h_u_cla24_and1575_y0, h_u_cla24_and1574_y0, h_u_cla24_and1576_y0);
  and_gate and_gate_h_u_cla24_and1577_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1577_y0);
  and_gate and_gate_h_u_cla24_and1578_y0(h_u_cla24_and1577_y0, h_u_cla24_and1576_y0, h_u_cla24_and1578_y0);
  and_gate and_gate_h_u_cla24_and1579_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1579_y0);
  and_gate and_gate_h_u_cla24_and1580_y0(h_u_cla24_and1579_y0, h_u_cla24_and1578_y0, h_u_cla24_and1580_y0);
  and_gate and_gate_h_u_cla24_and1581_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1581_y0);
  and_gate and_gate_h_u_cla24_and1582_y0(h_u_cla24_and1581_y0, h_u_cla24_and1580_y0, h_u_cla24_and1582_y0);
  and_gate and_gate_h_u_cla24_and1583_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1583_y0);
  and_gate and_gate_h_u_cla24_and1584_y0(h_u_cla24_and1583_y0, h_u_cla24_and1582_y0, h_u_cla24_and1584_y0);
  and_gate and_gate_h_u_cla24_and1585_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1585_y0);
  and_gate and_gate_h_u_cla24_and1586_y0(h_u_cla24_and1585_y0, h_u_cla24_and1584_y0, h_u_cla24_and1586_y0);
  and_gate and_gate_h_u_cla24_and1587_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1587_y0);
  and_gate and_gate_h_u_cla24_and1588_y0(h_u_cla24_and1587_y0, h_u_cla24_and1586_y0, h_u_cla24_and1588_y0);
  and_gate and_gate_h_u_cla24_and1589_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1589_y0);
  and_gate and_gate_h_u_cla24_and1590_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1590_y0);
  and_gate and_gate_h_u_cla24_and1591_y0(h_u_cla24_and1590_y0, h_u_cla24_and1589_y0, h_u_cla24_and1591_y0);
  and_gate and_gate_h_u_cla24_and1592_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1592_y0);
  and_gate and_gate_h_u_cla24_and1593_y0(h_u_cla24_and1592_y0, h_u_cla24_and1591_y0, h_u_cla24_and1593_y0);
  and_gate and_gate_h_u_cla24_and1594_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1594_y0);
  and_gate and_gate_h_u_cla24_and1595_y0(h_u_cla24_and1594_y0, h_u_cla24_and1593_y0, h_u_cla24_and1595_y0);
  and_gate and_gate_h_u_cla24_and1596_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1596_y0);
  and_gate and_gate_h_u_cla24_and1597_y0(h_u_cla24_and1596_y0, h_u_cla24_and1595_y0, h_u_cla24_and1597_y0);
  and_gate and_gate_h_u_cla24_and1598_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1598_y0);
  and_gate and_gate_h_u_cla24_and1599_y0(h_u_cla24_and1598_y0, h_u_cla24_and1597_y0, h_u_cla24_and1599_y0);
  and_gate and_gate_h_u_cla24_and1600_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1600_y0);
  and_gate and_gate_h_u_cla24_and1601_y0(h_u_cla24_and1600_y0, h_u_cla24_and1599_y0, h_u_cla24_and1601_y0);
  and_gate and_gate_h_u_cla24_and1602_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1602_y0);
  and_gate and_gate_h_u_cla24_and1603_y0(h_u_cla24_and1602_y0, h_u_cla24_and1601_y0, h_u_cla24_and1603_y0);
  and_gate and_gate_h_u_cla24_and1604_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1604_y0);
  and_gate and_gate_h_u_cla24_and1605_y0(h_u_cla24_and1604_y0, h_u_cla24_and1603_y0, h_u_cla24_and1605_y0);
  and_gate and_gate_h_u_cla24_and1606_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1606_y0);
  and_gate and_gate_h_u_cla24_and1607_y0(h_u_cla24_and1606_y0, h_u_cla24_and1605_y0, h_u_cla24_and1607_y0);
  and_gate and_gate_h_u_cla24_and1608_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1608_y0);
  and_gate and_gate_h_u_cla24_and1609_y0(h_u_cla24_and1608_y0, h_u_cla24_and1607_y0, h_u_cla24_and1609_y0);
  and_gate and_gate_h_u_cla24_and1610_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1610_y0);
  and_gate and_gate_h_u_cla24_and1611_y0(h_u_cla24_and1610_y0, h_u_cla24_and1609_y0, h_u_cla24_and1611_y0);
  and_gate and_gate_h_u_cla24_and1612_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1612_y0);
  and_gate and_gate_h_u_cla24_and1613_y0(h_u_cla24_and1612_y0, h_u_cla24_and1611_y0, h_u_cla24_and1613_y0);
  and_gate and_gate_h_u_cla24_and1614_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1614_y0);
  and_gate and_gate_h_u_cla24_and1615_y0(h_u_cla24_and1614_y0, h_u_cla24_and1613_y0, h_u_cla24_and1615_y0);
  and_gate and_gate_h_u_cla24_and1616_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1616_y0);
  and_gate and_gate_h_u_cla24_and1617_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1617_y0);
  and_gate and_gate_h_u_cla24_and1618_y0(h_u_cla24_and1617_y0, h_u_cla24_and1616_y0, h_u_cla24_and1618_y0);
  and_gate and_gate_h_u_cla24_and1619_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1619_y0);
  and_gate and_gate_h_u_cla24_and1620_y0(h_u_cla24_and1619_y0, h_u_cla24_and1618_y0, h_u_cla24_and1620_y0);
  and_gate and_gate_h_u_cla24_and1621_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1621_y0);
  and_gate and_gate_h_u_cla24_and1622_y0(h_u_cla24_and1621_y0, h_u_cla24_and1620_y0, h_u_cla24_and1622_y0);
  and_gate and_gate_h_u_cla24_and1623_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1623_y0);
  and_gate and_gate_h_u_cla24_and1624_y0(h_u_cla24_and1623_y0, h_u_cla24_and1622_y0, h_u_cla24_and1624_y0);
  and_gate and_gate_h_u_cla24_and1625_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1625_y0);
  and_gate and_gate_h_u_cla24_and1626_y0(h_u_cla24_and1625_y0, h_u_cla24_and1624_y0, h_u_cla24_and1626_y0);
  and_gate and_gate_h_u_cla24_and1627_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1627_y0);
  and_gate and_gate_h_u_cla24_and1628_y0(h_u_cla24_and1627_y0, h_u_cla24_and1626_y0, h_u_cla24_and1628_y0);
  and_gate and_gate_h_u_cla24_and1629_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1629_y0);
  and_gate and_gate_h_u_cla24_and1630_y0(h_u_cla24_and1629_y0, h_u_cla24_and1628_y0, h_u_cla24_and1630_y0);
  and_gate and_gate_h_u_cla24_and1631_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1631_y0);
  and_gate and_gate_h_u_cla24_and1632_y0(h_u_cla24_and1631_y0, h_u_cla24_and1630_y0, h_u_cla24_and1632_y0);
  and_gate and_gate_h_u_cla24_and1633_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1633_y0);
  and_gate and_gate_h_u_cla24_and1634_y0(h_u_cla24_and1633_y0, h_u_cla24_and1632_y0, h_u_cla24_and1634_y0);
  and_gate and_gate_h_u_cla24_and1635_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1635_y0);
  and_gate and_gate_h_u_cla24_and1636_y0(h_u_cla24_and1635_y0, h_u_cla24_and1634_y0, h_u_cla24_and1636_y0);
  and_gate and_gate_h_u_cla24_and1637_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1637_y0);
  and_gate and_gate_h_u_cla24_and1638_y0(h_u_cla24_and1637_y0, h_u_cla24_and1636_y0, h_u_cla24_and1638_y0);
  and_gate and_gate_h_u_cla24_and1639_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1639_y0);
  and_gate and_gate_h_u_cla24_and1640_y0(h_u_cla24_and1639_y0, h_u_cla24_and1638_y0, h_u_cla24_and1640_y0);
  and_gate and_gate_h_u_cla24_and1641_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1641_y0);
  and_gate and_gate_h_u_cla24_and1642_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1642_y0);
  and_gate and_gate_h_u_cla24_and1643_y0(h_u_cla24_and1642_y0, h_u_cla24_and1641_y0, h_u_cla24_and1643_y0);
  and_gate and_gate_h_u_cla24_and1644_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1644_y0);
  and_gate and_gate_h_u_cla24_and1645_y0(h_u_cla24_and1644_y0, h_u_cla24_and1643_y0, h_u_cla24_and1645_y0);
  and_gate and_gate_h_u_cla24_and1646_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1646_y0);
  and_gate and_gate_h_u_cla24_and1647_y0(h_u_cla24_and1646_y0, h_u_cla24_and1645_y0, h_u_cla24_and1647_y0);
  and_gate and_gate_h_u_cla24_and1648_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1648_y0);
  and_gate and_gate_h_u_cla24_and1649_y0(h_u_cla24_and1648_y0, h_u_cla24_and1647_y0, h_u_cla24_and1649_y0);
  and_gate and_gate_h_u_cla24_and1650_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1650_y0);
  and_gate and_gate_h_u_cla24_and1651_y0(h_u_cla24_and1650_y0, h_u_cla24_and1649_y0, h_u_cla24_and1651_y0);
  and_gate and_gate_h_u_cla24_and1652_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1652_y0);
  and_gate and_gate_h_u_cla24_and1653_y0(h_u_cla24_and1652_y0, h_u_cla24_and1651_y0, h_u_cla24_and1653_y0);
  and_gate and_gate_h_u_cla24_and1654_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1654_y0);
  and_gate and_gate_h_u_cla24_and1655_y0(h_u_cla24_and1654_y0, h_u_cla24_and1653_y0, h_u_cla24_and1655_y0);
  and_gate and_gate_h_u_cla24_and1656_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1656_y0);
  and_gate and_gate_h_u_cla24_and1657_y0(h_u_cla24_and1656_y0, h_u_cla24_and1655_y0, h_u_cla24_and1657_y0);
  and_gate and_gate_h_u_cla24_and1658_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1658_y0);
  and_gate and_gate_h_u_cla24_and1659_y0(h_u_cla24_and1658_y0, h_u_cla24_and1657_y0, h_u_cla24_and1659_y0);
  and_gate and_gate_h_u_cla24_and1660_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1660_y0);
  and_gate and_gate_h_u_cla24_and1661_y0(h_u_cla24_and1660_y0, h_u_cla24_and1659_y0, h_u_cla24_and1661_y0);
  and_gate and_gate_h_u_cla24_and1662_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1662_y0);
  and_gate and_gate_h_u_cla24_and1663_y0(h_u_cla24_and1662_y0, h_u_cla24_and1661_y0, h_u_cla24_and1663_y0);
  and_gate and_gate_h_u_cla24_and1664_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1664_y0);
  and_gate and_gate_h_u_cla24_and1665_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1665_y0);
  and_gate and_gate_h_u_cla24_and1666_y0(h_u_cla24_and1665_y0, h_u_cla24_and1664_y0, h_u_cla24_and1666_y0);
  and_gate and_gate_h_u_cla24_and1667_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1667_y0);
  and_gate and_gate_h_u_cla24_and1668_y0(h_u_cla24_and1667_y0, h_u_cla24_and1666_y0, h_u_cla24_and1668_y0);
  and_gate and_gate_h_u_cla24_and1669_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1669_y0);
  and_gate and_gate_h_u_cla24_and1670_y0(h_u_cla24_and1669_y0, h_u_cla24_and1668_y0, h_u_cla24_and1670_y0);
  and_gate and_gate_h_u_cla24_and1671_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1671_y0);
  and_gate and_gate_h_u_cla24_and1672_y0(h_u_cla24_and1671_y0, h_u_cla24_and1670_y0, h_u_cla24_and1672_y0);
  and_gate and_gate_h_u_cla24_and1673_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1673_y0);
  and_gate and_gate_h_u_cla24_and1674_y0(h_u_cla24_and1673_y0, h_u_cla24_and1672_y0, h_u_cla24_and1674_y0);
  and_gate and_gate_h_u_cla24_and1675_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1675_y0);
  and_gate and_gate_h_u_cla24_and1676_y0(h_u_cla24_and1675_y0, h_u_cla24_and1674_y0, h_u_cla24_and1676_y0);
  and_gate and_gate_h_u_cla24_and1677_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1677_y0);
  and_gate and_gate_h_u_cla24_and1678_y0(h_u_cla24_and1677_y0, h_u_cla24_and1676_y0, h_u_cla24_and1678_y0);
  and_gate and_gate_h_u_cla24_and1679_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1679_y0);
  and_gate and_gate_h_u_cla24_and1680_y0(h_u_cla24_and1679_y0, h_u_cla24_and1678_y0, h_u_cla24_and1680_y0);
  and_gate and_gate_h_u_cla24_and1681_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1681_y0);
  and_gate and_gate_h_u_cla24_and1682_y0(h_u_cla24_and1681_y0, h_u_cla24_and1680_y0, h_u_cla24_and1682_y0);
  and_gate and_gate_h_u_cla24_and1683_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1683_y0);
  and_gate and_gate_h_u_cla24_and1684_y0(h_u_cla24_and1683_y0, h_u_cla24_and1682_y0, h_u_cla24_and1684_y0);
  and_gate and_gate_h_u_cla24_and1685_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1685_y0);
  and_gate and_gate_h_u_cla24_and1686_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1686_y0);
  and_gate and_gate_h_u_cla24_and1687_y0(h_u_cla24_and1686_y0, h_u_cla24_and1685_y0, h_u_cla24_and1687_y0);
  and_gate and_gate_h_u_cla24_and1688_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1688_y0);
  and_gate and_gate_h_u_cla24_and1689_y0(h_u_cla24_and1688_y0, h_u_cla24_and1687_y0, h_u_cla24_and1689_y0);
  and_gate and_gate_h_u_cla24_and1690_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1690_y0);
  and_gate and_gate_h_u_cla24_and1691_y0(h_u_cla24_and1690_y0, h_u_cla24_and1689_y0, h_u_cla24_and1691_y0);
  and_gate and_gate_h_u_cla24_and1692_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1692_y0);
  and_gate and_gate_h_u_cla24_and1693_y0(h_u_cla24_and1692_y0, h_u_cla24_and1691_y0, h_u_cla24_and1693_y0);
  and_gate and_gate_h_u_cla24_and1694_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1694_y0);
  and_gate and_gate_h_u_cla24_and1695_y0(h_u_cla24_and1694_y0, h_u_cla24_and1693_y0, h_u_cla24_and1695_y0);
  and_gate and_gate_h_u_cla24_and1696_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1696_y0);
  and_gate and_gate_h_u_cla24_and1697_y0(h_u_cla24_and1696_y0, h_u_cla24_and1695_y0, h_u_cla24_and1697_y0);
  and_gate and_gate_h_u_cla24_and1698_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1698_y0);
  and_gate and_gate_h_u_cla24_and1699_y0(h_u_cla24_and1698_y0, h_u_cla24_and1697_y0, h_u_cla24_and1699_y0);
  and_gate and_gate_h_u_cla24_and1700_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1700_y0);
  and_gate and_gate_h_u_cla24_and1701_y0(h_u_cla24_and1700_y0, h_u_cla24_and1699_y0, h_u_cla24_and1701_y0);
  and_gate and_gate_h_u_cla24_and1702_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1702_y0);
  and_gate and_gate_h_u_cla24_and1703_y0(h_u_cla24_and1702_y0, h_u_cla24_and1701_y0, h_u_cla24_and1703_y0);
  and_gate and_gate_h_u_cla24_and1704_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1704_y0);
  and_gate and_gate_h_u_cla24_and1705_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1705_y0);
  and_gate and_gate_h_u_cla24_and1706_y0(h_u_cla24_and1705_y0, h_u_cla24_and1704_y0, h_u_cla24_and1706_y0);
  and_gate and_gate_h_u_cla24_and1707_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1707_y0);
  and_gate and_gate_h_u_cla24_and1708_y0(h_u_cla24_and1707_y0, h_u_cla24_and1706_y0, h_u_cla24_and1708_y0);
  and_gate and_gate_h_u_cla24_and1709_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1709_y0);
  and_gate and_gate_h_u_cla24_and1710_y0(h_u_cla24_and1709_y0, h_u_cla24_and1708_y0, h_u_cla24_and1710_y0);
  and_gate and_gate_h_u_cla24_and1711_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1711_y0);
  and_gate and_gate_h_u_cla24_and1712_y0(h_u_cla24_and1711_y0, h_u_cla24_and1710_y0, h_u_cla24_and1712_y0);
  and_gate and_gate_h_u_cla24_and1713_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1713_y0);
  and_gate and_gate_h_u_cla24_and1714_y0(h_u_cla24_and1713_y0, h_u_cla24_and1712_y0, h_u_cla24_and1714_y0);
  and_gate and_gate_h_u_cla24_and1715_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1715_y0);
  and_gate and_gate_h_u_cla24_and1716_y0(h_u_cla24_and1715_y0, h_u_cla24_and1714_y0, h_u_cla24_and1716_y0);
  and_gate and_gate_h_u_cla24_and1717_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1717_y0);
  and_gate and_gate_h_u_cla24_and1718_y0(h_u_cla24_and1717_y0, h_u_cla24_and1716_y0, h_u_cla24_and1718_y0);
  and_gate and_gate_h_u_cla24_and1719_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and1719_y0);
  and_gate and_gate_h_u_cla24_and1720_y0(h_u_cla24_and1719_y0, h_u_cla24_and1718_y0, h_u_cla24_and1720_y0);
  and_gate and_gate_h_u_cla24_and1721_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1721_y0);
  and_gate and_gate_h_u_cla24_and1722_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1722_y0);
  and_gate and_gate_h_u_cla24_and1723_y0(h_u_cla24_and1722_y0, h_u_cla24_and1721_y0, h_u_cla24_and1723_y0);
  and_gate and_gate_h_u_cla24_and1724_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1724_y0);
  and_gate and_gate_h_u_cla24_and1725_y0(h_u_cla24_and1724_y0, h_u_cla24_and1723_y0, h_u_cla24_and1725_y0);
  and_gate and_gate_h_u_cla24_and1726_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1726_y0);
  and_gate and_gate_h_u_cla24_and1727_y0(h_u_cla24_and1726_y0, h_u_cla24_and1725_y0, h_u_cla24_and1727_y0);
  and_gate and_gate_h_u_cla24_and1728_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1728_y0);
  and_gate and_gate_h_u_cla24_and1729_y0(h_u_cla24_and1728_y0, h_u_cla24_and1727_y0, h_u_cla24_and1729_y0);
  and_gate and_gate_h_u_cla24_and1730_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1730_y0);
  and_gate and_gate_h_u_cla24_and1731_y0(h_u_cla24_and1730_y0, h_u_cla24_and1729_y0, h_u_cla24_and1731_y0);
  and_gate and_gate_h_u_cla24_and1732_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1732_y0);
  and_gate and_gate_h_u_cla24_and1733_y0(h_u_cla24_and1732_y0, h_u_cla24_and1731_y0, h_u_cla24_and1733_y0);
  and_gate and_gate_h_u_cla24_and1734_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and1734_y0);
  and_gate and_gate_h_u_cla24_and1735_y0(h_u_cla24_and1734_y0, h_u_cla24_and1733_y0, h_u_cla24_and1735_y0);
  and_gate and_gate_h_u_cla24_and1736_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1736_y0);
  and_gate and_gate_h_u_cla24_and1737_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1737_y0);
  and_gate and_gate_h_u_cla24_and1738_y0(h_u_cla24_and1737_y0, h_u_cla24_and1736_y0, h_u_cla24_and1738_y0);
  and_gate and_gate_h_u_cla24_and1739_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1739_y0);
  and_gate and_gate_h_u_cla24_and1740_y0(h_u_cla24_and1739_y0, h_u_cla24_and1738_y0, h_u_cla24_and1740_y0);
  and_gate and_gate_h_u_cla24_and1741_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1741_y0);
  and_gate and_gate_h_u_cla24_and1742_y0(h_u_cla24_and1741_y0, h_u_cla24_and1740_y0, h_u_cla24_and1742_y0);
  and_gate and_gate_h_u_cla24_and1743_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1743_y0);
  and_gate and_gate_h_u_cla24_and1744_y0(h_u_cla24_and1743_y0, h_u_cla24_and1742_y0, h_u_cla24_and1744_y0);
  and_gate and_gate_h_u_cla24_and1745_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1745_y0);
  and_gate and_gate_h_u_cla24_and1746_y0(h_u_cla24_and1745_y0, h_u_cla24_and1744_y0, h_u_cla24_and1746_y0);
  and_gate and_gate_h_u_cla24_and1747_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and1747_y0);
  and_gate and_gate_h_u_cla24_and1748_y0(h_u_cla24_and1747_y0, h_u_cla24_and1746_y0, h_u_cla24_and1748_y0);
  and_gate and_gate_h_u_cla24_and1749_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1749_y0);
  and_gate and_gate_h_u_cla24_and1750_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1750_y0);
  and_gate and_gate_h_u_cla24_and1751_y0(h_u_cla24_and1750_y0, h_u_cla24_and1749_y0, h_u_cla24_and1751_y0);
  and_gate and_gate_h_u_cla24_and1752_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1752_y0);
  and_gate and_gate_h_u_cla24_and1753_y0(h_u_cla24_and1752_y0, h_u_cla24_and1751_y0, h_u_cla24_and1753_y0);
  and_gate and_gate_h_u_cla24_and1754_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1754_y0);
  and_gate and_gate_h_u_cla24_and1755_y0(h_u_cla24_and1754_y0, h_u_cla24_and1753_y0, h_u_cla24_and1755_y0);
  and_gate and_gate_h_u_cla24_and1756_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1756_y0);
  and_gate and_gate_h_u_cla24_and1757_y0(h_u_cla24_and1756_y0, h_u_cla24_and1755_y0, h_u_cla24_and1757_y0);
  and_gate and_gate_h_u_cla24_and1758_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and1758_y0);
  and_gate and_gate_h_u_cla24_and1759_y0(h_u_cla24_and1758_y0, h_u_cla24_and1757_y0, h_u_cla24_and1759_y0);
  and_gate and_gate_h_u_cla24_and1760_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1760_y0);
  and_gate and_gate_h_u_cla24_and1761_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1761_y0);
  and_gate and_gate_h_u_cla24_and1762_y0(h_u_cla24_and1761_y0, h_u_cla24_and1760_y0, h_u_cla24_and1762_y0);
  and_gate and_gate_h_u_cla24_and1763_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1763_y0);
  and_gate and_gate_h_u_cla24_and1764_y0(h_u_cla24_and1763_y0, h_u_cla24_and1762_y0, h_u_cla24_and1764_y0);
  and_gate and_gate_h_u_cla24_and1765_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1765_y0);
  and_gate and_gate_h_u_cla24_and1766_y0(h_u_cla24_and1765_y0, h_u_cla24_and1764_y0, h_u_cla24_and1766_y0);
  and_gate and_gate_h_u_cla24_and1767_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and1767_y0);
  and_gate and_gate_h_u_cla24_and1768_y0(h_u_cla24_and1767_y0, h_u_cla24_and1766_y0, h_u_cla24_and1768_y0);
  and_gate and_gate_h_u_cla24_and1769_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1769_y0);
  and_gate and_gate_h_u_cla24_and1770_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1770_y0);
  and_gate and_gate_h_u_cla24_and1771_y0(h_u_cla24_and1770_y0, h_u_cla24_and1769_y0, h_u_cla24_and1771_y0);
  and_gate and_gate_h_u_cla24_and1772_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1772_y0);
  and_gate and_gate_h_u_cla24_and1773_y0(h_u_cla24_and1772_y0, h_u_cla24_and1771_y0, h_u_cla24_and1773_y0);
  and_gate and_gate_h_u_cla24_and1774_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and1774_y0);
  and_gate and_gate_h_u_cla24_and1775_y0(h_u_cla24_and1774_y0, h_u_cla24_and1773_y0, h_u_cla24_and1775_y0);
  and_gate and_gate_h_u_cla24_and1776_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and1776_y0);
  and_gate and_gate_h_u_cla24_and1777_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and1777_y0);
  and_gate and_gate_h_u_cla24_and1778_y0(h_u_cla24_and1777_y0, h_u_cla24_and1776_y0, h_u_cla24_and1778_y0);
  and_gate and_gate_h_u_cla24_and1779_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and1779_y0);
  and_gate and_gate_h_u_cla24_and1780_y0(h_u_cla24_and1779_y0, h_u_cla24_and1778_y0, h_u_cla24_and1780_y0);
  and_gate and_gate_h_u_cla24_and1781_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and1781_y0);
  and_gate and_gate_h_u_cla24_and1782_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and1782_y0);
  and_gate and_gate_h_u_cla24_and1783_y0(h_u_cla24_and1782_y0, h_u_cla24_and1781_y0, h_u_cla24_and1783_y0);
  and_gate and_gate_h_u_cla24_and1784_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and1784_y0);
  or_gate or_gate_h_u_cla24_or136_y0(h_u_cla24_and1784_y0, h_u_cla24_and1528_y0, h_u_cla24_or136_y0);
  or_gate or_gate_h_u_cla24_or137_y0(h_u_cla24_or136_y0, h_u_cla24_and1559_y0, h_u_cla24_or137_y0);
  or_gate or_gate_h_u_cla24_or138_y0(h_u_cla24_or137_y0, h_u_cla24_and1588_y0, h_u_cla24_or138_y0);
  or_gate or_gate_h_u_cla24_or139_y0(h_u_cla24_or138_y0, h_u_cla24_and1615_y0, h_u_cla24_or139_y0);
  or_gate or_gate_h_u_cla24_or140_y0(h_u_cla24_or139_y0, h_u_cla24_and1640_y0, h_u_cla24_or140_y0);
  or_gate or_gate_h_u_cla24_or141_y0(h_u_cla24_or140_y0, h_u_cla24_and1663_y0, h_u_cla24_or141_y0);
  or_gate or_gate_h_u_cla24_or142_y0(h_u_cla24_or141_y0, h_u_cla24_and1684_y0, h_u_cla24_or142_y0);
  or_gate or_gate_h_u_cla24_or143_y0(h_u_cla24_or142_y0, h_u_cla24_and1703_y0, h_u_cla24_or143_y0);
  or_gate or_gate_h_u_cla24_or144_y0(h_u_cla24_or143_y0, h_u_cla24_and1720_y0, h_u_cla24_or144_y0);
  or_gate or_gate_h_u_cla24_or145_y0(h_u_cla24_or144_y0, h_u_cla24_and1735_y0, h_u_cla24_or145_y0);
  or_gate or_gate_h_u_cla24_or146_y0(h_u_cla24_or145_y0, h_u_cla24_and1748_y0, h_u_cla24_or146_y0);
  or_gate or_gate_h_u_cla24_or147_y0(h_u_cla24_or146_y0, h_u_cla24_and1759_y0, h_u_cla24_or147_y0);
  or_gate or_gate_h_u_cla24_or148_y0(h_u_cla24_or147_y0, h_u_cla24_and1768_y0, h_u_cla24_or148_y0);
  or_gate or_gate_h_u_cla24_or149_y0(h_u_cla24_or148_y0, h_u_cla24_and1775_y0, h_u_cla24_or149_y0);
  or_gate or_gate_h_u_cla24_or150_y0(h_u_cla24_or149_y0, h_u_cla24_and1780_y0, h_u_cla24_or150_y0);
  or_gate or_gate_h_u_cla24_or151_y0(h_u_cla24_or150_y0, h_u_cla24_and1783_y0, h_u_cla24_or151_y0);
  or_gate or_gate_h_u_cla24_or152_y0(h_u_cla24_pg_logic16_y1, h_u_cla24_or151_y0, h_u_cla24_or152_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic17_y0(a_17, b_17, h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_pg_logic17_y2);
  xor_gate xor_gate_h_u_cla24_xor17_y0(h_u_cla24_pg_logic17_y2, h_u_cla24_or152_y0, h_u_cla24_xor17_y0);
  and_gate and_gate_h_u_cla24_and1785_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and1785_y0);
  and_gate and_gate_h_u_cla24_and1786_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and1786_y0);
  and_gate and_gate_h_u_cla24_and1787_y0(h_u_cla24_and1786_y0, h_u_cla24_and1785_y0, h_u_cla24_and1787_y0);
  and_gate and_gate_h_u_cla24_and1788_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and1788_y0);
  and_gate and_gate_h_u_cla24_and1789_y0(h_u_cla24_and1788_y0, h_u_cla24_and1787_y0, h_u_cla24_and1789_y0);
  and_gate and_gate_h_u_cla24_and1790_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and1790_y0);
  and_gate and_gate_h_u_cla24_and1791_y0(h_u_cla24_and1790_y0, h_u_cla24_and1789_y0, h_u_cla24_and1791_y0);
  and_gate and_gate_h_u_cla24_and1792_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and1792_y0);
  and_gate and_gate_h_u_cla24_and1793_y0(h_u_cla24_and1792_y0, h_u_cla24_and1791_y0, h_u_cla24_and1793_y0);
  and_gate and_gate_h_u_cla24_and1794_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and1794_y0);
  and_gate and_gate_h_u_cla24_and1795_y0(h_u_cla24_and1794_y0, h_u_cla24_and1793_y0, h_u_cla24_and1795_y0);
  and_gate and_gate_h_u_cla24_and1796_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and1796_y0);
  and_gate and_gate_h_u_cla24_and1797_y0(h_u_cla24_and1796_y0, h_u_cla24_and1795_y0, h_u_cla24_and1797_y0);
  and_gate and_gate_h_u_cla24_and1798_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and1798_y0);
  and_gate and_gate_h_u_cla24_and1799_y0(h_u_cla24_and1798_y0, h_u_cla24_and1797_y0, h_u_cla24_and1799_y0);
  and_gate and_gate_h_u_cla24_and1800_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and1800_y0);
  and_gate and_gate_h_u_cla24_and1801_y0(h_u_cla24_and1800_y0, h_u_cla24_and1799_y0, h_u_cla24_and1801_y0);
  and_gate and_gate_h_u_cla24_and1802_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and1802_y0);
  and_gate and_gate_h_u_cla24_and1803_y0(h_u_cla24_and1802_y0, h_u_cla24_and1801_y0, h_u_cla24_and1803_y0);
  and_gate and_gate_h_u_cla24_and1804_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and1804_y0);
  and_gate and_gate_h_u_cla24_and1805_y0(h_u_cla24_and1804_y0, h_u_cla24_and1803_y0, h_u_cla24_and1805_y0);
  and_gate and_gate_h_u_cla24_and1806_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and1806_y0);
  and_gate and_gate_h_u_cla24_and1807_y0(h_u_cla24_and1806_y0, h_u_cla24_and1805_y0, h_u_cla24_and1807_y0);
  and_gate and_gate_h_u_cla24_and1808_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and1808_y0);
  and_gate and_gate_h_u_cla24_and1809_y0(h_u_cla24_and1808_y0, h_u_cla24_and1807_y0, h_u_cla24_and1809_y0);
  and_gate and_gate_h_u_cla24_and1810_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and1810_y0);
  and_gate and_gate_h_u_cla24_and1811_y0(h_u_cla24_and1810_y0, h_u_cla24_and1809_y0, h_u_cla24_and1811_y0);
  and_gate and_gate_h_u_cla24_and1812_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and1812_y0);
  and_gate and_gate_h_u_cla24_and1813_y0(h_u_cla24_and1812_y0, h_u_cla24_and1811_y0, h_u_cla24_and1813_y0);
  and_gate and_gate_h_u_cla24_and1814_y0(h_u_cla24_pg_logic15_y0, constant_wire_0, h_u_cla24_and1814_y0);
  and_gate and_gate_h_u_cla24_and1815_y0(h_u_cla24_and1814_y0, h_u_cla24_and1813_y0, h_u_cla24_and1815_y0);
  and_gate and_gate_h_u_cla24_and1816_y0(h_u_cla24_pg_logic16_y0, constant_wire_0, h_u_cla24_and1816_y0);
  and_gate and_gate_h_u_cla24_and1817_y0(h_u_cla24_and1816_y0, h_u_cla24_and1815_y0, h_u_cla24_and1817_y0);
  and_gate and_gate_h_u_cla24_and1818_y0(h_u_cla24_pg_logic17_y0, constant_wire_0, h_u_cla24_and1818_y0);
  and_gate and_gate_h_u_cla24_and1819_y0(h_u_cla24_and1818_y0, h_u_cla24_and1817_y0, h_u_cla24_and1819_y0);
  and_gate and_gate_h_u_cla24_and1820_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1820_y0);
  and_gate and_gate_h_u_cla24_and1821_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1821_y0);
  and_gate and_gate_h_u_cla24_and1822_y0(h_u_cla24_and1821_y0, h_u_cla24_and1820_y0, h_u_cla24_and1822_y0);
  and_gate and_gate_h_u_cla24_and1823_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1823_y0);
  and_gate and_gate_h_u_cla24_and1824_y0(h_u_cla24_and1823_y0, h_u_cla24_and1822_y0, h_u_cla24_and1824_y0);
  and_gate and_gate_h_u_cla24_and1825_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1825_y0);
  and_gate and_gate_h_u_cla24_and1826_y0(h_u_cla24_and1825_y0, h_u_cla24_and1824_y0, h_u_cla24_and1826_y0);
  and_gate and_gate_h_u_cla24_and1827_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1827_y0);
  and_gate and_gate_h_u_cla24_and1828_y0(h_u_cla24_and1827_y0, h_u_cla24_and1826_y0, h_u_cla24_and1828_y0);
  and_gate and_gate_h_u_cla24_and1829_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1829_y0);
  and_gate and_gate_h_u_cla24_and1830_y0(h_u_cla24_and1829_y0, h_u_cla24_and1828_y0, h_u_cla24_and1830_y0);
  and_gate and_gate_h_u_cla24_and1831_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1831_y0);
  and_gate and_gate_h_u_cla24_and1832_y0(h_u_cla24_and1831_y0, h_u_cla24_and1830_y0, h_u_cla24_and1832_y0);
  and_gate and_gate_h_u_cla24_and1833_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1833_y0);
  and_gate and_gate_h_u_cla24_and1834_y0(h_u_cla24_and1833_y0, h_u_cla24_and1832_y0, h_u_cla24_and1834_y0);
  and_gate and_gate_h_u_cla24_and1835_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1835_y0);
  and_gate and_gate_h_u_cla24_and1836_y0(h_u_cla24_and1835_y0, h_u_cla24_and1834_y0, h_u_cla24_and1836_y0);
  and_gate and_gate_h_u_cla24_and1837_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1837_y0);
  and_gate and_gate_h_u_cla24_and1838_y0(h_u_cla24_and1837_y0, h_u_cla24_and1836_y0, h_u_cla24_and1838_y0);
  and_gate and_gate_h_u_cla24_and1839_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1839_y0);
  and_gate and_gate_h_u_cla24_and1840_y0(h_u_cla24_and1839_y0, h_u_cla24_and1838_y0, h_u_cla24_and1840_y0);
  and_gate and_gate_h_u_cla24_and1841_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1841_y0);
  and_gate and_gate_h_u_cla24_and1842_y0(h_u_cla24_and1841_y0, h_u_cla24_and1840_y0, h_u_cla24_and1842_y0);
  and_gate and_gate_h_u_cla24_and1843_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1843_y0);
  and_gate and_gate_h_u_cla24_and1844_y0(h_u_cla24_and1843_y0, h_u_cla24_and1842_y0, h_u_cla24_and1844_y0);
  and_gate and_gate_h_u_cla24_and1845_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1845_y0);
  and_gate and_gate_h_u_cla24_and1846_y0(h_u_cla24_and1845_y0, h_u_cla24_and1844_y0, h_u_cla24_and1846_y0);
  and_gate and_gate_h_u_cla24_and1847_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1847_y0);
  and_gate and_gate_h_u_cla24_and1848_y0(h_u_cla24_and1847_y0, h_u_cla24_and1846_y0, h_u_cla24_and1848_y0);
  and_gate and_gate_h_u_cla24_and1849_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1849_y0);
  and_gate and_gate_h_u_cla24_and1850_y0(h_u_cla24_and1849_y0, h_u_cla24_and1848_y0, h_u_cla24_and1850_y0);
  and_gate and_gate_h_u_cla24_and1851_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and1851_y0);
  and_gate and_gate_h_u_cla24_and1852_y0(h_u_cla24_and1851_y0, h_u_cla24_and1850_y0, h_u_cla24_and1852_y0);
  and_gate and_gate_h_u_cla24_and1853_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1853_y0);
  and_gate and_gate_h_u_cla24_and1854_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1854_y0);
  and_gate and_gate_h_u_cla24_and1855_y0(h_u_cla24_and1854_y0, h_u_cla24_and1853_y0, h_u_cla24_and1855_y0);
  and_gate and_gate_h_u_cla24_and1856_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1856_y0);
  and_gate and_gate_h_u_cla24_and1857_y0(h_u_cla24_and1856_y0, h_u_cla24_and1855_y0, h_u_cla24_and1857_y0);
  and_gate and_gate_h_u_cla24_and1858_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1858_y0);
  and_gate and_gate_h_u_cla24_and1859_y0(h_u_cla24_and1858_y0, h_u_cla24_and1857_y0, h_u_cla24_and1859_y0);
  and_gate and_gate_h_u_cla24_and1860_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1860_y0);
  and_gate and_gate_h_u_cla24_and1861_y0(h_u_cla24_and1860_y0, h_u_cla24_and1859_y0, h_u_cla24_and1861_y0);
  and_gate and_gate_h_u_cla24_and1862_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1862_y0);
  and_gate and_gate_h_u_cla24_and1863_y0(h_u_cla24_and1862_y0, h_u_cla24_and1861_y0, h_u_cla24_and1863_y0);
  and_gate and_gate_h_u_cla24_and1864_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1864_y0);
  and_gate and_gate_h_u_cla24_and1865_y0(h_u_cla24_and1864_y0, h_u_cla24_and1863_y0, h_u_cla24_and1865_y0);
  and_gate and_gate_h_u_cla24_and1866_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1866_y0);
  and_gate and_gate_h_u_cla24_and1867_y0(h_u_cla24_and1866_y0, h_u_cla24_and1865_y0, h_u_cla24_and1867_y0);
  and_gate and_gate_h_u_cla24_and1868_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1868_y0);
  and_gate and_gate_h_u_cla24_and1869_y0(h_u_cla24_and1868_y0, h_u_cla24_and1867_y0, h_u_cla24_and1869_y0);
  and_gate and_gate_h_u_cla24_and1870_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1870_y0);
  and_gate and_gate_h_u_cla24_and1871_y0(h_u_cla24_and1870_y0, h_u_cla24_and1869_y0, h_u_cla24_and1871_y0);
  and_gate and_gate_h_u_cla24_and1872_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1872_y0);
  and_gate and_gate_h_u_cla24_and1873_y0(h_u_cla24_and1872_y0, h_u_cla24_and1871_y0, h_u_cla24_and1873_y0);
  and_gate and_gate_h_u_cla24_and1874_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1874_y0);
  and_gate and_gate_h_u_cla24_and1875_y0(h_u_cla24_and1874_y0, h_u_cla24_and1873_y0, h_u_cla24_and1875_y0);
  and_gate and_gate_h_u_cla24_and1876_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1876_y0);
  and_gate and_gate_h_u_cla24_and1877_y0(h_u_cla24_and1876_y0, h_u_cla24_and1875_y0, h_u_cla24_and1877_y0);
  and_gate and_gate_h_u_cla24_and1878_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1878_y0);
  and_gate and_gate_h_u_cla24_and1879_y0(h_u_cla24_and1878_y0, h_u_cla24_and1877_y0, h_u_cla24_and1879_y0);
  and_gate and_gate_h_u_cla24_and1880_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1880_y0);
  and_gate and_gate_h_u_cla24_and1881_y0(h_u_cla24_and1880_y0, h_u_cla24_and1879_y0, h_u_cla24_and1881_y0);
  and_gate and_gate_h_u_cla24_and1882_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and1882_y0);
  and_gate and_gate_h_u_cla24_and1883_y0(h_u_cla24_and1882_y0, h_u_cla24_and1881_y0, h_u_cla24_and1883_y0);
  and_gate and_gate_h_u_cla24_and1884_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1884_y0);
  and_gate and_gate_h_u_cla24_and1885_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1885_y0);
  and_gate and_gate_h_u_cla24_and1886_y0(h_u_cla24_and1885_y0, h_u_cla24_and1884_y0, h_u_cla24_and1886_y0);
  and_gate and_gate_h_u_cla24_and1887_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1887_y0);
  and_gate and_gate_h_u_cla24_and1888_y0(h_u_cla24_and1887_y0, h_u_cla24_and1886_y0, h_u_cla24_and1888_y0);
  and_gate and_gate_h_u_cla24_and1889_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1889_y0);
  and_gate and_gate_h_u_cla24_and1890_y0(h_u_cla24_and1889_y0, h_u_cla24_and1888_y0, h_u_cla24_and1890_y0);
  and_gate and_gate_h_u_cla24_and1891_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1891_y0);
  and_gate and_gate_h_u_cla24_and1892_y0(h_u_cla24_and1891_y0, h_u_cla24_and1890_y0, h_u_cla24_and1892_y0);
  and_gate and_gate_h_u_cla24_and1893_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1893_y0);
  and_gate and_gate_h_u_cla24_and1894_y0(h_u_cla24_and1893_y0, h_u_cla24_and1892_y0, h_u_cla24_and1894_y0);
  and_gate and_gate_h_u_cla24_and1895_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1895_y0);
  and_gate and_gate_h_u_cla24_and1896_y0(h_u_cla24_and1895_y0, h_u_cla24_and1894_y0, h_u_cla24_and1896_y0);
  and_gate and_gate_h_u_cla24_and1897_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1897_y0);
  and_gate and_gate_h_u_cla24_and1898_y0(h_u_cla24_and1897_y0, h_u_cla24_and1896_y0, h_u_cla24_and1898_y0);
  and_gate and_gate_h_u_cla24_and1899_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1899_y0);
  and_gate and_gate_h_u_cla24_and1900_y0(h_u_cla24_and1899_y0, h_u_cla24_and1898_y0, h_u_cla24_and1900_y0);
  and_gate and_gate_h_u_cla24_and1901_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1901_y0);
  and_gate and_gate_h_u_cla24_and1902_y0(h_u_cla24_and1901_y0, h_u_cla24_and1900_y0, h_u_cla24_and1902_y0);
  and_gate and_gate_h_u_cla24_and1903_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1903_y0);
  and_gate and_gate_h_u_cla24_and1904_y0(h_u_cla24_and1903_y0, h_u_cla24_and1902_y0, h_u_cla24_and1904_y0);
  and_gate and_gate_h_u_cla24_and1905_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1905_y0);
  and_gate and_gate_h_u_cla24_and1906_y0(h_u_cla24_and1905_y0, h_u_cla24_and1904_y0, h_u_cla24_and1906_y0);
  and_gate and_gate_h_u_cla24_and1907_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1907_y0);
  and_gate and_gate_h_u_cla24_and1908_y0(h_u_cla24_and1907_y0, h_u_cla24_and1906_y0, h_u_cla24_and1908_y0);
  and_gate and_gate_h_u_cla24_and1909_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1909_y0);
  and_gate and_gate_h_u_cla24_and1910_y0(h_u_cla24_and1909_y0, h_u_cla24_and1908_y0, h_u_cla24_and1910_y0);
  and_gate and_gate_h_u_cla24_and1911_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and1911_y0);
  and_gate and_gate_h_u_cla24_and1912_y0(h_u_cla24_and1911_y0, h_u_cla24_and1910_y0, h_u_cla24_and1912_y0);
  and_gate and_gate_h_u_cla24_and1913_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1913_y0);
  and_gate and_gate_h_u_cla24_and1914_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1914_y0);
  and_gate and_gate_h_u_cla24_and1915_y0(h_u_cla24_and1914_y0, h_u_cla24_and1913_y0, h_u_cla24_and1915_y0);
  and_gate and_gate_h_u_cla24_and1916_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1916_y0);
  and_gate and_gate_h_u_cla24_and1917_y0(h_u_cla24_and1916_y0, h_u_cla24_and1915_y0, h_u_cla24_and1917_y0);
  and_gate and_gate_h_u_cla24_and1918_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1918_y0);
  and_gate and_gate_h_u_cla24_and1919_y0(h_u_cla24_and1918_y0, h_u_cla24_and1917_y0, h_u_cla24_and1919_y0);
  and_gate and_gate_h_u_cla24_and1920_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1920_y0);
  and_gate and_gate_h_u_cla24_and1921_y0(h_u_cla24_and1920_y0, h_u_cla24_and1919_y0, h_u_cla24_and1921_y0);
  and_gate and_gate_h_u_cla24_and1922_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1922_y0);
  and_gate and_gate_h_u_cla24_and1923_y0(h_u_cla24_and1922_y0, h_u_cla24_and1921_y0, h_u_cla24_and1923_y0);
  and_gate and_gate_h_u_cla24_and1924_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1924_y0);
  and_gate and_gate_h_u_cla24_and1925_y0(h_u_cla24_and1924_y0, h_u_cla24_and1923_y0, h_u_cla24_and1925_y0);
  and_gate and_gate_h_u_cla24_and1926_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1926_y0);
  and_gate and_gate_h_u_cla24_and1927_y0(h_u_cla24_and1926_y0, h_u_cla24_and1925_y0, h_u_cla24_and1927_y0);
  and_gate and_gate_h_u_cla24_and1928_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1928_y0);
  and_gate and_gate_h_u_cla24_and1929_y0(h_u_cla24_and1928_y0, h_u_cla24_and1927_y0, h_u_cla24_and1929_y0);
  and_gate and_gate_h_u_cla24_and1930_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1930_y0);
  and_gate and_gate_h_u_cla24_and1931_y0(h_u_cla24_and1930_y0, h_u_cla24_and1929_y0, h_u_cla24_and1931_y0);
  and_gate and_gate_h_u_cla24_and1932_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1932_y0);
  and_gate and_gate_h_u_cla24_and1933_y0(h_u_cla24_and1932_y0, h_u_cla24_and1931_y0, h_u_cla24_and1933_y0);
  and_gate and_gate_h_u_cla24_and1934_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1934_y0);
  and_gate and_gate_h_u_cla24_and1935_y0(h_u_cla24_and1934_y0, h_u_cla24_and1933_y0, h_u_cla24_and1935_y0);
  and_gate and_gate_h_u_cla24_and1936_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1936_y0);
  and_gate and_gate_h_u_cla24_and1937_y0(h_u_cla24_and1936_y0, h_u_cla24_and1935_y0, h_u_cla24_and1937_y0);
  and_gate and_gate_h_u_cla24_and1938_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and1938_y0);
  and_gate and_gate_h_u_cla24_and1939_y0(h_u_cla24_and1938_y0, h_u_cla24_and1937_y0, h_u_cla24_and1939_y0);
  and_gate and_gate_h_u_cla24_and1940_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1940_y0);
  and_gate and_gate_h_u_cla24_and1941_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1941_y0);
  and_gate and_gate_h_u_cla24_and1942_y0(h_u_cla24_and1941_y0, h_u_cla24_and1940_y0, h_u_cla24_and1942_y0);
  and_gate and_gate_h_u_cla24_and1943_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1943_y0);
  and_gate and_gate_h_u_cla24_and1944_y0(h_u_cla24_and1943_y0, h_u_cla24_and1942_y0, h_u_cla24_and1944_y0);
  and_gate and_gate_h_u_cla24_and1945_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1945_y0);
  and_gate and_gate_h_u_cla24_and1946_y0(h_u_cla24_and1945_y0, h_u_cla24_and1944_y0, h_u_cla24_and1946_y0);
  and_gate and_gate_h_u_cla24_and1947_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1947_y0);
  and_gate and_gate_h_u_cla24_and1948_y0(h_u_cla24_and1947_y0, h_u_cla24_and1946_y0, h_u_cla24_and1948_y0);
  and_gate and_gate_h_u_cla24_and1949_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1949_y0);
  and_gate and_gate_h_u_cla24_and1950_y0(h_u_cla24_and1949_y0, h_u_cla24_and1948_y0, h_u_cla24_and1950_y0);
  and_gate and_gate_h_u_cla24_and1951_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1951_y0);
  and_gate and_gate_h_u_cla24_and1952_y0(h_u_cla24_and1951_y0, h_u_cla24_and1950_y0, h_u_cla24_and1952_y0);
  and_gate and_gate_h_u_cla24_and1953_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1953_y0);
  and_gate and_gate_h_u_cla24_and1954_y0(h_u_cla24_and1953_y0, h_u_cla24_and1952_y0, h_u_cla24_and1954_y0);
  and_gate and_gate_h_u_cla24_and1955_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1955_y0);
  and_gate and_gate_h_u_cla24_and1956_y0(h_u_cla24_and1955_y0, h_u_cla24_and1954_y0, h_u_cla24_and1956_y0);
  and_gate and_gate_h_u_cla24_and1957_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1957_y0);
  and_gate and_gate_h_u_cla24_and1958_y0(h_u_cla24_and1957_y0, h_u_cla24_and1956_y0, h_u_cla24_and1958_y0);
  and_gate and_gate_h_u_cla24_and1959_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1959_y0);
  and_gate and_gate_h_u_cla24_and1960_y0(h_u_cla24_and1959_y0, h_u_cla24_and1958_y0, h_u_cla24_and1960_y0);
  and_gate and_gate_h_u_cla24_and1961_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1961_y0);
  and_gate and_gate_h_u_cla24_and1962_y0(h_u_cla24_and1961_y0, h_u_cla24_and1960_y0, h_u_cla24_and1962_y0);
  and_gate and_gate_h_u_cla24_and1963_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and1963_y0);
  and_gate and_gate_h_u_cla24_and1964_y0(h_u_cla24_and1963_y0, h_u_cla24_and1962_y0, h_u_cla24_and1964_y0);
  and_gate and_gate_h_u_cla24_and1965_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1965_y0);
  and_gate and_gate_h_u_cla24_and1966_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1966_y0);
  and_gate and_gate_h_u_cla24_and1967_y0(h_u_cla24_and1966_y0, h_u_cla24_and1965_y0, h_u_cla24_and1967_y0);
  and_gate and_gate_h_u_cla24_and1968_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1968_y0);
  and_gate and_gate_h_u_cla24_and1969_y0(h_u_cla24_and1968_y0, h_u_cla24_and1967_y0, h_u_cla24_and1969_y0);
  and_gate and_gate_h_u_cla24_and1970_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1970_y0);
  and_gate and_gate_h_u_cla24_and1971_y0(h_u_cla24_and1970_y0, h_u_cla24_and1969_y0, h_u_cla24_and1971_y0);
  and_gate and_gate_h_u_cla24_and1972_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1972_y0);
  and_gate and_gate_h_u_cla24_and1973_y0(h_u_cla24_and1972_y0, h_u_cla24_and1971_y0, h_u_cla24_and1973_y0);
  and_gate and_gate_h_u_cla24_and1974_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1974_y0);
  and_gate and_gate_h_u_cla24_and1975_y0(h_u_cla24_and1974_y0, h_u_cla24_and1973_y0, h_u_cla24_and1975_y0);
  and_gate and_gate_h_u_cla24_and1976_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1976_y0);
  and_gate and_gate_h_u_cla24_and1977_y0(h_u_cla24_and1976_y0, h_u_cla24_and1975_y0, h_u_cla24_and1977_y0);
  and_gate and_gate_h_u_cla24_and1978_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1978_y0);
  and_gate and_gate_h_u_cla24_and1979_y0(h_u_cla24_and1978_y0, h_u_cla24_and1977_y0, h_u_cla24_and1979_y0);
  and_gate and_gate_h_u_cla24_and1980_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1980_y0);
  and_gate and_gate_h_u_cla24_and1981_y0(h_u_cla24_and1980_y0, h_u_cla24_and1979_y0, h_u_cla24_and1981_y0);
  and_gate and_gate_h_u_cla24_and1982_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1982_y0);
  and_gate and_gate_h_u_cla24_and1983_y0(h_u_cla24_and1982_y0, h_u_cla24_and1981_y0, h_u_cla24_and1983_y0);
  and_gate and_gate_h_u_cla24_and1984_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1984_y0);
  and_gate and_gate_h_u_cla24_and1985_y0(h_u_cla24_and1984_y0, h_u_cla24_and1983_y0, h_u_cla24_and1985_y0);
  and_gate and_gate_h_u_cla24_and1986_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and1986_y0);
  and_gate and_gate_h_u_cla24_and1987_y0(h_u_cla24_and1986_y0, h_u_cla24_and1985_y0, h_u_cla24_and1987_y0);
  and_gate and_gate_h_u_cla24_and1988_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1988_y0);
  and_gate and_gate_h_u_cla24_and1989_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1989_y0);
  and_gate and_gate_h_u_cla24_and1990_y0(h_u_cla24_and1989_y0, h_u_cla24_and1988_y0, h_u_cla24_and1990_y0);
  and_gate and_gate_h_u_cla24_and1991_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1991_y0);
  and_gate and_gate_h_u_cla24_and1992_y0(h_u_cla24_and1991_y0, h_u_cla24_and1990_y0, h_u_cla24_and1992_y0);
  and_gate and_gate_h_u_cla24_and1993_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1993_y0);
  and_gate and_gate_h_u_cla24_and1994_y0(h_u_cla24_and1993_y0, h_u_cla24_and1992_y0, h_u_cla24_and1994_y0);
  and_gate and_gate_h_u_cla24_and1995_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1995_y0);
  and_gate and_gate_h_u_cla24_and1996_y0(h_u_cla24_and1995_y0, h_u_cla24_and1994_y0, h_u_cla24_and1996_y0);
  and_gate and_gate_h_u_cla24_and1997_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1997_y0);
  and_gate and_gate_h_u_cla24_and1998_y0(h_u_cla24_and1997_y0, h_u_cla24_and1996_y0, h_u_cla24_and1998_y0);
  and_gate and_gate_h_u_cla24_and1999_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and1999_y0);
  and_gate and_gate_h_u_cla24_and2000_y0(h_u_cla24_and1999_y0, h_u_cla24_and1998_y0, h_u_cla24_and2000_y0);
  and_gate and_gate_h_u_cla24_and2001_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2001_y0);
  and_gate and_gate_h_u_cla24_and2002_y0(h_u_cla24_and2001_y0, h_u_cla24_and2000_y0, h_u_cla24_and2002_y0);
  and_gate and_gate_h_u_cla24_and2003_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2003_y0);
  and_gate and_gate_h_u_cla24_and2004_y0(h_u_cla24_and2003_y0, h_u_cla24_and2002_y0, h_u_cla24_and2004_y0);
  and_gate and_gate_h_u_cla24_and2005_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2005_y0);
  and_gate and_gate_h_u_cla24_and2006_y0(h_u_cla24_and2005_y0, h_u_cla24_and2004_y0, h_u_cla24_and2006_y0);
  and_gate and_gate_h_u_cla24_and2007_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2007_y0);
  and_gate and_gate_h_u_cla24_and2008_y0(h_u_cla24_and2007_y0, h_u_cla24_and2006_y0, h_u_cla24_and2008_y0);
  and_gate and_gate_h_u_cla24_and2009_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2009_y0);
  and_gate and_gate_h_u_cla24_and2010_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2010_y0);
  and_gate and_gate_h_u_cla24_and2011_y0(h_u_cla24_and2010_y0, h_u_cla24_and2009_y0, h_u_cla24_and2011_y0);
  and_gate and_gate_h_u_cla24_and2012_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2012_y0);
  and_gate and_gate_h_u_cla24_and2013_y0(h_u_cla24_and2012_y0, h_u_cla24_and2011_y0, h_u_cla24_and2013_y0);
  and_gate and_gate_h_u_cla24_and2014_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2014_y0);
  and_gate and_gate_h_u_cla24_and2015_y0(h_u_cla24_and2014_y0, h_u_cla24_and2013_y0, h_u_cla24_and2015_y0);
  and_gate and_gate_h_u_cla24_and2016_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2016_y0);
  and_gate and_gate_h_u_cla24_and2017_y0(h_u_cla24_and2016_y0, h_u_cla24_and2015_y0, h_u_cla24_and2017_y0);
  and_gate and_gate_h_u_cla24_and2018_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2018_y0);
  and_gate and_gate_h_u_cla24_and2019_y0(h_u_cla24_and2018_y0, h_u_cla24_and2017_y0, h_u_cla24_and2019_y0);
  and_gate and_gate_h_u_cla24_and2020_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2020_y0);
  and_gate and_gate_h_u_cla24_and2021_y0(h_u_cla24_and2020_y0, h_u_cla24_and2019_y0, h_u_cla24_and2021_y0);
  and_gate and_gate_h_u_cla24_and2022_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2022_y0);
  and_gate and_gate_h_u_cla24_and2023_y0(h_u_cla24_and2022_y0, h_u_cla24_and2021_y0, h_u_cla24_and2023_y0);
  and_gate and_gate_h_u_cla24_and2024_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2024_y0);
  and_gate and_gate_h_u_cla24_and2025_y0(h_u_cla24_and2024_y0, h_u_cla24_and2023_y0, h_u_cla24_and2025_y0);
  and_gate and_gate_h_u_cla24_and2026_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2026_y0);
  and_gate and_gate_h_u_cla24_and2027_y0(h_u_cla24_and2026_y0, h_u_cla24_and2025_y0, h_u_cla24_and2027_y0);
  and_gate and_gate_h_u_cla24_and2028_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2028_y0);
  and_gate and_gate_h_u_cla24_and2029_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2029_y0);
  and_gate and_gate_h_u_cla24_and2030_y0(h_u_cla24_and2029_y0, h_u_cla24_and2028_y0, h_u_cla24_and2030_y0);
  and_gate and_gate_h_u_cla24_and2031_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2031_y0);
  and_gate and_gate_h_u_cla24_and2032_y0(h_u_cla24_and2031_y0, h_u_cla24_and2030_y0, h_u_cla24_and2032_y0);
  and_gate and_gate_h_u_cla24_and2033_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2033_y0);
  and_gate and_gate_h_u_cla24_and2034_y0(h_u_cla24_and2033_y0, h_u_cla24_and2032_y0, h_u_cla24_and2034_y0);
  and_gate and_gate_h_u_cla24_and2035_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2035_y0);
  and_gate and_gate_h_u_cla24_and2036_y0(h_u_cla24_and2035_y0, h_u_cla24_and2034_y0, h_u_cla24_and2036_y0);
  and_gate and_gate_h_u_cla24_and2037_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2037_y0);
  and_gate and_gate_h_u_cla24_and2038_y0(h_u_cla24_and2037_y0, h_u_cla24_and2036_y0, h_u_cla24_and2038_y0);
  and_gate and_gate_h_u_cla24_and2039_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2039_y0);
  and_gate and_gate_h_u_cla24_and2040_y0(h_u_cla24_and2039_y0, h_u_cla24_and2038_y0, h_u_cla24_and2040_y0);
  and_gate and_gate_h_u_cla24_and2041_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2041_y0);
  and_gate and_gate_h_u_cla24_and2042_y0(h_u_cla24_and2041_y0, h_u_cla24_and2040_y0, h_u_cla24_and2042_y0);
  and_gate and_gate_h_u_cla24_and2043_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2043_y0);
  and_gate and_gate_h_u_cla24_and2044_y0(h_u_cla24_and2043_y0, h_u_cla24_and2042_y0, h_u_cla24_and2044_y0);
  and_gate and_gate_h_u_cla24_and2045_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2045_y0);
  and_gate and_gate_h_u_cla24_and2046_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2046_y0);
  and_gate and_gate_h_u_cla24_and2047_y0(h_u_cla24_and2046_y0, h_u_cla24_and2045_y0, h_u_cla24_and2047_y0);
  and_gate and_gate_h_u_cla24_and2048_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2048_y0);
  and_gate and_gate_h_u_cla24_and2049_y0(h_u_cla24_and2048_y0, h_u_cla24_and2047_y0, h_u_cla24_and2049_y0);
  and_gate and_gate_h_u_cla24_and2050_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2050_y0);
  and_gate and_gate_h_u_cla24_and2051_y0(h_u_cla24_and2050_y0, h_u_cla24_and2049_y0, h_u_cla24_and2051_y0);
  and_gate and_gate_h_u_cla24_and2052_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2052_y0);
  and_gate and_gate_h_u_cla24_and2053_y0(h_u_cla24_and2052_y0, h_u_cla24_and2051_y0, h_u_cla24_and2053_y0);
  and_gate and_gate_h_u_cla24_and2054_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2054_y0);
  and_gate and_gate_h_u_cla24_and2055_y0(h_u_cla24_and2054_y0, h_u_cla24_and2053_y0, h_u_cla24_and2055_y0);
  and_gate and_gate_h_u_cla24_and2056_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2056_y0);
  and_gate and_gate_h_u_cla24_and2057_y0(h_u_cla24_and2056_y0, h_u_cla24_and2055_y0, h_u_cla24_and2057_y0);
  and_gate and_gate_h_u_cla24_and2058_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2058_y0);
  and_gate and_gate_h_u_cla24_and2059_y0(h_u_cla24_and2058_y0, h_u_cla24_and2057_y0, h_u_cla24_and2059_y0);
  and_gate and_gate_h_u_cla24_and2060_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2060_y0);
  and_gate and_gate_h_u_cla24_and2061_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2061_y0);
  and_gate and_gate_h_u_cla24_and2062_y0(h_u_cla24_and2061_y0, h_u_cla24_and2060_y0, h_u_cla24_and2062_y0);
  and_gate and_gate_h_u_cla24_and2063_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2063_y0);
  and_gate and_gate_h_u_cla24_and2064_y0(h_u_cla24_and2063_y0, h_u_cla24_and2062_y0, h_u_cla24_and2064_y0);
  and_gate and_gate_h_u_cla24_and2065_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2065_y0);
  and_gate and_gate_h_u_cla24_and2066_y0(h_u_cla24_and2065_y0, h_u_cla24_and2064_y0, h_u_cla24_and2066_y0);
  and_gate and_gate_h_u_cla24_and2067_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2067_y0);
  and_gate and_gate_h_u_cla24_and2068_y0(h_u_cla24_and2067_y0, h_u_cla24_and2066_y0, h_u_cla24_and2068_y0);
  and_gate and_gate_h_u_cla24_and2069_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2069_y0);
  and_gate and_gate_h_u_cla24_and2070_y0(h_u_cla24_and2069_y0, h_u_cla24_and2068_y0, h_u_cla24_and2070_y0);
  and_gate and_gate_h_u_cla24_and2071_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2071_y0);
  and_gate and_gate_h_u_cla24_and2072_y0(h_u_cla24_and2071_y0, h_u_cla24_and2070_y0, h_u_cla24_and2072_y0);
  and_gate and_gate_h_u_cla24_and2073_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2073_y0);
  and_gate and_gate_h_u_cla24_and2074_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2074_y0);
  and_gate and_gate_h_u_cla24_and2075_y0(h_u_cla24_and2074_y0, h_u_cla24_and2073_y0, h_u_cla24_and2075_y0);
  and_gate and_gate_h_u_cla24_and2076_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2076_y0);
  and_gate and_gate_h_u_cla24_and2077_y0(h_u_cla24_and2076_y0, h_u_cla24_and2075_y0, h_u_cla24_and2077_y0);
  and_gate and_gate_h_u_cla24_and2078_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2078_y0);
  and_gate and_gate_h_u_cla24_and2079_y0(h_u_cla24_and2078_y0, h_u_cla24_and2077_y0, h_u_cla24_and2079_y0);
  and_gate and_gate_h_u_cla24_and2080_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2080_y0);
  and_gate and_gate_h_u_cla24_and2081_y0(h_u_cla24_and2080_y0, h_u_cla24_and2079_y0, h_u_cla24_and2081_y0);
  and_gate and_gate_h_u_cla24_and2082_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2082_y0);
  and_gate and_gate_h_u_cla24_and2083_y0(h_u_cla24_and2082_y0, h_u_cla24_and2081_y0, h_u_cla24_and2083_y0);
  and_gate and_gate_h_u_cla24_and2084_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2084_y0);
  and_gate and_gate_h_u_cla24_and2085_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2085_y0);
  and_gate and_gate_h_u_cla24_and2086_y0(h_u_cla24_and2085_y0, h_u_cla24_and2084_y0, h_u_cla24_and2086_y0);
  and_gate and_gate_h_u_cla24_and2087_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2087_y0);
  and_gate and_gate_h_u_cla24_and2088_y0(h_u_cla24_and2087_y0, h_u_cla24_and2086_y0, h_u_cla24_and2088_y0);
  and_gate and_gate_h_u_cla24_and2089_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2089_y0);
  and_gate and_gate_h_u_cla24_and2090_y0(h_u_cla24_and2089_y0, h_u_cla24_and2088_y0, h_u_cla24_and2090_y0);
  and_gate and_gate_h_u_cla24_and2091_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2091_y0);
  and_gate and_gate_h_u_cla24_and2092_y0(h_u_cla24_and2091_y0, h_u_cla24_and2090_y0, h_u_cla24_and2092_y0);
  and_gate and_gate_h_u_cla24_and2093_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2093_y0);
  and_gate and_gate_h_u_cla24_and2094_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2094_y0);
  and_gate and_gate_h_u_cla24_and2095_y0(h_u_cla24_and2094_y0, h_u_cla24_and2093_y0, h_u_cla24_and2095_y0);
  and_gate and_gate_h_u_cla24_and2096_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2096_y0);
  and_gate and_gate_h_u_cla24_and2097_y0(h_u_cla24_and2096_y0, h_u_cla24_and2095_y0, h_u_cla24_and2097_y0);
  and_gate and_gate_h_u_cla24_and2098_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2098_y0);
  and_gate and_gate_h_u_cla24_and2099_y0(h_u_cla24_and2098_y0, h_u_cla24_and2097_y0, h_u_cla24_and2099_y0);
  and_gate and_gate_h_u_cla24_and2100_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2100_y0);
  and_gate and_gate_h_u_cla24_and2101_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2101_y0);
  and_gate and_gate_h_u_cla24_and2102_y0(h_u_cla24_and2101_y0, h_u_cla24_and2100_y0, h_u_cla24_and2102_y0);
  and_gate and_gate_h_u_cla24_and2103_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2103_y0);
  and_gate and_gate_h_u_cla24_and2104_y0(h_u_cla24_and2103_y0, h_u_cla24_and2102_y0, h_u_cla24_and2104_y0);
  and_gate and_gate_h_u_cla24_and2105_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and2105_y0);
  and_gate and_gate_h_u_cla24_and2106_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and2106_y0);
  and_gate and_gate_h_u_cla24_and2107_y0(h_u_cla24_and2106_y0, h_u_cla24_and2105_y0, h_u_cla24_and2107_y0);
  and_gate and_gate_h_u_cla24_and2108_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and2108_y0);
  or_gate or_gate_h_u_cla24_or153_y0(h_u_cla24_and2108_y0, h_u_cla24_and1819_y0, h_u_cla24_or153_y0);
  or_gate or_gate_h_u_cla24_or154_y0(h_u_cla24_or153_y0, h_u_cla24_and1852_y0, h_u_cla24_or154_y0);
  or_gate or_gate_h_u_cla24_or155_y0(h_u_cla24_or154_y0, h_u_cla24_and1883_y0, h_u_cla24_or155_y0);
  or_gate or_gate_h_u_cla24_or156_y0(h_u_cla24_or155_y0, h_u_cla24_and1912_y0, h_u_cla24_or156_y0);
  or_gate or_gate_h_u_cla24_or157_y0(h_u_cla24_or156_y0, h_u_cla24_and1939_y0, h_u_cla24_or157_y0);
  or_gate or_gate_h_u_cla24_or158_y0(h_u_cla24_or157_y0, h_u_cla24_and1964_y0, h_u_cla24_or158_y0);
  or_gate or_gate_h_u_cla24_or159_y0(h_u_cla24_or158_y0, h_u_cla24_and1987_y0, h_u_cla24_or159_y0);
  or_gate or_gate_h_u_cla24_or160_y0(h_u_cla24_or159_y0, h_u_cla24_and2008_y0, h_u_cla24_or160_y0);
  or_gate or_gate_h_u_cla24_or161_y0(h_u_cla24_or160_y0, h_u_cla24_and2027_y0, h_u_cla24_or161_y0);
  or_gate or_gate_h_u_cla24_or162_y0(h_u_cla24_or161_y0, h_u_cla24_and2044_y0, h_u_cla24_or162_y0);
  or_gate or_gate_h_u_cla24_or163_y0(h_u_cla24_or162_y0, h_u_cla24_and2059_y0, h_u_cla24_or163_y0);
  or_gate or_gate_h_u_cla24_or164_y0(h_u_cla24_or163_y0, h_u_cla24_and2072_y0, h_u_cla24_or164_y0);
  or_gate or_gate_h_u_cla24_or165_y0(h_u_cla24_or164_y0, h_u_cla24_and2083_y0, h_u_cla24_or165_y0);
  or_gate or_gate_h_u_cla24_or166_y0(h_u_cla24_or165_y0, h_u_cla24_and2092_y0, h_u_cla24_or166_y0);
  or_gate or_gate_h_u_cla24_or167_y0(h_u_cla24_or166_y0, h_u_cla24_and2099_y0, h_u_cla24_or167_y0);
  or_gate or_gate_h_u_cla24_or168_y0(h_u_cla24_or167_y0, h_u_cla24_and2104_y0, h_u_cla24_or168_y0);
  or_gate or_gate_h_u_cla24_or169_y0(h_u_cla24_or168_y0, h_u_cla24_and2107_y0, h_u_cla24_or169_y0);
  or_gate or_gate_h_u_cla24_or170_y0(h_u_cla24_pg_logic17_y1, h_u_cla24_or169_y0, h_u_cla24_or170_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic18_y0(a_18, b_18, h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_pg_logic18_y2);
  xor_gate xor_gate_h_u_cla24_xor18_y0(h_u_cla24_pg_logic18_y2, h_u_cla24_or170_y0, h_u_cla24_xor18_y0);
  and_gate and_gate_h_u_cla24_and2109_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and2109_y0);
  and_gate and_gate_h_u_cla24_and2110_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and2110_y0);
  and_gate and_gate_h_u_cla24_and2111_y0(h_u_cla24_and2110_y0, h_u_cla24_and2109_y0, h_u_cla24_and2111_y0);
  and_gate and_gate_h_u_cla24_and2112_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and2112_y0);
  and_gate and_gate_h_u_cla24_and2113_y0(h_u_cla24_and2112_y0, h_u_cla24_and2111_y0, h_u_cla24_and2113_y0);
  and_gate and_gate_h_u_cla24_and2114_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and2114_y0);
  and_gate and_gate_h_u_cla24_and2115_y0(h_u_cla24_and2114_y0, h_u_cla24_and2113_y0, h_u_cla24_and2115_y0);
  and_gate and_gate_h_u_cla24_and2116_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and2116_y0);
  and_gate and_gate_h_u_cla24_and2117_y0(h_u_cla24_and2116_y0, h_u_cla24_and2115_y0, h_u_cla24_and2117_y0);
  and_gate and_gate_h_u_cla24_and2118_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and2118_y0);
  and_gate and_gate_h_u_cla24_and2119_y0(h_u_cla24_and2118_y0, h_u_cla24_and2117_y0, h_u_cla24_and2119_y0);
  and_gate and_gate_h_u_cla24_and2120_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and2120_y0);
  and_gate and_gate_h_u_cla24_and2121_y0(h_u_cla24_and2120_y0, h_u_cla24_and2119_y0, h_u_cla24_and2121_y0);
  and_gate and_gate_h_u_cla24_and2122_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and2122_y0);
  and_gate and_gate_h_u_cla24_and2123_y0(h_u_cla24_and2122_y0, h_u_cla24_and2121_y0, h_u_cla24_and2123_y0);
  and_gate and_gate_h_u_cla24_and2124_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and2124_y0);
  and_gate and_gate_h_u_cla24_and2125_y0(h_u_cla24_and2124_y0, h_u_cla24_and2123_y0, h_u_cla24_and2125_y0);
  and_gate and_gate_h_u_cla24_and2126_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and2126_y0);
  and_gate and_gate_h_u_cla24_and2127_y0(h_u_cla24_and2126_y0, h_u_cla24_and2125_y0, h_u_cla24_and2127_y0);
  and_gate and_gate_h_u_cla24_and2128_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and2128_y0);
  and_gate and_gate_h_u_cla24_and2129_y0(h_u_cla24_and2128_y0, h_u_cla24_and2127_y0, h_u_cla24_and2129_y0);
  and_gate and_gate_h_u_cla24_and2130_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and2130_y0);
  and_gate and_gate_h_u_cla24_and2131_y0(h_u_cla24_and2130_y0, h_u_cla24_and2129_y0, h_u_cla24_and2131_y0);
  and_gate and_gate_h_u_cla24_and2132_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and2132_y0);
  and_gate and_gate_h_u_cla24_and2133_y0(h_u_cla24_and2132_y0, h_u_cla24_and2131_y0, h_u_cla24_and2133_y0);
  and_gate and_gate_h_u_cla24_and2134_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and2134_y0);
  and_gate and_gate_h_u_cla24_and2135_y0(h_u_cla24_and2134_y0, h_u_cla24_and2133_y0, h_u_cla24_and2135_y0);
  and_gate and_gate_h_u_cla24_and2136_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and2136_y0);
  and_gate and_gate_h_u_cla24_and2137_y0(h_u_cla24_and2136_y0, h_u_cla24_and2135_y0, h_u_cla24_and2137_y0);
  and_gate and_gate_h_u_cla24_and2138_y0(h_u_cla24_pg_logic15_y0, constant_wire_0, h_u_cla24_and2138_y0);
  and_gate and_gate_h_u_cla24_and2139_y0(h_u_cla24_and2138_y0, h_u_cla24_and2137_y0, h_u_cla24_and2139_y0);
  and_gate and_gate_h_u_cla24_and2140_y0(h_u_cla24_pg_logic16_y0, constant_wire_0, h_u_cla24_and2140_y0);
  and_gate and_gate_h_u_cla24_and2141_y0(h_u_cla24_and2140_y0, h_u_cla24_and2139_y0, h_u_cla24_and2141_y0);
  and_gate and_gate_h_u_cla24_and2142_y0(h_u_cla24_pg_logic17_y0, constant_wire_0, h_u_cla24_and2142_y0);
  and_gate and_gate_h_u_cla24_and2143_y0(h_u_cla24_and2142_y0, h_u_cla24_and2141_y0, h_u_cla24_and2143_y0);
  and_gate and_gate_h_u_cla24_and2144_y0(h_u_cla24_pg_logic18_y0, constant_wire_0, h_u_cla24_and2144_y0);
  and_gate and_gate_h_u_cla24_and2145_y0(h_u_cla24_and2144_y0, h_u_cla24_and2143_y0, h_u_cla24_and2145_y0);
  and_gate and_gate_h_u_cla24_and2146_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2146_y0);
  and_gate and_gate_h_u_cla24_and2147_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2147_y0);
  and_gate and_gate_h_u_cla24_and2148_y0(h_u_cla24_and2147_y0, h_u_cla24_and2146_y0, h_u_cla24_and2148_y0);
  and_gate and_gate_h_u_cla24_and2149_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2149_y0);
  and_gate and_gate_h_u_cla24_and2150_y0(h_u_cla24_and2149_y0, h_u_cla24_and2148_y0, h_u_cla24_and2150_y0);
  and_gate and_gate_h_u_cla24_and2151_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2151_y0);
  and_gate and_gate_h_u_cla24_and2152_y0(h_u_cla24_and2151_y0, h_u_cla24_and2150_y0, h_u_cla24_and2152_y0);
  and_gate and_gate_h_u_cla24_and2153_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2153_y0);
  and_gate and_gate_h_u_cla24_and2154_y0(h_u_cla24_and2153_y0, h_u_cla24_and2152_y0, h_u_cla24_and2154_y0);
  and_gate and_gate_h_u_cla24_and2155_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2155_y0);
  and_gate and_gate_h_u_cla24_and2156_y0(h_u_cla24_and2155_y0, h_u_cla24_and2154_y0, h_u_cla24_and2156_y0);
  and_gate and_gate_h_u_cla24_and2157_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2157_y0);
  and_gate and_gate_h_u_cla24_and2158_y0(h_u_cla24_and2157_y0, h_u_cla24_and2156_y0, h_u_cla24_and2158_y0);
  and_gate and_gate_h_u_cla24_and2159_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2159_y0);
  and_gate and_gate_h_u_cla24_and2160_y0(h_u_cla24_and2159_y0, h_u_cla24_and2158_y0, h_u_cla24_and2160_y0);
  and_gate and_gate_h_u_cla24_and2161_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2161_y0);
  and_gate and_gate_h_u_cla24_and2162_y0(h_u_cla24_and2161_y0, h_u_cla24_and2160_y0, h_u_cla24_and2162_y0);
  and_gate and_gate_h_u_cla24_and2163_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2163_y0);
  and_gate and_gate_h_u_cla24_and2164_y0(h_u_cla24_and2163_y0, h_u_cla24_and2162_y0, h_u_cla24_and2164_y0);
  and_gate and_gate_h_u_cla24_and2165_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2165_y0);
  and_gate and_gate_h_u_cla24_and2166_y0(h_u_cla24_and2165_y0, h_u_cla24_and2164_y0, h_u_cla24_and2166_y0);
  and_gate and_gate_h_u_cla24_and2167_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2167_y0);
  and_gate and_gate_h_u_cla24_and2168_y0(h_u_cla24_and2167_y0, h_u_cla24_and2166_y0, h_u_cla24_and2168_y0);
  and_gate and_gate_h_u_cla24_and2169_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2169_y0);
  and_gate and_gate_h_u_cla24_and2170_y0(h_u_cla24_and2169_y0, h_u_cla24_and2168_y0, h_u_cla24_and2170_y0);
  and_gate and_gate_h_u_cla24_and2171_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2171_y0);
  and_gate and_gate_h_u_cla24_and2172_y0(h_u_cla24_and2171_y0, h_u_cla24_and2170_y0, h_u_cla24_and2172_y0);
  and_gate and_gate_h_u_cla24_and2173_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2173_y0);
  and_gate and_gate_h_u_cla24_and2174_y0(h_u_cla24_and2173_y0, h_u_cla24_and2172_y0, h_u_cla24_and2174_y0);
  and_gate and_gate_h_u_cla24_and2175_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2175_y0);
  and_gate and_gate_h_u_cla24_and2176_y0(h_u_cla24_and2175_y0, h_u_cla24_and2174_y0, h_u_cla24_and2176_y0);
  and_gate and_gate_h_u_cla24_and2177_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2177_y0);
  and_gate and_gate_h_u_cla24_and2178_y0(h_u_cla24_and2177_y0, h_u_cla24_and2176_y0, h_u_cla24_and2178_y0);
  and_gate and_gate_h_u_cla24_and2179_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2179_y0);
  and_gate and_gate_h_u_cla24_and2180_y0(h_u_cla24_and2179_y0, h_u_cla24_and2178_y0, h_u_cla24_and2180_y0);
  and_gate and_gate_h_u_cla24_and2181_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2181_y0);
  and_gate and_gate_h_u_cla24_and2182_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2182_y0);
  and_gate and_gate_h_u_cla24_and2183_y0(h_u_cla24_and2182_y0, h_u_cla24_and2181_y0, h_u_cla24_and2183_y0);
  and_gate and_gate_h_u_cla24_and2184_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2184_y0);
  and_gate and_gate_h_u_cla24_and2185_y0(h_u_cla24_and2184_y0, h_u_cla24_and2183_y0, h_u_cla24_and2185_y0);
  and_gate and_gate_h_u_cla24_and2186_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2186_y0);
  and_gate and_gate_h_u_cla24_and2187_y0(h_u_cla24_and2186_y0, h_u_cla24_and2185_y0, h_u_cla24_and2187_y0);
  and_gate and_gate_h_u_cla24_and2188_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2188_y0);
  and_gate and_gate_h_u_cla24_and2189_y0(h_u_cla24_and2188_y0, h_u_cla24_and2187_y0, h_u_cla24_and2189_y0);
  and_gate and_gate_h_u_cla24_and2190_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2190_y0);
  and_gate and_gate_h_u_cla24_and2191_y0(h_u_cla24_and2190_y0, h_u_cla24_and2189_y0, h_u_cla24_and2191_y0);
  and_gate and_gate_h_u_cla24_and2192_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2192_y0);
  and_gate and_gate_h_u_cla24_and2193_y0(h_u_cla24_and2192_y0, h_u_cla24_and2191_y0, h_u_cla24_and2193_y0);
  and_gate and_gate_h_u_cla24_and2194_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2194_y0);
  and_gate and_gate_h_u_cla24_and2195_y0(h_u_cla24_and2194_y0, h_u_cla24_and2193_y0, h_u_cla24_and2195_y0);
  and_gate and_gate_h_u_cla24_and2196_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2196_y0);
  and_gate and_gate_h_u_cla24_and2197_y0(h_u_cla24_and2196_y0, h_u_cla24_and2195_y0, h_u_cla24_and2197_y0);
  and_gate and_gate_h_u_cla24_and2198_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2198_y0);
  and_gate and_gate_h_u_cla24_and2199_y0(h_u_cla24_and2198_y0, h_u_cla24_and2197_y0, h_u_cla24_and2199_y0);
  and_gate and_gate_h_u_cla24_and2200_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2200_y0);
  and_gate and_gate_h_u_cla24_and2201_y0(h_u_cla24_and2200_y0, h_u_cla24_and2199_y0, h_u_cla24_and2201_y0);
  and_gate and_gate_h_u_cla24_and2202_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2202_y0);
  and_gate and_gate_h_u_cla24_and2203_y0(h_u_cla24_and2202_y0, h_u_cla24_and2201_y0, h_u_cla24_and2203_y0);
  and_gate and_gate_h_u_cla24_and2204_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2204_y0);
  and_gate and_gate_h_u_cla24_and2205_y0(h_u_cla24_and2204_y0, h_u_cla24_and2203_y0, h_u_cla24_and2205_y0);
  and_gate and_gate_h_u_cla24_and2206_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2206_y0);
  and_gate and_gate_h_u_cla24_and2207_y0(h_u_cla24_and2206_y0, h_u_cla24_and2205_y0, h_u_cla24_and2207_y0);
  and_gate and_gate_h_u_cla24_and2208_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2208_y0);
  and_gate and_gate_h_u_cla24_and2209_y0(h_u_cla24_and2208_y0, h_u_cla24_and2207_y0, h_u_cla24_and2209_y0);
  and_gate and_gate_h_u_cla24_and2210_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2210_y0);
  and_gate and_gate_h_u_cla24_and2211_y0(h_u_cla24_and2210_y0, h_u_cla24_and2209_y0, h_u_cla24_and2211_y0);
  and_gate and_gate_h_u_cla24_and2212_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2212_y0);
  and_gate and_gate_h_u_cla24_and2213_y0(h_u_cla24_and2212_y0, h_u_cla24_and2211_y0, h_u_cla24_and2213_y0);
  and_gate and_gate_h_u_cla24_and2214_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2214_y0);
  and_gate and_gate_h_u_cla24_and2215_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2215_y0);
  and_gate and_gate_h_u_cla24_and2216_y0(h_u_cla24_and2215_y0, h_u_cla24_and2214_y0, h_u_cla24_and2216_y0);
  and_gate and_gate_h_u_cla24_and2217_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2217_y0);
  and_gate and_gate_h_u_cla24_and2218_y0(h_u_cla24_and2217_y0, h_u_cla24_and2216_y0, h_u_cla24_and2218_y0);
  and_gate and_gate_h_u_cla24_and2219_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2219_y0);
  and_gate and_gate_h_u_cla24_and2220_y0(h_u_cla24_and2219_y0, h_u_cla24_and2218_y0, h_u_cla24_and2220_y0);
  and_gate and_gate_h_u_cla24_and2221_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2221_y0);
  and_gate and_gate_h_u_cla24_and2222_y0(h_u_cla24_and2221_y0, h_u_cla24_and2220_y0, h_u_cla24_and2222_y0);
  and_gate and_gate_h_u_cla24_and2223_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2223_y0);
  and_gate and_gate_h_u_cla24_and2224_y0(h_u_cla24_and2223_y0, h_u_cla24_and2222_y0, h_u_cla24_and2224_y0);
  and_gate and_gate_h_u_cla24_and2225_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2225_y0);
  and_gate and_gate_h_u_cla24_and2226_y0(h_u_cla24_and2225_y0, h_u_cla24_and2224_y0, h_u_cla24_and2226_y0);
  and_gate and_gate_h_u_cla24_and2227_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2227_y0);
  and_gate and_gate_h_u_cla24_and2228_y0(h_u_cla24_and2227_y0, h_u_cla24_and2226_y0, h_u_cla24_and2228_y0);
  and_gate and_gate_h_u_cla24_and2229_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2229_y0);
  and_gate and_gate_h_u_cla24_and2230_y0(h_u_cla24_and2229_y0, h_u_cla24_and2228_y0, h_u_cla24_and2230_y0);
  and_gate and_gate_h_u_cla24_and2231_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2231_y0);
  and_gate and_gate_h_u_cla24_and2232_y0(h_u_cla24_and2231_y0, h_u_cla24_and2230_y0, h_u_cla24_and2232_y0);
  and_gate and_gate_h_u_cla24_and2233_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2233_y0);
  and_gate and_gate_h_u_cla24_and2234_y0(h_u_cla24_and2233_y0, h_u_cla24_and2232_y0, h_u_cla24_and2234_y0);
  and_gate and_gate_h_u_cla24_and2235_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2235_y0);
  and_gate and_gate_h_u_cla24_and2236_y0(h_u_cla24_and2235_y0, h_u_cla24_and2234_y0, h_u_cla24_and2236_y0);
  and_gate and_gate_h_u_cla24_and2237_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2237_y0);
  and_gate and_gate_h_u_cla24_and2238_y0(h_u_cla24_and2237_y0, h_u_cla24_and2236_y0, h_u_cla24_and2238_y0);
  and_gate and_gate_h_u_cla24_and2239_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2239_y0);
  and_gate and_gate_h_u_cla24_and2240_y0(h_u_cla24_and2239_y0, h_u_cla24_and2238_y0, h_u_cla24_and2240_y0);
  and_gate and_gate_h_u_cla24_and2241_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2241_y0);
  and_gate and_gate_h_u_cla24_and2242_y0(h_u_cla24_and2241_y0, h_u_cla24_and2240_y0, h_u_cla24_and2242_y0);
  and_gate and_gate_h_u_cla24_and2243_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2243_y0);
  and_gate and_gate_h_u_cla24_and2244_y0(h_u_cla24_and2243_y0, h_u_cla24_and2242_y0, h_u_cla24_and2244_y0);
  and_gate and_gate_h_u_cla24_and2245_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2245_y0);
  and_gate and_gate_h_u_cla24_and2246_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2246_y0);
  and_gate and_gate_h_u_cla24_and2247_y0(h_u_cla24_and2246_y0, h_u_cla24_and2245_y0, h_u_cla24_and2247_y0);
  and_gate and_gate_h_u_cla24_and2248_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2248_y0);
  and_gate and_gate_h_u_cla24_and2249_y0(h_u_cla24_and2248_y0, h_u_cla24_and2247_y0, h_u_cla24_and2249_y0);
  and_gate and_gate_h_u_cla24_and2250_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2250_y0);
  and_gate and_gate_h_u_cla24_and2251_y0(h_u_cla24_and2250_y0, h_u_cla24_and2249_y0, h_u_cla24_and2251_y0);
  and_gate and_gate_h_u_cla24_and2252_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2252_y0);
  and_gate and_gate_h_u_cla24_and2253_y0(h_u_cla24_and2252_y0, h_u_cla24_and2251_y0, h_u_cla24_and2253_y0);
  and_gate and_gate_h_u_cla24_and2254_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2254_y0);
  and_gate and_gate_h_u_cla24_and2255_y0(h_u_cla24_and2254_y0, h_u_cla24_and2253_y0, h_u_cla24_and2255_y0);
  and_gate and_gate_h_u_cla24_and2256_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2256_y0);
  and_gate and_gate_h_u_cla24_and2257_y0(h_u_cla24_and2256_y0, h_u_cla24_and2255_y0, h_u_cla24_and2257_y0);
  and_gate and_gate_h_u_cla24_and2258_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2258_y0);
  and_gate and_gate_h_u_cla24_and2259_y0(h_u_cla24_and2258_y0, h_u_cla24_and2257_y0, h_u_cla24_and2259_y0);
  and_gate and_gate_h_u_cla24_and2260_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2260_y0);
  and_gate and_gate_h_u_cla24_and2261_y0(h_u_cla24_and2260_y0, h_u_cla24_and2259_y0, h_u_cla24_and2261_y0);
  and_gate and_gate_h_u_cla24_and2262_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2262_y0);
  and_gate and_gate_h_u_cla24_and2263_y0(h_u_cla24_and2262_y0, h_u_cla24_and2261_y0, h_u_cla24_and2263_y0);
  and_gate and_gate_h_u_cla24_and2264_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2264_y0);
  and_gate and_gate_h_u_cla24_and2265_y0(h_u_cla24_and2264_y0, h_u_cla24_and2263_y0, h_u_cla24_and2265_y0);
  and_gate and_gate_h_u_cla24_and2266_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2266_y0);
  and_gate and_gate_h_u_cla24_and2267_y0(h_u_cla24_and2266_y0, h_u_cla24_and2265_y0, h_u_cla24_and2267_y0);
  and_gate and_gate_h_u_cla24_and2268_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2268_y0);
  and_gate and_gate_h_u_cla24_and2269_y0(h_u_cla24_and2268_y0, h_u_cla24_and2267_y0, h_u_cla24_and2269_y0);
  and_gate and_gate_h_u_cla24_and2270_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2270_y0);
  and_gate and_gate_h_u_cla24_and2271_y0(h_u_cla24_and2270_y0, h_u_cla24_and2269_y0, h_u_cla24_and2271_y0);
  and_gate and_gate_h_u_cla24_and2272_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2272_y0);
  and_gate and_gate_h_u_cla24_and2273_y0(h_u_cla24_and2272_y0, h_u_cla24_and2271_y0, h_u_cla24_and2273_y0);
  and_gate and_gate_h_u_cla24_and2274_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2274_y0);
  and_gate and_gate_h_u_cla24_and2275_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2275_y0);
  and_gate and_gate_h_u_cla24_and2276_y0(h_u_cla24_and2275_y0, h_u_cla24_and2274_y0, h_u_cla24_and2276_y0);
  and_gate and_gate_h_u_cla24_and2277_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2277_y0);
  and_gate and_gate_h_u_cla24_and2278_y0(h_u_cla24_and2277_y0, h_u_cla24_and2276_y0, h_u_cla24_and2278_y0);
  and_gate and_gate_h_u_cla24_and2279_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2279_y0);
  and_gate and_gate_h_u_cla24_and2280_y0(h_u_cla24_and2279_y0, h_u_cla24_and2278_y0, h_u_cla24_and2280_y0);
  and_gate and_gate_h_u_cla24_and2281_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2281_y0);
  and_gate and_gate_h_u_cla24_and2282_y0(h_u_cla24_and2281_y0, h_u_cla24_and2280_y0, h_u_cla24_and2282_y0);
  and_gate and_gate_h_u_cla24_and2283_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2283_y0);
  and_gate and_gate_h_u_cla24_and2284_y0(h_u_cla24_and2283_y0, h_u_cla24_and2282_y0, h_u_cla24_and2284_y0);
  and_gate and_gate_h_u_cla24_and2285_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2285_y0);
  and_gate and_gate_h_u_cla24_and2286_y0(h_u_cla24_and2285_y0, h_u_cla24_and2284_y0, h_u_cla24_and2286_y0);
  and_gate and_gate_h_u_cla24_and2287_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2287_y0);
  and_gate and_gate_h_u_cla24_and2288_y0(h_u_cla24_and2287_y0, h_u_cla24_and2286_y0, h_u_cla24_and2288_y0);
  and_gate and_gate_h_u_cla24_and2289_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2289_y0);
  and_gate and_gate_h_u_cla24_and2290_y0(h_u_cla24_and2289_y0, h_u_cla24_and2288_y0, h_u_cla24_and2290_y0);
  and_gate and_gate_h_u_cla24_and2291_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2291_y0);
  and_gate and_gate_h_u_cla24_and2292_y0(h_u_cla24_and2291_y0, h_u_cla24_and2290_y0, h_u_cla24_and2292_y0);
  and_gate and_gate_h_u_cla24_and2293_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2293_y0);
  and_gate and_gate_h_u_cla24_and2294_y0(h_u_cla24_and2293_y0, h_u_cla24_and2292_y0, h_u_cla24_and2294_y0);
  and_gate and_gate_h_u_cla24_and2295_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2295_y0);
  and_gate and_gate_h_u_cla24_and2296_y0(h_u_cla24_and2295_y0, h_u_cla24_and2294_y0, h_u_cla24_and2296_y0);
  and_gate and_gate_h_u_cla24_and2297_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2297_y0);
  and_gate and_gate_h_u_cla24_and2298_y0(h_u_cla24_and2297_y0, h_u_cla24_and2296_y0, h_u_cla24_and2298_y0);
  and_gate and_gate_h_u_cla24_and2299_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2299_y0);
  and_gate and_gate_h_u_cla24_and2300_y0(h_u_cla24_and2299_y0, h_u_cla24_and2298_y0, h_u_cla24_and2300_y0);
  and_gate and_gate_h_u_cla24_and2301_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2301_y0);
  and_gate and_gate_h_u_cla24_and2302_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2302_y0);
  and_gate and_gate_h_u_cla24_and2303_y0(h_u_cla24_and2302_y0, h_u_cla24_and2301_y0, h_u_cla24_and2303_y0);
  and_gate and_gate_h_u_cla24_and2304_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2304_y0);
  and_gate and_gate_h_u_cla24_and2305_y0(h_u_cla24_and2304_y0, h_u_cla24_and2303_y0, h_u_cla24_and2305_y0);
  and_gate and_gate_h_u_cla24_and2306_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2306_y0);
  and_gate and_gate_h_u_cla24_and2307_y0(h_u_cla24_and2306_y0, h_u_cla24_and2305_y0, h_u_cla24_and2307_y0);
  and_gate and_gate_h_u_cla24_and2308_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2308_y0);
  and_gate and_gate_h_u_cla24_and2309_y0(h_u_cla24_and2308_y0, h_u_cla24_and2307_y0, h_u_cla24_and2309_y0);
  and_gate and_gate_h_u_cla24_and2310_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2310_y0);
  and_gate and_gate_h_u_cla24_and2311_y0(h_u_cla24_and2310_y0, h_u_cla24_and2309_y0, h_u_cla24_and2311_y0);
  and_gate and_gate_h_u_cla24_and2312_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2312_y0);
  and_gate and_gate_h_u_cla24_and2313_y0(h_u_cla24_and2312_y0, h_u_cla24_and2311_y0, h_u_cla24_and2313_y0);
  and_gate and_gate_h_u_cla24_and2314_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2314_y0);
  and_gate and_gate_h_u_cla24_and2315_y0(h_u_cla24_and2314_y0, h_u_cla24_and2313_y0, h_u_cla24_and2315_y0);
  and_gate and_gate_h_u_cla24_and2316_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2316_y0);
  and_gate and_gate_h_u_cla24_and2317_y0(h_u_cla24_and2316_y0, h_u_cla24_and2315_y0, h_u_cla24_and2317_y0);
  and_gate and_gate_h_u_cla24_and2318_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2318_y0);
  and_gate and_gate_h_u_cla24_and2319_y0(h_u_cla24_and2318_y0, h_u_cla24_and2317_y0, h_u_cla24_and2319_y0);
  and_gate and_gate_h_u_cla24_and2320_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2320_y0);
  and_gate and_gate_h_u_cla24_and2321_y0(h_u_cla24_and2320_y0, h_u_cla24_and2319_y0, h_u_cla24_and2321_y0);
  and_gate and_gate_h_u_cla24_and2322_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2322_y0);
  and_gate and_gate_h_u_cla24_and2323_y0(h_u_cla24_and2322_y0, h_u_cla24_and2321_y0, h_u_cla24_and2323_y0);
  and_gate and_gate_h_u_cla24_and2324_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2324_y0);
  and_gate and_gate_h_u_cla24_and2325_y0(h_u_cla24_and2324_y0, h_u_cla24_and2323_y0, h_u_cla24_and2325_y0);
  and_gate and_gate_h_u_cla24_and2326_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2326_y0);
  and_gate and_gate_h_u_cla24_and2327_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2327_y0);
  and_gate and_gate_h_u_cla24_and2328_y0(h_u_cla24_and2327_y0, h_u_cla24_and2326_y0, h_u_cla24_and2328_y0);
  and_gate and_gate_h_u_cla24_and2329_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2329_y0);
  and_gate and_gate_h_u_cla24_and2330_y0(h_u_cla24_and2329_y0, h_u_cla24_and2328_y0, h_u_cla24_and2330_y0);
  and_gate and_gate_h_u_cla24_and2331_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2331_y0);
  and_gate and_gate_h_u_cla24_and2332_y0(h_u_cla24_and2331_y0, h_u_cla24_and2330_y0, h_u_cla24_and2332_y0);
  and_gate and_gate_h_u_cla24_and2333_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2333_y0);
  and_gate and_gate_h_u_cla24_and2334_y0(h_u_cla24_and2333_y0, h_u_cla24_and2332_y0, h_u_cla24_and2334_y0);
  and_gate and_gate_h_u_cla24_and2335_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2335_y0);
  and_gate and_gate_h_u_cla24_and2336_y0(h_u_cla24_and2335_y0, h_u_cla24_and2334_y0, h_u_cla24_and2336_y0);
  and_gate and_gate_h_u_cla24_and2337_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2337_y0);
  and_gate and_gate_h_u_cla24_and2338_y0(h_u_cla24_and2337_y0, h_u_cla24_and2336_y0, h_u_cla24_and2338_y0);
  and_gate and_gate_h_u_cla24_and2339_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2339_y0);
  and_gate and_gate_h_u_cla24_and2340_y0(h_u_cla24_and2339_y0, h_u_cla24_and2338_y0, h_u_cla24_and2340_y0);
  and_gate and_gate_h_u_cla24_and2341_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2341_y0);
  and_gate and_gate_h_u_cla24_and2342_y0(h_u_cla24_and2341_y0, h_u_cla24_and2340_y0, h_u_cla24_and2342_y0);
  and_gate and_gate_h_u_cla24_and2343_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2343_y0);
  and_gate and_gate_h_u_cla24_and2344_y0(h_u_cla24_and2343_y0, h_u_cla24_and2342_y0, h_u_cla24_and2344_y0);
  and_gate and_gate_h_u_cla24_and2345_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2345_y0);
  and_gate and_gate_h_u_cla24_and2346_y0(h_u_cla24_and2345_y0, h_u_cla24_and2344_y0, h_u_cla24_and2346_y0);
  and_gate and_gate_h_u_cla24_and2347_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2347_y0);
  and_gate and_gate_h_u_cla24_and2348_y0(h_u_cla24_and2347_y0, h_u_cla24_and2346_y0, h_u_cla24_and2348_y0);
  and_gate and_gate_h_u_cla24_and2349_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2349_y0);
  and_gate and_gate_h_u_cla24_and2350_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2350_y0);
  and_gate and_gate_h_u_cla24_and2351_y0(h_u_cla24_and2350_y0, h_u_cla24_and2349_y0, h_u_cla24_and2351_y0);
  and_gate and_gate_h_u_cla24_and2352_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2352_y0);
  and_gate and_gate_h_u_cla24_and2353_y0(h_u_cla24_and2352_y0, h_u_cla24_and2351_y0, h_u_cla24_and2353_y0);
  and_gate and_gate_h_u_cla24_and2354_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2354_y0);
  and_gate and_gate_h_u_cla24_and2355_y0(h_u_cla24_and2354_y0, h_u_cla24_and2353_y0, h_u_cla24_and2355_y0);
  and_gate and_gate_h_u_cla24_and2356_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2356_y0);
  and_gate and_gate_h_u_cla24_and2357_y0(h_u_cla24_and2356_y0, h_u_cla24_and2355_y0, h_u_cla24_and2357_y0);
  and_gate and_gate_h_u_cla24_and2358_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2358_y0);
  and_gate and_gate_h_u_cla24_and2359_y0(h_u_cla24_and2358_y0, h_u_cla24_and2357_y0, h_u_cla24_and2359_y0);
  and_gate and_gate_h_u_cla24_and2360_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2360_y0);
  and_gate and_gate_h_u_cla24_and2361_y0(h_u_cla24_and2360_y0, h_u_cla24_and2359_y0, h_u_cla24_and2361_y0);
  and_gate and_gate_h_u_cla24_and2362_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2362_y0);
  and_gate and_gate_h_u_cla24_and2363_y0(h_u_cla24_and2362_y0, h_u_cla24_and2361_y0, h_u_cla24_and2363_y0);
  and_gate and_gate_h_u_cla24_and2364_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2364_y0);
  and_gate and_gate_h_u_cla24_and2365_y0(h_u_cla24_and2364_y0, h_u_cla24_and2363_y0, h_u_cla24_and2365_y0);
  and_gate and_gate_h_u_cla24_and2366_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2366_y0);
  and_gate and_gate_h_u_cla24_and2367_y0(h_u_cla24_and2366_y0, h_u_cla24_and2365_y0, h_u_cla24_and2367_y0);
  and_gate and_gate_h_u_cla24_and2368_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2368_y0);
  and_gate and_gate_h_u_cla24_and2369_y0(h_u_cla24_and2368_y0, h_u_cla24_and2367_y0, h_u_cla24_and2369_y0);
  and_gate and_gate_h_u_cla24_and2370_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2370_y0);
  and_gate and_gate_h_u_cla24_and2371_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2371_y0);
  and_gate and_gate_h_u_cla24_and2372_y0(h_u_cla24_and2371_y0, h_u_cla24_and2370_y0, h_u_cla24_and2372_y0);
  and_gate and_gate_h_u_cla24_and2373_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2373_y0);
  and_gate and_gate_h_u_cla24_and2374_y0(h_u_cla24_and2373_y0, h_u_cla24_and2372_y0, h_u_cla24_and2374_y0);
  and_gate and_gate_h_u_cla24_and2375_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2375_y0);
  and_gate and_gate_h_u_cla24_and2376_y0(h_u_cla24_and2375_y0, h_u_cla24_and2374_y0, h_u_cla24_and2376_y0);
  and_gate and_gate_h_u_cla24_and2377_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2377_y0);
  and_gate and_gate_h_u_cla24_and2378_y0(h_u_cla24_and2377_y0, h_u_cla24_and2376_y0, h_u_cla24_and2378_y0);
  and_gate and_gate_h_u_cla24_and2379_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2379_y0);
  and_gate and_gate_h_u_cla24_and2380_y0(h_u_cla24_and2379_y0, h_u_cla24_and2378_y0, h_u_cla24_and2380_y0);
  and_gate and_gate_h_u_cla24_and2381_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2381_y0);
  and_gate and_gate_h_u_cla24_and2382_y0(h_u_cla24_and2381_y0, h_u_cla24_and2380_y0, h_u_cla24_and2382_y0);
  and_gate and_gate_h_u_cla24_and2383_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2383_y0);
  and_gate and_gate_h_u_cla24_and2384_y0(h_u_cla24_and2383_y0, h_u_cla24_and2382_y0, h_u_cla24_and2384_y0);
  and_gate and_gate_h_u_cla24_and2385_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2385_y0);
  and_gate and_gate_h_u_cla24_and2386_y0(h_u_cla24_and2385_y0, h_u_cla24_and2384_y0, h_u_cla24_and2386_y0);
  and_gate and_gate_h_u_cla24_and2387_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2387_y0);
  and_gate and_gate_h_u_cla24_and2388_y0(h_u_cla24_and2387_y0, h_u_cla24_and2386_y0, h_u_cla24_and2388_y0);
  and_gate and_gate_h_u_cla24_and2389_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2389_y0);
  and_gate and_gate_h_u_cla24_and2390_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2390_y0);
  and_gate and_gate_h_u_cla24_and2391_y0(h_u_cla24_and2390_y0, h_u_cla24_and2389_y0, h_u_cla24_and2391_y0);
  and_gate and_gate_h_u_cla24_and2392_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2392_y0);
  and_gate and_gate_h_u_cla24_and2393_y0(h_u_cla24_and2392_y0, h_u_cla24_and2391_y0, h_u_cla24_and2393_y0);
  and_gate and_gate_h_u_cla24_and2394_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2394_y0);
  and_gate and_gate_h_u_cla24_and2395_y0(h_u_cla24_and2394_y0, h_u_cla24_and2393_y0, h_u_cla24_and2395_y0);
  and_gate and_gate_h_u_cla24_and2396_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2396_y0);
  and_gate and_gate_h_u_cla24_and2397_y0(h_u_cla24_and2396_y0, h_u_cla24_and2395_y0, h_u_cla24_and2397_y0);
  and_gate and_gate_h_u_cla24_and2398_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2398_y0);
  and_gate and_gate_h_u_cla24_and2399_y0(h_u_cla24_and2398_y0, h_u_cla24_and2397_y0, h_u_cla24_and2399_y0);
  and_gate and_gate_h_u_cla24_and2400_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2400_y0);
  and_gate and_gate_h_u_cla24_and2401_y0(h_u_cla24_and2400_y0, h_u_cla24_and2399_y0, h_u_cla24_and2401_y0);
  and_gate and_gate_h_u_cla24_and2402_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2402_y0);
  and_gate and_gate_h_u_cla24_and2403_y0(h_u_cla24_and2402_y0, h_u_cla24_and2401_y0, h_u_cla24_and2403_y0);
  and_gate and_gate_h_u_cla24_and2404_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2404_y0);
  and_gate and_gate_h_u_cla24_and2405_y0(h_u_cla24_and2404_y0, h_u_cla24_and2403_y0, h_u_cla24_and2405_y0);
  and_gate and_gate_h_u_cla24_and2406_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2406_y0);
  and_gate and_gate_h_u_cla24_and2407_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2407_y0);
  and_gate and_gate_h_u_cla24_and2408_y0(h_u_cla24_and2407_y0, h_u_cla24_and2406_y0, h_u_cla24_and2408_y0);
  and_gate and_gate_h_u_cla24_and2409_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2409_y0);
  and_gate and_gate_h_u_cla24_and2410_y0(h_u_cla24_and2409_y0, h_u_cla24_and2408_y0, h_u_cla24_and2410_y0);
  and_gate and_gate_h_u_cla24_and2411_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2411_y0);
  and_gate and_gate_h_u_cla24_and2412_y0(h_u_cla24_and2411_y0, h_u_cla24_and2410_y0, h_u_cla24_and2412_y0);
  and_gate and_gate_h_u_cla24_and2413_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2413_y0);
  and_gate and_gate_h_u_cla24_and2414_y0(h_u_cla24_and2413_y0, h_u_cla24_and2412_y0, h_u_cla24_and2414_y0);
  and_gate and_gate_h_u_cla24_and2415_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2415_y0);
  and_gate and_gate_h_u_cla24_and2416_y0(h_u_cla24_and2415_y0, h_u_cla24_and2414_y0, h_u_cla24_and2416_y0);
  and_gate and_gate_h_u_cla24_and2417_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2417_y0);
  and_gate and_gate_h_u_cla24_and2418_y0(h_u_cla24_and2417_y0, h_u_cla24_and2416_y0, h_u_cla24_and2418_y0);
  and_gate and_gate_h_u_cla24_and2419_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2419_y0);
  and_gate and_gate_h_u_cla24_and2420_y0(h_u_cla24_and2419_y0, h_u_cla24_and2418_y0, h_u_cla24_and2420_y0);
  and_gate and_gate_h_u_cla24_and2421_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2421_y0);
  and_gate and_gate_h_u_cla24_and2422_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2422_y0);
  and_gate and_gate_h_u_cla24_and2423_y0(h_u_cla24_and2422_y0, h_u_cla24_and2421_y0, h_u_cla24_and2423_y0);
  and_gate and_gate_h_u_cla24_and2424_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2424_y0);
  and_gate and_gate_h_u_cla24_and2425_y0(h_u_cla24_and2424_y0, h_u_cla24_and2423_y0, h_u_cla24_and2425_y0);
  and_gate and_gate_h_u_cla24_and2426_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2426_y0);
  and_gate and_gate_h_u_cla24_and2427_y0(h_u_cla24_and2426_y0, h_u_cla24_and2425_y0, h_u_cla24_and2427_y0);
  and_gate and_gate_h_u_cla24_and2428_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2428_y0);
  and_gate and_gate_h_u_cla24_and2429_y0(h_u_cla24_and2428_y0, h_u_cla24_and2427_y0, h_u_cla24_and2429_y0);
  and_gate and_gate_h_u_cla24_and2430_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2430_y0);
  and_gate and_gate_h_u_cla24_and2431_y0(h_u_cla24_and2430_y0, h_u_cla24_and2429_y0, h_u_cla24_and2431_y0);
  and_gate and_gate_h_u_cla24_and2432_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2432_y0);
  and_gate and_gate_h_u_cla24_and2433_y0(h_u_cla24_and2432_y0, h_u_cla24_and2431_y0, h_u_cla24_and2433_y0);
  and_gate and_gate_h_u_cla24_and2434_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2434_y0);
  and_gate and_gate_h_u_cla24_and2435_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2435_y0);
  and_gate and_gate_h_u_cla24_and2436_y0(h_u_cla24_and2435_y0, h_u_cla24_and2434_y0, h_u_cla24_and2436_y0);
  and_gate and_gate_h_u_cla24_and2437_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2437_y0);
  and_gate and_gate_h_u_cla24_and2438_y0(h_u_cla24_and2437_y0, h_u_cla24_and2436_y0, h_u_cla24_and2438_y0);
  and_gate and_gate_h_u_cla24_and2439_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2439_y0);
  and_gate and_gate_h_u_cla24_and2440_y0(h_u_cla24_and2439_y0, h_u_cla24_and2438_y0, h_u_cla24_and2440_y0);
  and_gate and_gate_h_u_cla24_and2441_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2441_y0);
  and_gate and_gate_h_u_cla24_and2442_y0(h_u_cla24_and2441_y0, h_u_cla24_and2440_y0, h_u_cla24_and2442_y0);
  and_gate and_gate_h_u_cla24_and2443_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2443_y0);
  and_gate and_gate_h_u_cla24_and2444_y0(h_u_cla24_and2443_y0, h_u_cla24_and2442_y0, h_u_cla24_and2444_y0);
  and_gate and_gate_h_u_cla24_and2445_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2445_y0);
  and_gate and_gate_h_u_cla24_and2446_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2446_y0);
  and_gate and_gate_h_u_cla24_and2447_y0(h_u_cla24_and2446_y0, h_u_cla24_and2445_y0, h_u_cla24_and2447_y0);
  and_gate and_gate_h_u_cla24_and2448_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2448_y0);
  and_gate and_gate_h_u_cla24_and2449_y0(h_u_cla24_and2448_y0, h_u_cla24_and2447_y0, h_u_cla24_and2449_y0);
  and_gate and_gate_h_u_cla24_and2450_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2450_y0);
  and_gate and_gate_h_u_cla24_and2451_y0(h_u_cla24_and2450_y0, h_u_cla24_and2449_y0, h_u_cla24_and2451_y0);
  and_gate and_gate_h_u_cla24_and2452_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2452_y0);
  and_gate and_gate_h_u_cla24_and2453_y0(h_u_cla24_and2452_y0, h_u_cla24_and2451_y0, h_u_cla24_and2453_y0);
  and_gate and_gate_h_u_cla24_and2454_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2454_y0);
  and_gate and_gate_h_u_cla24_and2455_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2455_y0);
  and_gate and_gate_h_u_cla24_and2456_y0(h_u_cla24_and2455_y0, h_u_cla24_and2454_y0, h_u_cla24_and2456_y0);
  and_gate and_gate_h_u_cla24_and2457_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2457_y0);
  and_gate and_gate_h_u_cla24_and2458_y0(h_u_cla24_and2457_y0, h_u_cla24_and2456_y0, h_u_cla24_and2458_y0);
  and_gate and_gate_h_u_cla24_and2459_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2459_y0);
  and_gate and_gate_h_u_cla24_and2460_y0(h_u_cla24_and2459_y0, h_u_cla24_and2458_y0, h_u_cla24_and2460_y0);
  and_gate and_gate_h_u_cla24_and2461_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and2461_y0);
  and_gate and_gate_h_u_cla24_and2462_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and2462_y0);
  and_gate and_gate_h_u_cla24_and2463_y0(h_u_cla24_and2462_y0, h_u_cla24_and2461_y0, h_u_cla24_and2463_y0);
  and_gate and_gate_h_u_cla24_and2464_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and2464_y0);
  and_gate and_gate_h_u_cla24_and2465_y0(h_u_cla24_and2464_y0, h_u_cla24_and2463_y0, h_u_cla24_and2465_y0);
  and_gate and_gate_h_u_cla24_and2466_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and2466_y0);
  and_gate and_gate_h_u_cla24_and2467_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and2467_y0);
  and_gate and_gate_h_u_cla24_and2468_y0(h_u_cla24_and2467_y0, h_u_cla24_and2466_y0, h_u_cla24_and2468_y0);
  and_gate and_gate_h_u_cla24_and2469_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and2469_y0);
  or_gate or_gate_h_u_cla24_or171_y0(h_u_cla24_and2469_y0, h_u_cla24_and2145_y0, h_u_cla24_or171_y0);
  or_gate or_gate_h_u_cla24_or172_y0(h_u_cla24_or171_y0, h_u_cla24_and2180_y0, h_u_cla24_or172_y0);
  or_gate or_gate_h_u_cla24_or173_y0(h_u_cla24_or172_y0, h_u_cla24_and2213_y0, h_u_cla24_or173_y0);
  or_gate or_gate_h_u_cla24_or174_y0(h_u_cla24_or173_y0, h_u_cla24_and2244_y0, h_u_cla24_or174_y0);
  or_gate or_gate_h_u_cla24_or175_y0(h_u_cla24_or174_y0, h_u_cla24_and2273_y0, h_u_cla24_or175_y0);
  or_gate or_gate_h_u_cla24_or176_y0(h_u_cla24_or175_y0, h_u_cla24_and2300_y0, h_u_cla24_or176_y0);
  or_gate or_gate_h_u_cla24_or177_y0(h_u_cla24_or176_y0, h_u_cla24_and2325_y0, h_u_cla24_or177_y0);
  or_gate or_gate_h_u_cla24_or178_y0(h_u_cla24_or177_y0, h_u_cla24_and2348_y0, h_u_cla24_or178_y0);
  or_gate or_gate_h_u_cla24_or179_y0(h_u_cla24_or178_y0, h_u_cla24_and2369_y0, h_u_cla24_or179_y0);
  or_gate or_gate_h_u_cla24_or180_y0(h_u_cla24_or179_y0, h_u_cla24_and2388_y0, h_u_cla24_or180_y0);
  or_gate or_gate_h_u_cla24_or181_y0(h_u_cla24_or180_y0, h_u_cla24_and2405_y0, h_u_cla24_or181_y0);
  or_gate or_gate_h_u_cla24_or182_y0(h_u_cla24_or181_y0, h_u_cla24_and2420_y0, h_u_cla24_or182_y0);
  or_gate or_gate_h_u_cla24_or183_y0(h_u_cla24_or182_y0, h_u_cla24_and2433_y0, h_u_cla24_or183_y0);
  or_gate or_gate_h_u_cla24_or184_y0(h_u_cla24_or183_y0, h_u_cla24_and2444_y0, h_u_cla24_or184_y0);
  or_gate or_gate_h_u_cla24_or185_y0(h_u_cla24_or184_y0, h_u_cla24_and2453_y0, h_u_cla24_or185_y0);
  or_gate or_gate_h_u_cla24_or186_y0(h_u_cla24_or185_y0, h_u_cla24_and2460_y0, h_u_cla24_or186_y0);
  or_gate or_gate_h_u_cla24_or187_y0(h_u_cla24_or186_y0, h_u_cla24_and2465_y0, h_u_cla24_or187_y0);
  or_gate or_gate_h_u_cla24_or188_y0(h_u_cla24_or187_y0, h_u_cla24_and2468_y0, h_u_cla24_or188_y0);
  or_gate or_gate_h_u_cla24_or189_y0(h_u_cla24_pg_logic18_y1, h_u_cla24_or188_y0, h_u_cla24_or189_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic19_y0(a_19, b_19, h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_pg_logic19_y2);
  xor_gate xor_gate_h_u_cla24_xor19_y0(h_u_cla24_pg_logic19_y2, h_u_cla24_or189_y0, h_u_cla24_xor19_y0);
  and_gate and_gate_h_u_cla24_and2470_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and2470_y0);
  and_gate and_gate_h_u_cla24_and2471_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and2471_y0);
  and_gate and_gate_h_u_cla24_and2472_y0(h_u_cla24_and2471_y0, h_u_cla24_and2470_y0, h_u_cla24_and2472_y0);
  and_gate and_gate_h_u_cla24_and2473_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and2473_y0);
  and_gate and_gate_h_u_cla24_and2474_y0(h_u_cla24_and2473_y0, h_u_cla24_and2472_y0, h_u_cla24_and2474_y0);
  and_gate and_gate_h_u_cla24_and2475_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and2475_y0);
  and_gate and_gate_h_u_cla24_and2476_y0(h_u_cla24_and2475_y0, h_u_cla24_and2474_y0, h_u_cla24_and2476_y0);
  and_gate and_gate_h_u_cla24_and2477_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and2477_y0);
  and_gate and_gate_h_u_cla24_and2478_y0(h_u_cla24_and2477_y0, h_u_cla24_and2476_y0, h_u_cla24_and2478_y0);
  and_gate and_gate_h_u_cla24_and2479_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and2479_y0);
  and_gate and_gate_h_u_cla24_and2480_y0(h_u_cla24_and2479_y0, h_u_cla24_and2478_y0, h_u_cla24_and2480_y0);
  and_gate and_gate_h_u_cla24_and2481_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and2481_y0);
  and_gate and_gate_h_u_cla24_and2482_y0(h_u_cla24_and2481_y0, h_u_cla24_and2480_y0, h_u_cla24_and2482_y0);
  and_gate and_gate_h_u_cla24_and2483_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and2483_y0);
  and_gate and_gate_h_u_cla24_and2484_y0(h_u_cla24_and2483_y0, h_u_cla24_and2482_y0, h_u_cla24_and2484_y0);
  and_gate and_gate_h_u_cla24_and2485_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and2485_y0);
  and_gate and_gate_h_u_cla24_and2486_y0(h_u_cla24_and2485_y0, h_u_cla24_and2484_y0, h_u_cla24_and2486_y0);
  and_gate and_gate_h_u_cla24_and2487_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and2487_y0);
  and_gate and_gate_h_u_cla24_and2488_y0(h_u_cla24_and2487_y0, h_u_cla24_and2486_y0, h_u_cla24_and2488_y0);
  and_gate and_gate_h_u_cla24_and2489_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and2489_y0);
  and_gate and_gate_h_u_cla24_and2490_y0(h_u_cla24_and2489_y0, h_u_cla24_and2488_y0, h_u_cla24_and2490_y0);
  and_gate and_gate_h_u_cla24_and2491_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and2491_y0);
  and_gate and_gate_h_u_cla24_and2492_y0(h_u_cla24_and2491_y0, h_u_cla24_and2490_y0, h_u_cla24_and2492_y0);
  and_gate and_gate_h_u_cla24_and2493_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and2493_y0);
  and_gate and_gate_h_u_cla24_and2494_y0(h_u_cla24_and2493_y0, h_u_cla24_and2492_y0, h_u_cla24_and2494_y0);
  and_gate and_gate_h_u_cla24_and2495_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and2495_y0);
  and_gate and_gate_h_u_cla24_and2496_y0(h_u_cla24_and2495_y0, h_u_cla24_and2494_y0, h_u_cla24_and2496_y0);
  and_gate and_gate_h_u_cla24_and2497_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and2497_y0);
  and_gate and_gate_h_u_cla24_and2498_y0(h_u_cla24_and2497_y0, h_u_cla24_and2496_y0, h_u_cla24_and2498_y0);
  and_gate and_gate_h_u_cla24_and2499_y0(h_u_cla24_pg_logic15_y0, constant_wire_0, h_u_cla24_and2499_y0);
  and_gate and_gate_h_u_cla24_and2500_y0(h_u_cla24_and2499_y0, h_u_cla24_and2498_y0, h_u_cla24_and2500_y0);
  and_gate and_gate_h_u_cla24_and2501_y0(h_u_cla24_pg_logic16_y0, constant_wire_0, h_u_cla24_and2501_y0);
  and_gate and_gate_h_u_cla24_and2502_y0(h_u_cla24_and2501_y0, h_u_cla24_and2500_y0, h_u_cla24_and2502_y0);
  and_gate and_gate_h_u_cla24_and2503_y0(h_u_cla24_pg_logic17_y0, constant_wire_0, h_u_cla24_and2503_y0);
  and_gate and_gate_h_u_cla24_and2504_y0(h_u_cla24_and2503_y0, h_u_cla24_and2502_y0, h_u_cla24_and2504_y0);
  and_gate and_gate_h_u_cla24_and2505_y0(h_u_cla24_pg_logic18_y0, constant_wire_0, h_u_cla24_and2505_y0);
  and_gate and_gate_h_u_cla24_and2506_y0(h_u_cla24_and2505_y0, h_u_cla24_and2504_y0, h_u_cla24_and2506_y0);
  and_gate and_gate_h_u_cla24_and2507_y0(h_u_cla24_pg_logic19_y0, constant_wire_0, h_u_cla24_and2507_y0);
  and_gate and_gate_h_u_cla24_and2508_y0(h_u_cla24_and2507_y0, h_u_cla24_and2506_y0, h_u_cla24_and2508_y0);
  and_gate and_gate_h_u_cla24_and2509_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2509_y0);
  and_gate and_gate_h_u_cla24_and2510_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2510_y0);
  and_gate and_gate_h_u_cla24_and2511_y0(h_u_cla24_and2510_y0, h_u_cla24_and2509_y0, h_u_cla24_and2511_y0);
  and_gate and_gate_h_u_cla24_and2512_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2512_y0);
  and_gate and_gate_h_u_cla24_and2513_y0(h_u_cla24_and2512_y0, h_u_cla24_and2511_y0, h_u_cla24_and2513_y0);
  and_gate and_gate_h_u_cla24_and2514_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2514_y0);
  and_gate and_gate_h_u_cla24_and2515_y0(h_u_cla24_and2514_y0, h_u_cla24_and2513_y0, h_u_cla24_and2515_y0);
  and_gate and_gate_h_u_cla24_and2516_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2516_y0);
  and_gate and_gate_h_u_cla24_and2517_y0(h_u_cla24_and2516_y0, h_u_cla24_and2515_y0, h_u_cla24_and2517_y0);
  and_gate and_gate_h_u_cla24_and2518_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2518_y0);
  and_gate and_gate_h_u_cla24_and2519_y0(h_u_cla24_and2518_y0, h_u_cla24_and2517_y0, h_u_cla24_and2519_y0);
  and_gate and_gate_h_u_cla24_and2520_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2520_y0);
  and_gate and_gate_h_u_cla24_and2521_y0(h_u_cla24_and2520_y0, h_u_cla24_and2519_y0, h_u_cla24_and2521_y0);
  and_gate and_gate_h_u_cla24_and2522_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2522_y0);
  and_gate and_gate_h_u_cla24_and2523_y0(h_u_cla24_and2522_y0, h_u_cla24_and2521_y0, h_u_cla24_and2523_y0);
  and_gate and_gate_h_u_cla24_and2524_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2524_y0);
  and_gate and_gate_h_u_cla24_and2525_y0(h_u_cla24_and2524_y0, h_u_cla24_and2523_y0, h_u_cla24_and2525_y0);
  and_gate and_gate_h_u_cla24_and2526_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2526_y0);
  and_gate and_gate_h_u_cla24_and2527_y0(h_u_cla24_and2526_y0, h_u_cla24_and2525_y0, h_u_cla24_and2527_y0);
  and_gate and_gate_h_u_cla24_and2528_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2528_y0);
  and_gate and_gate_h_u_cla24_and2529_y0(h_u_cla24_and2528_y0, h_u_cla24_and2527_y0, h_u_cla24_and2529_y0);
  and_gate and_gate_h_u_cla24_and2530_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2530_y0);
  and_gate and_gate_h_u_cla24_and2531_y0(h_u_cla24_and2530_y0, h_u_cla24_and2529_y0, h_u_cla24_and2531_y0);
  and_gate and_gate_h_u_cla24_and2532_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2532_y0);
  and_gate and_gate_h_u_cla24_and2533_y0(h_u_cla24_and2532_y0, h_u_cla24_and2531_y0, h_u_cla24_and2533_y0);
  and_gate and_gate_h_u_cla24_and2534_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2534_y0);
  and_gate and_gate_h_u_cla24_and2535_y0(h_u_cla24_and2534_y0, h_u_cla24_and2533_y0, h_u_cla24_and2535_y0);
  and_gate and_gate_h_u_cla24_and2536_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2536_y0);
  and_gate and_gate_h_u_cla24_and2537_y0(h_u_cla24_and2536_y0, h_u_cla24_and2535_y0, h_u_cla24_and2537_y0);
  and_gate and_gate_h_u_cla24_and2538_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2538_y0);
  and_gate and_gate_h_u_cla24_and2539_y0(h_u_cla24_and2538_y0, h_u_cla24_and2537_y0, h_u_cla24_and2539_y0);
  and_gate and_gate_h_u_cla24_and2540_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2540_y0);
  and_gate and_gate_h_u_cla24_and2541_y0(h_u_cla24_and2540_y0, h_u_cla24_and2539_y0, h_u_cla24_and2541_y0);
  and_gate and_gate_h_u_cla24_and2542_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2542_y0);
  and_gate and_gate_h_u_cla24_and2543_y0(h_u_cla24_and2542_y0, h_u_cla24_and2541_y0, h_u_cla24_and2543_y0);
  and_gate and_gate_h_u_cla24_and2544_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2544_y0);
  and_gate and_gate_h_u_cla24_and2545_y0(h_u_cla24_and2544_y0, h_u_cla24_and2543_y0, h_u_cla24_and2545_y0);
  and_gate and_gate_h_u_cla24_and2546_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2546_y0);
  and_gate and_gate_h_u_cla24_and2547_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2547_y0);
  and_gate and_gate_h_u_cla24_and2548_y0(h_u_cla24_and2547_y0, h_u_cla24_and2546_y0, h_u_cla24_and2548_y0);
  and_gate and_gate_h_u_cla24_and2549_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2549_y0);
  and_gate and_gate_h_u_cla24_and2550_y0(h_u_cla24_and2549_y0, h_u_cla24_and2548_y0, h_u_cla24_and2550_y0);
  and_gate and_gate_h_u_cla24_and2551_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2551_y0);
  and_gate and_gate_h_u_cla24_and2552_y0(h_u_cla24_and2551_y0, h_u_cla24_and2550_y0, h_u_cla24_and2552_y0);
  and_gate and_gate_h_u_cla24_and2553_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2553_y0);
  and_gate and_gate_h_u_cla24_and2554_y0(h_u_cla24_and2553_y0, h_u_cla24_and2552_y0, h_u_cla24_and2554_y0);
  and_gate and_gate_h_u_cla24_and2555_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2555_y0);
  and_gate and_gate_h_u_cla24_and2556_y0(h_u_cla24_and2555_y0, h_u_cla24_and2554_y0, h_u_cla24_and2556_y0);
  and_gate and_gate_h_u_cla24_and2557_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2557_y0);
  and_gate and_gate_h_u_cla24_and2558_y0(h_u_cla24_and2557_y0, h_u_cla24_and2556_y0, h_u_cla24_and2558_y0);
  and_gate and_gate_h_u_cla24_and2559_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2559_y0);
  and_gate and_gate_h_u_cla24_and2560_y0(h_u_cla24_and2559_y0, h_u_cla24_and2558_y0, h_u_cla24_and2560_y0);
  and_gate and_gate_h_u_cla24_and2561_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2561_y0);
  and_gate and_gate_h_u_cla24_and2562_y0(h_u_cla24_and2561_y0, h_u_cla24_and2560_y0, h_u_cla24_and2562_y0);
  and_gate and_gate_h_u_cla24_and2563_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2563_y0);
  and_gate and_gate_h_u_cla24_and2564_y0(h_u_cla24_and2563_y0, h_u_cla24_and2562_y0, h_u_cla24_and2564_y0);
  and_gate and_gate_h_u_cla24_and2565_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2565_y0);
  and_gate and_gate_h_u_cla24_and2566_y0(h_u_cla24_and2565_y0, h_u_cla24_and2564_y0, h_u_cla24_and2566_y0);
  and_gate and_gate_h_u_cla24_and2567_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2567_y0);
  and_gate and_gate_h_u_cla24_and2568_y0(h_u_cla24_and2567_y0, h_u_cla24_and2566_y0, h_u_cla24_and2568_y0);
  and_gate and_gate_h_u_cla24_and2569_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2569_y0);
  and_gate and_gate_h_u_cla24_and2570_y0(h_u_cla24_and2569_y0, h_u_cla24_and2568_y0, h_u_cla24_and2570_y0);
  and_gate and_gate_h_u_cla24_and2571_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2571_y0);
  and_gate and_gate_h_u_cla24_and2572_y0(h_u_cla24_and2571_y0, h_u_cla24_and2570_y0, h_u_cla24_and2572_y0);
  and_gate and_gate_h_u_cla24_and2573_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2573_y0);
  and_gate and_gate_h_u_cla24_and2574_y0(h_u_cla24_and2573_y0, h_u_cla24_and2572_y0, h_u_cla24_and2574_y0);
  and_gate and_gate_h_u_cla24_and2575_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2575_y0);
  and_gate and_gate_h_u_cla24_and2576_y0(h_u_cla24_and2575_y0, h_u_cla24_and2574_y0, h_u_cla24_and2576_y0);
  and_gate and_gate_h_u_cla24_and2577_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2577_y0);
  and_gate and_gate_h_u_cla24_and2578_y0(h_u_cla24_and2577_y0, h_u_cla24_and2576_y0, h_u_cla24_and2578_y0);
  and_gate and_gate_h_u_cla24_and2579_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2579_y0);
  and_gate and_gate_h_u_cla24_and2580_y0(h_u_cla24_and2579_y0, h_u_cla24_and2578_y0, h_u_cla24_and2580_y0);
  and_gate and_gate_h_u_cla24_and2581_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2581_y0);
  and_gate and_gate_h_u_cla24_and2582_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2582_y0);
  and_gate and_gate_h_u_cla24_and2583_y0(h_u_cla24_and2582_y0, h_u_cla24_and2581_y0, h_u_cla24_and2583_y0);
  and_gate and_gate_h_u_cla24_and2584_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2584_y0);
  and_gate and_gate_h_u_cla24_and2585_y0(h_u_cla24_and2584_y0, h_u_cla24_and2583_y0, h_u_cla24_and2585_y0);
  and_gate and_gate_h_u_cla24_and2586_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2586_y0);
  and_gate and_gate_h_u_cla24_and2587_y0(h_u_cla24_and2586_y0, h_u_cla24_and2585_y0, h_u_cla24_and2587_y0);
  and_gate and_gate_h_u_cla24_and2588_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2588_y0);
  and_gate and_gate_h_u_cla24_and2589_y0(h_u_cla24_and2588_y0, h_u_cla24_and2587_y0, h_u_cla24_and2589_y0);
  and_gate and_gate_h_u_cla24_and2590_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2590_y0);
  and_gate and_gate_h_u_cla24_and2591_y0(h_u_cla24_and2590_y0, h_u_cla24_and2589_y0, h_u_cla24_and2591_y0);
  and_gate and_gate_h_u_cla24_and2592_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2592_y0);
  and_gate and_gate_h_u_cla24_and2593_y0(h_u_cla24_and2592_y0, h_u_cla24_and2591_y0, h_u_cla24_and2593_y0);
  and_gate and_gate_h_u_cla24_and2594_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2594_y0);
  and_gate and_gate_h_u_cla24_and2595_y0(h_u_cla24_and2594_y0, h_u_cla24_and2593_y0, h_u_cla24_and2595_y0);
  and_gate and_gate_h_u_cla24_and2596_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2596_y0);
  and_gate and_gate_h_u_cla24_and2597_y0(h_u_cla24_and2596_y0, h_u_cla24_and2595_y0, h_u_cla24_and2597_y0);
  and_gate and_gate_h_u_cla24_and2598_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2598_y0);
  and_gate and_gate_h_u_cla24_and2599_y0(h_u_cla24_and2598_y0, h_u_cla24_and2597_y0, h_u_cla24_and2599_y0);
  and_gate and_gate_h_u_cla24_and2600_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2600_y0);
  and_gate and_gate_h_u_cla24_and2601_y0(h_u_cla24_and2600_y0, h_u_cla24_and2599_y0, h_u_cla24_and2601_y0);
  and_gate and_gate_h_u_cla24_and2602_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2602_y0);
  and_gate and_gate_h_u_cla24_and2603_y0(h_u_cla24_and2602_y0, h_u_cla24_and2601_y0, h_u_cla24_and2603_y0);
  and_gate and_gate_h_u_cla24_and2604_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2604_y0);
  and_gate and_gate_h_u_cla24_and2605_y0(h_u_cla24_and2604_y0, h_u_cla24_and2603_y0, h_u_cla24_and2605_y0);
  and_gate and_gate_h_u_cla24_and2606_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2606_y0);
  and_gate and_gate_h_u_cla24_and2607_y0(h_u_cla24_and2606_y0, h_u_cla24_and2605_y0, h_u_cla24_and2607_y0);
  and_gate and_gate_h_u_cla24_and2608_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2608_y0);
  and_gate and_gate_h_u_cla24_and2609_y0(h_u_cla24_and2608_y0, h_u_cla24_and2607_y0, h_u_cla24_and2609_y0);
  and_gate and_gate_h_u_cla24_and2610_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2610_y0);
  and_gate and_gate_h_u_cla24_and2611_y0(h_u_cla24_and2610_y0, h_u_cla24_and2609_y0, h_u_cla24_and2611_y0);
  and_gate and_gate_h_u_cla24_and2612_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2612_y0);
  and_gate and_gate_h_u_cla24_and2613_y0(h_u_cla24_and2612_y0, h_u_cla24_and2611_y0, h_u_cla24_and2613_y0);
  and_gate and_gate_h_u_cla24_and2614_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2614_y0);
  and_gate and_gate_h_u_cla24_and2615_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2615_y0);
  and_gate and_gate_h_u_cla24_and2616_y0(h_u_cla24_and2615_y0, h_u_cla24_and2614_y0, h_u_cla24_and2616_y0);
  and_gate and_gate_h_u_cla24_and2617_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2617_y0);
  and_gate and_gate_h_u_cla24_and2618_y0(h_u_cla24_and2617_y0, h_u_cla24_and2616_y0, h_u_cla24_and2618_y0);
  and_gate and_gate_h_u_cla24_and2619_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2619_y0);
  and_gate and_gate_h_u_cla24_and2620_y0(h_u_cla24_and2619_y0, h_u_cla24_and2618_y0, h_u_cla24_and2620_y0);
  and_gate and_gate_h_u_cla24_and2621_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2621_y0);
  and_gate and_gate_h_u_cla24_and2622_y0(h_u_cla24_and2621_y0, h_u_cla24_and2620_y0, h_u_cla24_and2622_y0);
  and_gate and_gate_h_u_cla24_and2623_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2623_y0);
  and_gate and_gate_h_u_cla24_and2624_y0(h_u_cla24_and2623_y0, h_u_cla24_and2622_y0, h_u_cla24_and2624_y0);
  and_gate and_gate_h_u_cla24_and2625_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2625_y0);
  and_gate and_gate_h_u_cla24_and2626_y0(h_u_cla24_and2625_y0, h_u_cla24_and2624_y0, h_u_cla24_and2626_y0);
  and_gate and_gate_h_u_cla24_and2627_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2627_y0);
  and_gate and_gate_h_u_cla24_and2628_y0(h_u_cla24_and2627_y0, h_u_cla24_and2626_y0, h_u_cla24_and2628_y0);
  and_gate and_gate_h_u_cla24_and2629_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2629_y0);
  and_gate and_gate_h_u_cla24_and2630_y0(h_u_cla24_and2629_y0, h_u_cla24_and2628_y0, h_u_cla24_and2630_y0);
  and_gate and_gate_h_u_cla24_and2631_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2631_y0);
  and_gate and_gate_h_u_cla24_and2632_y0(h_u_cla24_and2631_y0, h_u_cla24_and2630_y0, h_u_cla24_and2632_y0);
  and_gate and_gate_h_u_cla24_and2633_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2633_y0);
  and_gate and_gate_h_u_cla24_and2634_y0(h_u_cla24_and2633_y0, h_u_cla24_and2632_y0, h_u_cla24_and2634_y0);
  and_gate and_gate_h_u_cla24_and2635_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2635_y0);
  and_gate and_gate_h_u_cla24_and2636_y0(h_u_cla24_and2635_y0, h_u_cla24_and2634_y0, h_u_cla24_and2636_y0);
  and_gate and_gate_h_u_cla24_and2637_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2637_y0);
  and_gate and_gate_h_u_cla24_and2638_y0(h_u_cla24_and2637_y0, h_u_cla24_and2636_y0, h_u_cla24_and2638_y0);
  and_gate and_gate_h_u_cla24_and2639_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2639_y0);
  and_gate and_gate_h_u_cla24_and2640_y0(h_u_cla24_and2639_y0, h_u_cla24_and2638_y0, h_u_cla24_and2640_y0);
  and_gate and_gate_h_u_cla24_and2641_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2641_y0);
  and_gate and_gate_h_u_cla24_and2642_y0(h_u_cla24_and2641_y0, h_u_cla24_and2640_y0, h_u_cla24_and2642_y0);
  and_gate and_gate_h_u_cla24_and2643_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and2643_y0);
  and_gate and_gate_h_u_cla24_and2644_y0(h_u_cla24_and2643_y0, h_u_cla24_and2642_y0, h_u_cla24_and2644_y0);
  and_gate and_gate_h_u_cla24_and2645_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2645_y0);
  and_gate and_gate_h_u_cla24_and2646_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2646_y0);
  and_gate and_gate_h_u_cla24_and2647_y0(h_u_cla24_and2646_y0, h_u_cla24_and2645_y0, h_u_cla24_and2647_y0);
  and_gate and_gate_h_u_cla24_and2648_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2648_y0);
  and_gate and_gate_h_u_cla24_and2649_y0(h_u_cla24_and2648_y0, h_u_cla24_and2647_y0, h_u_cla24_and2649_y0);
  and_gate and_gate_h_u_cla24_and2650_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2650_y0);
  and_gate and_gate_h_u_cla24_and2651_y0(h_u_cla24_and2650_y0, h_u_cla24_and2649_y0, h_u_cla24_and2651_y0);
  and_gate and_gate_h_u_cla24_and2652_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2652_y0);
  and_gate and_gate_h_u_cla24_and2653_y0(h_u_cla24_and2652_y0, h_u_cla24_and2651_y0, h_u_cla24_and2653_y0);
  and_gate and_gate_h_u_cla24_and2654_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2654_y0);
  and_gate and_gate_h_u_cla24_and2655_y0(h_u_cla24_and2654_y0, h_u_cla24_and2653_y0, h_u_cla24_and2655_y0);
  and_gate and_gate_h_u_cla24_and2656_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2656_y0);
  and_gate and_gate_h_u_cla24_and2657_y0(h_u_cla24_and2656_y0, h_u_cla24_and2655_y0, h_u_cla24_and2657_y0);
  and_gate and_gate_h_u_cla24_and2658_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2658_y0);
  and_gate and_gate_h_u_cla24_and2659_y0(h_u_cla24_and2658_y0, h_u_cla24_and2657_y0, h_u_cla24_and2659_y0);
  and_gate and_gate_h_u_cla24_and2660_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2660_y0);
  and_gate and_gate_h_u_cla24_and2661_y0(h_u_cla24_and2660_y0, h_u_cla24_and2659_y0, h_u_cla24_and2661_y0);
  and_gate and_gate_h_u_cla24_and2662_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2662_y0);
  and_gate and_gate_h_u_cla24_and2663_y0(h_u_cla24_and2662_y0, h_u_cla24_and2661_y0, h_u_cla24_and2663_y0);
  and_gate and_gate_h_u_cla24_and2664_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2664_y0);
  and_gate and_gate_h_u_cla24_and2665_y0(h_u_cla24_and2664_y0, h_u_cla24_and2663_y0, h_u_cla24_and2665_y0);
  and_gate and_gate_h_u_cla24_and2666_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2666_y0);
  and_gate and_gate_h_u_cla24_and2667_y0(h_u_cla24_and2666_y0, h_u_cla24_and2665_y0, h_u_cla24_and2667_y0);
  and_gate and_gate_h_u_cla24_and2668_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2668_y0);
  and_gate and_gate_h_u_cla24_and2669_y0(h_u_cla24_and2668_y0, h_u_cla24_and2667_y0, h_u_cla24_and2669_y0);
  and_gate and_gate_h_u_cla24_and2670_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2670_y0);
  and_gate and_gate_h_u_cla24_and2671_y0(h_u_cla24_and2670_y0, h_u_cla24_and2669_y0, h_u_cla24_and2671_y0);
  and_gate and_gate_h_u_cla24_and2672_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and2672_y0);
  and_gate and_gate_h_u_cla24_and2673_y0(h_u_cla24_and2672_y0, h_u_cla24_and2671_y0, h_u_cla24_and2673_y0);
  and_gate and_gate_h_u_cla24_and2674_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2674_y0);
  and_gate and_gate_h_u_cla24_and2675_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2675_y0);
  and_gate and_gate_h_u_cla24_and2676_y0(h_u_cla24_and2675_y0, h_u_cla24_and2674_y0, h_u_cla24_and2676_y0);
  and_gate and_gate_h_u_cla24_and2677_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2677_y0);
  and_gate and_gate_h_u_cla24_and2678_y0(h_u_cla24_and2677_y0, h_u_cla24_and2676_y0, h_u_cla24_and2678_y0);
  and_gate and_gate_h_u_cla24_and2679_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2679_y0);
  and_gate and_gate_h_u_cla24_and2680_y0(h_u_cla24_and2679_y0, h_u_cla24_and2678_y0, h_u_cla24_and2680_y0);
  and_gate and_gate_h_u_cla24_and2681_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2681_y0);
  and_gate and_gate_h_u_cla24_and2682_y0(h_u_cla24_and2681_y0, h_u_cla24_and2680_y0, h_u_cla24_and2682_y0);
  and_gate and_gate_h_u_cla24_and2683_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2683_y0);
  and_gate and_gate_h_u_cla24_and2684_y0(h_u_cla24_and2683_y0, h_u_cla24_and2682_y0, h_u_cla24_and2684_y0);
  and_gate and_gate_h_u_cla24_and2685_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2685_y0);
  and_gate and_gate_h_u_cla24_and2686_y0(h_u_cla24_and2685_y0, h_u_cla24_and2684_y0, h_u_cla24_and2686_y0);
  and_gate and_gate_h_u_cla24_and2687_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2687_y0);
  and_gate and_gate_h_u_cla24_and2688_y0(h_u_cla24_and2687_y0, h_u_cla24_and2686_y0, h_u_cla24_and2688_y0);
  and_gate and_gate_h_u_cla24_and2689_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2689_y0);
  and_gate and_gate_h_u_cla24_and2690_y0(h_u_cla24_and2689_y0, h_u_cla24_and2688_y0, h_u_cla24_and2690_y0);
  and_gate and_gate_h_u_cla24_and2691_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2691_y0);
  and_gate and_gate_h_u_cla24_and2692_y0(h_u_cla24_and2691_y0, h_u_cla24_and2690_y0, h_u_cla24_and2692_y0);
  and_gate and_gate_h_u_cla24_and2693_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2693_y0);
  and_gate and_gate_h_u_cla24_and2694_y0(h_u_cla24_and2693_y0, h_u_cla24_and2692_y0, h_u_cla24_and2694_y0);
  and_gate and_gate_h_u_cla24_and2695_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2695_y0);
  and_gate and_gate_h_u_cla24_and2696_y0(h_u_cla24_and2695_y0, h_u_cla24_and2694_y0, h_u_cla24_and2696_y0);
  and_gate and_gate_h_u_cla24_and2697_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2697_y0);
  and_gate and_gate_h_u_cla24_and2698_y0(h_u_cla24_and2697_y0, h_u_cla24_and2696_y0, h_u_cla24_and2698_y0);
  and_gate and_gate_h_u_cla24_and2699_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and2699_y0);
  and_gate and_gate_h_u_cla24_and2700_y0(h_u_cla24_and2699_y0, h_u_cla24_and2698_y0, h_u_cla24_and2700_y0);
  and_gate and_gate_h_u_cla24_and2701_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2701_y0);
  and_gate and_gate_h_u_cla24_and2702_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2702_y0);
  and_gate and_gate_h_u_cla24_and2703_y0(h_u_cla24_and2702_y0, h_u_cla24_and2701_y0, h_u_cla24_and2703_y0);
  and_gate and_gate_h_u_cla24_and2704_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2704_y0);
  and_gate and_gate_h_u_cla24_and2705_y0(h_u_cla24_and2704_y0, h_u_cla24_and2703_y0, h_u_cla24_and2705_y0);
  and_gate and_gate_h_u_cla24_and2706_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2706_y0);
  and_gate and_gate_h_u_cla24_and2707_y0(h_u_cla24_and2706_y0, h_u_cla24_and2705_y0, h_u_cla24_and2707_y0);
  and_gate and_gate_h_u_cla24_and2708_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2708_y0);
  and_gate and_gate_h_u_cla24_and2709_y0(h_u_cla24_and2708_y0, h_u_cla24_and2707_y0, h_u_cla24_and2709_y0);
  and_gate and_gate_h_u_cla24_and2710_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2710_y0);
  and_gate and_gate_h_u_cla24_and2711_y0(h_u_cla24_and2710_y0, h_u_cla24_and2709_y0, h_u_cla24_and2711_y0);
  and_gate and_gate_h_u_cla24_and2712_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2712_y0);
  and_gate and_gate_h_u_cla24_and2713_y0(h_u_cla24_and2712_y0, h_u_cla24_and2711_y0, h_u_cla24_and2713_y0);
  and_gate and_gate_h_u_cla24_and2714_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2714_y0);
  and_gate and_gate_h_u_cla24_and2715_y0(h_u_cla24_and2714_y0, h_u_cla24_and2713_y0, h_u_cla24_and2715_y0);
  and_gate and_gate_h_u_cla24_and2716_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2716_y0);
  and_gate and_gate_h_u_cla24_and2717_y0(h_u_cla24_and2716_y0, h_u_cla24_and2715_y0, h_u_cla24_and2717_y0);
  and_gate and_gate_h_u_cla24_and2718_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2718_y0);
  and_gate and_gate_h_u_cla24_and2719_y0(h_u_cla24_and2718_y0, h_u_cla24_and2717_y0, h_u_cla24_and2719_y0);
  and_gate and_gate_h_u_cla24_and2720_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2720_y0);
  and_gate and_gate_h_u_cla24_and2721_y0(h_u_cla24_and2720_y0, h_u_cla24_and2719_y0, h_u_cla24_and2721_y0);
  and_gate and_gate_h_u_cla24_and2722_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2722_y0);
  and_gate and_gate_h_u_cla24_and2723_y0(h_u_cla24_and2722_y0, h_u_cla24_and2721_y0, h_u_cla24_and2723_y0);
  and_gate and_gate_h_u_cla24_and2724_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and2724_y0);
  and_gate and_gate_h_u_cla24_and2725_y0(h_u_cla24_and2724_y0, h_u_cla24_and2723_y0, h_u_cla24_and2725_y0);
  and_gate and_gate_h_u_cla24_and2726_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2726_y0);
  and_gate and_gate_h_u_cla24_and2727_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2727_y0);
  and_gate and_gate_h_u_cla24_and2728_y0(h_u_cla24_and2727_y0, h_u_cla24_and2726_y0, h_u_cla24_and2728_y0);
  and_gate and_gate_h_u_cla24_and2729_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2729_y0);
  and_gate and_gate_h_u_cla24_and2730_y0(h_u_cla24_and2729_y0, h_u_cla24_and2728_y0, h_u_cla24_and2730_y0);
  and_gate and_gate_h_u_cla24_and2731_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2731_y0);
  and_gate and_gate_h_u_cla24_and2732_y0(h_u_cla24_and2731_y0, h_u_cla24_and2730_y0, h_u_cla24_and2732_y0);
  and_gate and_gate_h_u_cla24_and2733_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2733_y0);
  and_gate and_gate_h_u_cla24_and2734_y0(h_u_cla24_and2733_y0, h_u_cla24_and2732_y0, h_u_cla24_and2734_y0);
  and_gate and_gate_h_u_cla24_and2735_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2735_y0);
  and_gate and_gate_h_u_cla24_and2736_y0(h_u_cla24_and2735_y0, h_u_cla24_and2734_y0, h_u_cla24_and2736_y0);
  and_gate and_gate_h_u_cla24_and2737_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2737_y0);
  and_gate and_gate_h_u_cla24_and2738_y0(h_u_cla24_and2737_y0, h_u_cla24_and2736_y0, h_u_cla24_and2738_y0);
  and_gate and_gate_h_u_cla24_and2739_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2739_y0);
  and_gate and_gate_h_u_cla24_and2740_y0(h_u_cla24_and2739_y0, h_u_cla24_and2738_y0, h_u_cla24_and2740_y0);
  and_gate and_gate_h_u_cla24_and2741_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2741_y0);
  and_gate and_gate_h_u_cla24_and2742_y0(h_u_cla24_and2741_y0, h_u_cla24_and2740_y0, h_u_cla24_and2742_y0);
  and_gate and_gate_h_u_cla24_and2743_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2743_y0);
  and_gate and_gate_h_u_cla24_and2744_y0(h_u_cla24_and2743_y0, h_u_cla24_and2742_y0, h_u_cla24_and2744_y0);
  and_gate and_gate_h_u_cla24_and2745_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2745_y0);
  and_gate and_gate_h_u_cla24_and2746_y0(h_u_cla24_and2745_y0, h_u_cla24_and2744_y0, h_u_cla24_and2746_y0);
  and_gate and_gate_h_u_cla24_and2747_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and2747_y0);
  and_gate and_gate_h_u_cla24_and2748_y0(h_u_cla24_and2747_y0, h_u_cla24_and2746_y0, h_u_cla24_and2748_y0);
  and_gate and_gate_h_u_cla24_and2749_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2749_y0);
  and_gate and_gate_h_u_cla24_and2750_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2750_y0);
  and_gate and_gate_h_u_cla24_and2751_y0(h_u_cla24_and2750_y0, h_u_cla24_and2749_y0, h_u_cla24_and2751_y0);
  and_gate and_gate_h_u_cla24_and2752_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2752_y0);
  and_gate and_gate_h_u_cla24_and2753_y0(h_u_cla24_and2752_y0, h_u_cla24_and2751_y0, h_u_cla24_and2753_y0);
  and_gate and_gate_h_u_cla24_and2754_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2754_y0);
  and_gate and_gate_h_u_cla24_and2755_y0(h_u_cla24_and2754_y0, h_u_cla24_and2753_y0, h_u_cla24_and2755_y0);
  and_gate and_gate_h_u_cla24_and2756_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2756_y0);
  and_gate and_gate_h_u_cla24_and2757_y0(h_u_cla24_and2756_y0, h_u_cla24_and2755_y0, h_u_cla24_and2757_y0);
  and_gate and_gate_h_u_cla24_and2758_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2758_y0);
  and_gate and_gate_h_u_cla24_and2759_y0(h_u_cla24_and2758_y0, h_u_cla24_and2757_y0, h_u_cla24_and2759_y0);
  and_gate and_gate_h_u_cla24_and2760_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2760_y0);
  and_gate and_gate_h_u_cla24_and2761_y0(h_u_cla24_and2760_y0, h_u_cla24_and2759_y0, h_u_cla24_and2761_y0);
  and_gate and_gate_h_u_cla24_and2762_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2762_y0);
  and_gate and_gate_h_u_cla24_and2763_y0(h_u_cla24_and2762_y0, h_u_cla24_and2761_y0, h_u_cla24_and2763_y0);
  and_gate and_gate_h_u_cla24_and2764_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2764_y0);
  and_gate and_gate_h_u_cla24_and2765_y0(h_u_cla24_and2764_y0, h_u_cla24_and2763_y0, h_u_cla24_and2765_y0);
  and_gate and_gate_h_u_cla24_and2766_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2766_y0);
  and_gate and_gate_h_u_cla24_and2767_y0(h_u_cla24_and2766_y0, h_u_cla24_and2765_y0, h_u_cla24_and2767_y0);
  and_gate and_gate_h_u_cla24_and2768_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and2768_y0);
  and_gate and_gate_h_u_cla24_and2769_y0(h_u_cla24_and2768_y0, h_u_cla24_and2767_y0, h_u_cla24_and2769_y0);
  and_gate and_gate_h_u_cla24_and2770_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2770_y0);
  and_gate and_gate_h_u_cla24_and2771_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2771_y0);
  and_gate and_gate_h_u_cla24_and2772_y0(h_u_cla24_and2771_y0, h_u_cla24_and2770_y0, h_u_cla24_and2772_y0);
  and_gate and_gate_h_u_cla24_and2773_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2773_y0);
  and_gate and_gate_h_u_cla24_and2774_y0(h_u_cla24_and2773_y0, h_u_cla24_and2772_y0, h_u_cla24_and2774_y0);
  and_gate and_gate_h_u_cla24_and2775_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2775_y0);
  and_gate and_gate_h_u_cla24_and2776_y0(h_u_cla24_and2775_y0, h_u_cla24_and2774_y0, h_u_cla24_and2776_y0);
  and_gate and_gate_h_u_cla24_and2777_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2777_y0);
  and_gate and_gate_h_u_cla24_and2778_y0(h_u_cla24_and2777_y0, h_u_cla24_and2776_y0, h_u_cla24_and2778_y0);
  and_gate and_gate_h_u_cla24_and2779_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2779_y0);
  and_gate and_gate_h_u_cla24_and2780_y0(h_u_cla24_and2779_y0, h_u_cla24_and2778_y0, h_u_cla24_and2780_y0);
  and_gate and_gate_h_u_cla24_and2781_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2781_y0);
  and_gate and_gate_h_u_cla24_and2782_y0(h_u_cla24_and2781_y0, h_u_cla24_and2780_y0, h_u_cla24_and2782_y0);
  and_gate and_gate_h_u_cla24_and2783_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2783_y0);
  and_gate and_gate_h_u_cla24_and2784_y0(h_u_cla24_and2783_y0, h_u_cla24_and2782_y0, h_u_cla24_and2784_y0);
  and_gate and_gate_h_u_cla24_and2785_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2785_y0);
  and_gate and_gate_h_u_cla24_and2786_y0(h_u_cla24_and2785_y0, h_u_cla24_and2784_y0, h_u_cla24_and2786_y0);
  and_gate and_gate_h_u_cla24_and2787_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and2787_y0);
  and_gate and_gate_h_u_cla24_and2788_y0(h_u_cla24_and2787_y0, h_u_cla24_and2786_y0, h_u_cla24_and2788_y0);
  and_gate and_gate_h_u_cla24_and2789_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2789_y0);
  and_gate and_gate_h_u_cla24_and2790_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2790_y0);
  and_gate and_gate_h_u_cla24_and2791_y0(h_u_cla24_and2790_y0, h_u_cla24_and2789_y0, h_u_cla24_and2791_y0);
  and_gate and_gate_h_u_cla24_and2792_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2792_y0);
  and_gate and_gate_h_u_cla24_and2793_y0(h_u_cla24_and2792_y0, h_u_cla24_and2791_y0, h_u_cla24_and2793_y0);
  and_gate and_gate_h_u_cla24_and2794_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2794_y0);
  and_gate and_gate_h_u_cla24_and2795_y0(h_u_cla24_and2794_y0, h_u_cla24_and2793_y0, h_u_cla24_and2795_y0);
  and_gate and_gate_h_u_cla24_and2796_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2796_y0);
  and_gate and_gate_h_u_cla24_and2797_y0(h_u_cla24_and2796_y0, h_u_cla24_and2795_y0, h_u_cla24_and2797_y0);
  and_gate and_gate_h_u_cla24_and2798_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2798_y0);
  and_gate and_gate_h_u_cla24_and2799_y0(h_u_cla24_and2798_y0, h_u_cla24_and2797_y0, h_u_cla24_and2799_y0);
  and_gate and_gate_h_u_cla24_and2800_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2800_y0);
  and_gate and_gate_h_u_cla24_and2801_y0(h_u_cla24_and2800_y0, h_u_cla24_and2799_y0, h_u_cla24_and2801_y0);
  and_gate and_gate_h_u_cla24_and2802_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2802_y0);
  and_gate and_gate_h_u_cla24_and2803_y0(h_u_cla24_and2802_y0, h_u_cla24_and2801_y0, h_u_cla24_and2803_y0);
  and_gate and_gate_h_u_cla24_and2804_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and2804_y0);
  and_gate and_gate_h_u_cla24_and2805_y0(h_u_cla24_and2804_y0, h_u_cla24_and2803_y0, h_u_cla24_and2805_y0);
  and_gate and_gate_h_u_cla24_and2806_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2806_y0);
  and_gate and_gate_h_u_cla24_and2807_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2807_y0);
  and_gate and_gate_h_u_cla24_and2808_y0(h_u_cla24_and2807_y0, h_u_cla24_and2806_y0, h_u_cla24_and2808_y0);
  and_gate and_gate_h_u_cla24_and2809_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2809_y0);
  and_gate and_gate_h_u_cla24_and2810_y0(h_u_cla24_and2809_y0, h_u_cla24_and2808_y0, h_u_cla24_and2810_y0);
  and_gate and_gate_h_u_cla24_and2811_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2811_y0);
  and_gate and_gate_h_u_cla24_and2812_y0(h_u_cla24_and2811_y0, h_u_cla24_and2810_y0, h_u_cla24_and2812_y0);
  and_gate and_gate_h_u_cla24_and2813_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2813_y0);
  and_gate and_gate_h_u_cla24_and2814_y0(h_u_cla24_and2813_y0, h_u_cla24_and2812_y0, h_u_cla24_and2814_y0);
  and_gate and_gate_h_u_cla24_and2815_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2815_y0);
  and_gate and_gate_h_u_cla24_and2816_y0(h_u_cla24_and2815_y0, h_u_cla24_and2814_y0, h_u_cla24_and2816_y0);
  and_gate and_gate_h_u_cla24_and2817_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2817_y0);
  and_gate and_gate_h_u_cla24_and2818_y0(h_u_cla24_and2817_y0, h_u_cla24_and2816_y0, h_u_cla24_and2818_y0);
  and_gate and_gate_h_u_cla24_and2819_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and2819_y0);
  and_gate and_gate_h_u_cla24_and2820_y0(h_u_cla24_and2819_y0, h_u_cla24_and2818_y0, h_u_cla24_and2820_y0);
  and_gate and_gate_h_u_cla24_and2821_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2821_y0);
  and_gate and_gate_h_u_cla24_and2822_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2822_y0);
  and_gate and_gate_h_u_cla24_and2823_y0(h_u_cla24_and2822_y0, h_u_cla24_and2821_y0, h_u_cla24_and2823_y0);
  and_gate and_gate_h_u_cla24_and2824_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2824_y0);
  and_gate and_gate_h_u_cla24_and2825_y0(h_u_cla24_and2824_y0, h_u_cla24_and2823_y0, h_u_cla24_and2825_y0);
  and_gate and_gate_h_u_cla24_and2826_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2826_y0);
  and_gate and_gate_h_u_cla24_and2827_y0(h_u_cla24_and2826_y0, h_u_cla24_and2825_y0, h_u_cla24_and2827_y0);
  and_gate and_gate_h_u_cla24_and2828_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2828_y0);
  and_gate and_gate_h_u_cla24_and2829_y0(h_u_cla24_and2828_y0, h_u_cla24_and2827_y0, h_u_cla24_and2829_y0);
  and_gate and_gate_h_u_cla24_and2830_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2830_y0);
  and_gate and_gate_h_u_cla24_and2831_y0(h_u_cla24_and2830_y0, h_u_cla24_and2829_y0, h_u_cla24_and2831_y0);
  and_gate and_gate_h_u_cla24_and2832_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and2832_y0);
  and_gate and_gate_h_u_cla24_and2833_y0(h_u_cla24_and2832_y0, h_u_cla24_and2831_y0, h_u_cla24_and2833_y0);
  and_gate and_gate_h_u_cla24_and2834_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2834_y0);
  and_gate and_gate_h_u_cla24_and2835_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2835_y0);
  and_gate and_gate_h_u_cla24_and2836_y0(h_u_cla24_and2835_y0, h_u_cla24_and2834_y0, h_u_cla24_and2836_y0);
  and_gate and_gate_h_u_cla24_and2837_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2837_y0);
  and_gate and_gate_h_u_cla24_and2838_y0(h_u_cla24_and2837_y0, h_u_cla24_and2836_y0, h_u_cla24_and2838_y0);
  and_gate and_gate_h_u_cla24_and2839_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2839_y0);
  and_gate and_gate_h_u_cla24_and2840_y0(h_u_cla24_and2839_y0, h_u_cla24_and2838_y0, h_u_cla24_and2840_y0);
  and_gate and_gate_h_u_cla24_and2841_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2841_y0);
  and_gate and_gate_h_u_cla24_and2842_y0(h_u_cla24_and2841_y0, h_u_cla24_and2840_y0, h_u_cla24_and2842_y0);
  and_gate and_gate_h_u_cla24_and2843_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and2843_y0);
  and_gate and_gate_h_u_cla24_and2844_y0(h_u_cla24_and2843_y0, h_u_cla24_and2842_y0, h_u_cla24_and2844_y0);
  and_gate and_gate_h_u_cla24_and2845_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2845_y0);
  and_gate and_gate_h_u_cla24_and2846_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2846_y0);
  and_gate and_gate_h_u_cla24_and2847_y0(h_u_cla24_and2846_y0, h_u_cla24_and2845_y0, h_u_cla24_and2847_y0);
  and_gate and_gate_h_u_cla24_and2848_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2848_y0);
  and_gate and_gate_h_u_cla24_and2849_y0(h_u_cla24_and2848_y0, h_u_cla24_and2847_y0, h_u_cla24_and2849_y0);
  and_gate and_gate_h_u_cla24_and2850_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2850_y0);
  and_gate and_gate_h_u_cla24_and2851_y0(h_u_cla24_and2850_y0, h_u_cla24_and2849_y0, h_u_cla24_and2851_y0);
  and_gate and_gate_h_u_cla24_and2852_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and2852_y0);
  and_gate and_gate_h_u_cla24_and2853_y0(h_u_cla24_and2852_y0, h_u_cla24_and2851_y0, h_u_cla24_and2853_y0);
  and_gate and_gate_h_u_cla24_and2854_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and2854_y0);
  and_gate and_gate_h_u_cla24_and2855_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and2855_y0);
  and_gate and_gate_h_u_cla24_and2856_y0(h_u_cla24_and2855_y0, h_u_cla24_and2854_y0, h_u_cla24_and2856_y0);
  and_gate and_gate_h_u_cla24_and2857_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and2857_y0);
  and_gate and_gate_h_u_cla24_and2858_y0(h_u_cla24_and2857_y0, h_u_cla24_and2856_y0, h_u_cla24_and2858_y0);
  and_gate and_gate_h_u_cla24_and2859_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and2859_y0);
  and_gate and_gate_h_u_cla24_and2860_y0(h_u_cla24_and2859_y0, h_u_cla24_and2858_y0, h_u_cla24_and2860_y0);
  and_gate and_gate_h_u_cla24_and2861_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and2861_y0);
  and_gate and_gate_h_u_cla24_and2862_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and2862_y0);
  and_gate and_gate_h_u_cla24_and2863_y0(h_u_cla24_and2862_y0, h_u_cla24_and2861_y0, h_u_cla24_and2863_y0);
  and_gate and_gate_h_u_cla24_and2864_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and2864_y0);
  and_gate and_gate_h_u_cla24_and2865_y0(h_u_cla24_and2864_y0, h_u_cla24_and2863_y0, h_u_cla24_and2865_y0);
  and_gate and_gate_h_u_cla24_and2866_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and2866_y0);
  and_gate and_gate_h_u_cla24_and2867_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and2867_y0);
  and_gate and_gate_h_u_cla24_and2868_y0(h_u_cla24_and2867_y0, h_u_cla24_and2866_y0, h_u_cla24_and2868_y0);
  and_gate and_gate_h_u_cla24_and2869_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and2869_y0);
  or_gate or_gate_h_u_cla24_or190_y0(h_u_cla24_and2869_y0, h_u_cla24_and2508_y0, h_u_cla24_or190_y0);
  or_gate or_gate_h_u_cla24_or191_y0(h_u_cla24_or190_y0, h_u_cla24_and2545_y0, h_u_cla24_or191_y0);
  or_gate or_gate_h_u_cla24_or192_y0(h_u_cla24_or191_y0, h_u_cla24_and2580_y0, h_u_cla24_or192_y0);
  or_gate or_gate_h_u_cla24_or193_y0(h_u_cla24_or192_y0, h_u_cla24_and2613_y0, h_u_cla24_or193_y0);
  or_gate or_gate_h_u_cla24_or194_y0(h_u_cla24_or193_y0, h_u_cla24_and2644_y0, h_u_cla24_or194_y0);
  or_gate or_gate_h_u_cla24_or195_y0(h_u_cla24_or194_y0, h_u_cla24_and2673_y0, h_u_cla24_or195_y0);
  or_gate or_gate_h_u_cla24_or196_y0(h_u_cla24_or195_y0, h_u_cla24_and2700_y0, h_u_cla24_or196_y0);
  or_gate or_gate_h_u_cla24_or197_y0(h_u_cla24_or196_y0, h_u_cla24_and2725_y0, h_u_cla24_or197_y0);
  or_gate or_gate_h_u_cla24_or198_y0(h_u_cla24_or197_y0, h_u_cla24_and2748_y0, h_u_cla24_or198_y0);
  or_gate or_gate_h_u_cla24_or199_y0(h_u_cla24_or198_y0, h_u_cla24_and2769_y0, h_u_cla24_or199_y0);
  or_gate or_gate_h_u_cla24_or200_y0(h_u_cla24_or199_y0, h_u_cla24_and2788_y0, h_u_cla24_or200_y0);
  or_gate or_gate_h_u_cla24_or201_y0(h_u_cla24_or200_y0, h_u_cla24_and2805_y0, h_u_cla24_or201_y0);
  or_gate or_gate_h_u_cla24_or202_y0(h_u_cla24_or201_y0, h_u_cla24_and2820_y0, h_u_cla24_or202_y0);
  or_gate or_gate_h_u_cla24_or203_y0(h_u_cla24_or202_y0, h_u_cla24_and2833_y0, h_u_cla24_or203_y0);
  or_gate or_gate_h_u_cla24_or204_y0(h_u_cla24_or203_y0, h_u_cla24_and2844_y0, h_u_cla24_or204_y0);
  or_gate or_gate_h_u_cla24_or205_y0(h_u_cla24_or204_y0, h_u_cla24_and2853_y0, h_u_cla24_or205_y0);
  or_gate or_gate_h_u_cla24_or206_y0(h_u_cla24_or205_y0, h_u_cla24_and2860_y0, h_u_cla24_or206_y0);
  or_gate or_gate_h_u_cla24_or207_y0(h_u_cla24_or206_y0, h_u_cla24_and2865_y0, h_u_cla24_or207_y0);
  or_gate or_gate_h_u_cla24_or208_y0(h_u_cla24_or207_y0, h_u_cla24_and2868_y0, h_u_cla24_or208_y0);
  or_gate or_gate_h_u_cla24_or209_y0(h_u_cla24_pg_logic19_y1, h_u_cla24_or208_y0, h_u_cla24_or209_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic20_y0(a_20, b_20, h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic20_y1, h_u_cla24_pg_logic20_y2);
  xor_gate xor_gate_h_u_cla24_xor20_y0(h_u_cla24_pg_logic20_y2, h_u_cla24_or209_y0, h_u_cla24_xor20_y0);
  and_gate and_gate_h_u_cla24_and2870_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and2870_y0);
  and_gate and_gate_h_u_cla24_and2871_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and2871_y0);
  and_gate and_gate_h_u_cla24_and2872_y0(h_u_cla24_and2871_y0, h_u_cla24_and2870_y0, h_u_cla24_and2872_y0);
  and_gate and_gate_h_u_cla24_and2873_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and2873_y0);
  and_gate and_gate_h_u_cla24_and2874_y0(h_u_cla24_and2873_y0, h_u_cla24_and2872_y0, h_u_cla24_and2874_y0);
  and_gate and_gate_h_u_cla24_and2875_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and2875_y0);
  and_gate and_gate_h_u_cla24_and2876_y0(h_u_cla24_and2875_y0, h_u_cla24_and2874_y0, h_u_cla24_and2876_y0);
  and_gate and_gate_h_u_cla24_and2877_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and2877_y0);
  and_gate and_gate_h_u_cla24_and2878_y0(h_u_cla24_and2877_y0, h_u_cla24_and2876_y0, h_u_cla24_and2878_y0);
  and_gate and_gate_h_u_cla24_and2879_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and2879_y0);
  and_gate and_gate_h_u_cla24_and2880_y0(h_u_cla24_and2879_y0, h_u_cla24_and2878_y0, h_u_cla24_and2880_y0);
  and_gate and_gate_h_u_cla24_and2881_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and2881_y0);
  and_gate and_gate_h_u_cla24_and2882_y0(h_u_cla24_and2881_y0, h_u_cla24_and2880_y0, h_u_cla24_and2882_y0);
  and_gate and_gate_h_u_cla24_and2883_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and2883_y0);
  and_gate and_gate_h_u_cla24_and2884_y0(h_u_cla24_and2883_y0, h_u_cla24_and2882_y0, h_u_cla24_and2884_y0);
  and_gate and_gate_h_u_cla24_and2885_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and2885_y0);
  and_gate and_gate_h_u_cla24_and2886_y0(h_u_cla24_and2885_y0, h_u_cla24_and2884_y0, h_u_cla24_and2886_y0);
  and_gate and_gate_h_u_cla24_and2887_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and2887_y0);
  and_gate and_gate_h_u_cla24_and2888_y0(h_u_cla24_and2887_y0, h_u_cla24_and2886_y0, h_u_cla24_and2888_y0);
  and_gate and_gate_h_u_cla24_and2889_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and2889_y0);
  and_gate and_gate_h_u_cla24_and2890_y0(h_u_cla24_and2889_y0, h_u_cla24_and2888_y0, h_u_cla24_and2890_y0);
  and_gate and_gate_h_u_cla24_and2891_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and2891_y0);
  and_gate and_gate_h_u_cla24_and2892_y0(h_u_cla24_and2891_y0, h_u_cla24_and2890_y0, h_u_cla24_and2892_y0);
  and_gate and_gate_h_u_cla24_and2893_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and2893_y0);
  and_gate and_gate_h_u_cla24_and2894_y0(h_u_cla24_and2893_y0, h_u_cla24_and2892_y0, h_u_cla24_and2894_y0);
  and_gate and_gate_h_u_cla24_and2895_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and2895_y0);
  and_gate and_gate_h_u_cla24_and2896_y0(h_u_cla24_and2895_y0, h_u_cla24_and2894_y0, h_u_cla24_and2896_y0);
  and_gate and_gate_h_u_cla24_and2897_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and2897_y0);
  and_gate and_gate_h_u_cla24_and2898_y0(h_u_cla24_and2897_y0, h_u_cla24_and2896_y0, h_u_cla24_and2898_y0);
  and_gate and_gate_h_u_cla24_and2899_y0(h_u_cla24_pg_logic15_y0, constant_wire_0, h_u_cla24_and2899_y0);
  and_gate and_gate_h_u_cla24_and2900_y0(h_u_cla24_and2899_y0, h_u_cla24_and2898_y0, h_u_cla24_and2900_y0);
  and_gate and_gate_h_u_cla24_and2901_y0(h_u_cla24_pg_logic16_y0, constant_wire_0, h_u_cla24_and2901_y0);
  and_gate and_gate_h_u_cla24_and2902_y0(h_u_cla24_and2901_y0, h_u_cla24_and2900_y0, h_u_cla24_and2902_y0);
  and_gate and_gate_h_u_cla24_and2903_y0(h_u_cla24_pg_logic17_y0, constant_wire_0, h_u_cla24_and2903_y0);
  and_gate and_gate_h_u_cla24_and2904_y0(h_u_cla24_and2903_y0, h_u_cla24_and2902_y0, h_u_cla24_and2904_y0);
  and_gate and_gate_h_u_cla24_and2905_y0(h_u_cla24_pg_logic18_y0, constant_wire_0, h_u_cla24_and2905_y0);
  and_gate and_gate_h_u_cla24_and2906_y0(h_u_cla24_and2905_y0, h_u_cla24_and2904_y0, h_u_cla24_and2906_y0);
  and_gate and_gate_h_u_cla24_and2907_y0(h_u_cla24_pg_logic19_y0, constant_wire_0, h_u_cla24_and2907_y0);
  and_gate and_gate_h_u_cla24_and2908_y0(h_u_cla24_and2907_y0, h_u_cla24_and2906_y0, h_u_cla24_and2908_y0);
  and_gate and_gate_h_u_cla24_and2909_y0(h_u_cla24_pg_logic20_y0, constant_wire_0, h_u_cla24_and2909_y0);
  and_gate and_gate_h_u_cla24_and2910_y0(h_u_cla24_and2909_y0, h_u_cla24_and2908_y0, h_u_cla24_and2910_y0);
  and_gate and_gate_h_u_cla24_and2911_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2911_y0);
  and_gate and_gate_h_u_cla24_and2912_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2912_y0);
  and_gate and_gate_h_u_cla24_and2913_y0(h_u_cla24_and2912_y0, h_u_cla24_and2911_y0, h_u_cla24_and2913_y0);
  and_gate and_gate_h_u_cla24_and2914_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2914_y0);
  and_gate and_gate_h_u_cla24_and2915_y0(h_u_cla24_and2914_y0, h_u_cla24_and2913_y0, h_u_cla24_and2915_y0);
  and_gate and_gate_h_u_cla24_and2916_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2916_y0);
  and_gate and_gate_h_u_cla24_and2917_y0(h_u_cla24_and2916_y0, h_u_cla24_and2915_y0, h_u_cla24_and2917_y0);
  and_gate and_gate_h_u_cla24_and2918_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2918_y0);
  and_gate and_gate_h_u_cla24_and2919_y0(h_u_cla24_and2918_y0, h_u_cla24_and2917_y0, h_u_cla24_and2919_y0);
  and_gate and_gate_h_u_cla24_and2920_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2920_y0);
  and_gate and_gate_h_u_cla24_and2921_y0(h_u_cla24_and2920_y0, h_u_cla24_and2919_y0, h_u_cla24_and2921_y0);
  and_gate and_gate_h_u_cla24_and2922_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2922_y0);
  and_gate and_gate_h_u_cla24_and2923_y0(h_u_cla24_and2922_y0, h_u_cla24_and2921_y0, h_u_cla24_and2923_y0);
  and_gate and_gate_h_u_cla24_and2924_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2924_y0);
  and_gate and_gate_h_u_cla24_and2925_y0(h_u_cla24_and2924_y0, h_u_cla24_and2923_y0, h_u_cla24_and2925_y0);
  and_gate and_gate_h_u_cla24_and2926_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2926_y0);
  and_gate and_gate_h_u_cla24_and2927_y0(h_u_cla24_and2926_y0, h_u_cla24_and2925_y0, h_u_cla24_and2927_y0);
  and_gate and_gate_h_u_cla24_and2928_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2928_y0);
  and_gate and_gate_h_u_cla24_and2929_y0(h_u_cla24_and2928_y0, h_u_cla24_and2927_y0, h_u_cla24_and2929_y0);
  and_gate and_gate_h_u_cla24_and2930_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2930_y0);
  and_gate and_gate_h_u_cla24_and2931_y0(h_u_cla24_and2930_y0, h_u_cla24_and2929_y0, h_u_cla24_and2931_y0);
  and_gate and_gate_h_u_cla24_and2932_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2932_y0);
  and_gate and_gate_h_u_cla24_and2933_y0(h_u_cla24_and2932_y0, h_u_cla24_and2931_y0, h_u_cla24_and2933_y0);
  and_gate and_gate_h_u_cla24_and2934_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2934_y0);
  and_gate and_gate_h_u_cla24_and2935_y0(h_u_cla24_and2934_y0, h_u_cla24_and2933_y0, h_u_cla24_and2935_y0);
  and_gate and_gate_h_u_cla24_and2936_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2936_y0);
  and_gate and_gate_h_u_cla24_and2937_y0(h_u_cla24_and2936_y0, h_u_cla24_and2935_y0, h_u_cla24_and2937_y0);
  and_gate and_gate_h_u_cla24_and2938_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2938_y0);
  and_gate and_gate_h_u_cla24_and2939_y0(h_u_cla24_and2938_y0, h_u_cla24_and2937_y0, h_u_cla24_and2939_y0);
  and_gate and_gate_h_u_cla24_and2940_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2940_y0);
  and_gate and_gate_h_u_cla24_and2941_y0(h_u_cla24_and2940_y0, h_u_cla24_and2939_y0, h_u_cla24_and2941_y0);
  and_gate and_gate_h_u_cla24_and2942_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2942_y0);
  and_gate and_gate_h_u_cla24_and2943_y0(h_u_cla24_and2942_y0, h_u_cla24_and2941_y0, h_u_cla24_and2943_y0);
  and_gate and_gate_h_u_cla24_and2944_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2944_y0);
  and_gate and_gate_h_u_cla24_and2945_y0(h_u_cla24_and2944_y0, h_u_cla24_and2943_y0, h_u_cla24_and2945_y0);
  and_gate and_gate_h_u_cla24_and2946_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2946_y0);
  and_gate and_gate_h_u_cla24_and2947_y0(h_u_cla24_and2946_y0, h_u_cla24_and2945_y0, h_u_cla24_and2947_y0);
  and_gate and_gate_h_u_cla24_and2948_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and2948_y0);
  and_gate and_gate_h_u_cla24_and2949_y0(h_u_cla24_and2948_y0, h_u_cla24_and2947_y0, h_u_cla24_and2949_y0);
  and_gate and_gate_h_u_cla24_and2950_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2950_y0);
  and_gate and_gate_h_u_cla24_and2951_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2951_y0);
  and_gate and_gate_h_u_cla24_and2952_y0(h_u_cla24_and2951_y0, h_u_cla24_and2950_y0, h_u_cla24_and2952_y0);
  and_gate and_gate_h_u_cla24_and2953_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2953_y0);
  and_gate and_gate_h_u_cla24_and2954_y0(h_u_cla24_and2953_y0, h_u_cla24_and2952_y0, h_u_cla24_and2954_y0);
  and_gate and_gate_h_u_cla24_and2955_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2955_y0);
  and_gate and_gate_h_u_cla24_and2956_y0(h_u_cla24_and2955_y0, h_u_cla24_and2954_y0, h_u_cla24_and2956_y0);
  and_gate and_gate_h_u_cla24_and2957_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2957_y0);
  and_gate and_gate_h_u_cla24_and2958_y0(h_u_cla24_and2957_y0, h_u_cla24_and2956_y0, h_u_cla24_and2958_y0);
  and_gate and_gate_h_u_cla24_and2959_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2959_y0);
  and_gate and_gate_h_u_cla24_and2960_y0(h_u_cla24_and2959_y0, h_u_cla24_and2958_y0, h_u_cla24_and2960_y0);
  and_gate and_gate_h_u_cla24_and2961_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2961_y0);
  and_gate and_gate_h_u_cla24_and2962_y0(h_u_cla24_and2961_y0, h_u_cla24_and2960_y0, h_u_cla24_and2962_y0);
  and_gate and_gate_h_u_cla24_and2963_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2963_y0);
  and_gate and_gate_h_u_cla24_and2964_y0(h_u_cla24_and2963_y0, h_u_cla24_and2962_y0, h_u_cla24_and2964_y0);
  and_gate and_gate_h_u_cla24_and2965_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2965_y0);
  and_gate and_gate_h_u_cla24_and2966_y0(h_u_cla24_and2965_y0, h_u_cla24_and2964_y0, h_u_cla24_and2966_y0);
  and_gate and_gate_h_u_cla24_and2967_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2967_y0);
  and_gate and_gate_h_u_cla24_and2968_y0(h_u_cla24_and2967_y0, h_u_cla24_and2966_y0, h_u_cla24_and2968_y0);
  and_gate and_gate_h_u_cla24_and2969_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2969_y0);
  and_gate and_gate_h_u_cla24_and2970_y0(h_u_cla24_and2969_y0, h_u_cla24_and2968_y0, h_u_cla24_and2970_y0);
  and_gate and_gate_h_u_cla24_and2971_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2971_y0);
  and_gate and_gate_h_u_cla24_and2972_y0(h_u_cla24_and2971_y0, h_u_cla24_and2970_y0, h_u_cla24_and2972_y0);
  and_gate and_gate_h_u_cla24_and2973_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2973_y0);
  and_gate and_gate_h_u_cla24_and2974_y0(h_u_cla24_and2973_y0, h_u_cla24_and2972_y0, h_u_cla24_and2974_y0);
  and_gate and_gate_h_u_cla24_and2975_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2975_y0);
  and_gate and_gate_h_u_cla24_and2976_y0(h_u_cla24_and2975_y0, h_u_cla24_and2974_y0, h_u_cla24_and2976_y0);
  and_gate and_gate_h_u_cla24_and2977_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2977_y0);
  and_gate and_gate_h_u_cla24_and2978_y0(h_u_cla24_and2977_y0, h_u_cla24_and2976_y0, h_u_cla24_and2978_y0);
  and_gate and_gate_h_u_cla24_and2979_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2979_y0);
  and_gate and_gate_h_u_cla24_and2980_y0(h_u_cla24_and2979_y0, h_u_cla24_and2978_y0, h_u_cla24_and2980_y0);
  and_gate and_gate_h_u_cla24_and2981_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2981_y0);
  and_gate and_gate_h_u_cla24_and2982_y0(h_u_cla24_and2981_y0, h_u_cla24_and2980_y0, h_u_cla24_and2982_y0);
  and_gate and_gate_h_u_cla24_and2983_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2983_y0);
  and_gate and_gate_h_u_cla24_and2984_y0(h_u_cla24_and2983_y0, h_u_cla24_and2982_y0, h_u_cla24_and2984_y0);
  and_gate and_gate_h_u_cla24_and2985_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and2985_y0);
  and_gate and_gate_h_u_cla24_and2986_y0(h_u_cla24_and2985_y0, h_u_cla24_and2984_y0, h_u_cla24_and2986_y0);
  and_gate and_gate_h_u_cla24_and2987_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2987_y0);
  and_gate and_gate_h_u_cla24_and2988_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2988_y0);
  and_gate and_gate_h_u_cla24_and2989_y0(h_u_cla24_and2988_y0, h_u_cla24_and2987_y0, h_u_cla24_and2989_y0);
  and_gate and_gate_h_u_cla24_and2990_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2990_y0);
  and_gate and_gate_h_u_cla24_and2991_y0(h_u_cla24_and2990_y0, h_u_cla24_and2989_y0, h_u_cla24_and2991_y0);
  and_gate and_gate_h_u_cla24_and2992_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2992_y0);
  and_gate and_gate_h_u_cla24_and2993_y0(h_u_cla24_and2992_y0, h_u_cla24_and2991_y0, h_u_cla24_and2993_y0);
  and_gate and_gate_h_u_cla24_and2994_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2994_y0);
  and_gate and_gate_h_u_cla24_and2995_y0(h_u_cla24_and2994_y0, h_u_cla24_and2993_y0, h_u_cla24_and2995_y0);
  and_gate and_gate_h_u_cla24_and2996_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2996_y0);
  and_gate and_gate_h_u_cla24_and2997_y0(h_u_cla24_and2996_y0, h_u_cla24_and2995_y0, h_u_cla24_and2997_y0);
  and_gate and_gate_h_u_cla24_and2998_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and2998_y0);
  and_gate and_gate_h_u_cla24_and2999_y0(h_u_cla24_and2998_y0, h_u_cla24_and2997_y0, h_u_cla24_and2999_y0);
  and_gate and_gate_h_u_cla24_and3000_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3000_y0);
  and_gate and_gate_h_u_cla24_and3001_y0(h_u_cla24_and3000_y0, h_u_cla24_and2999_y0, h_u_cla24_and3001_y0);
  and_gate and_gate_h_u_cla24_and3002_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3002_y0);
  and_gate and_gate_h_u_cla24_and3003_y0(h_u_cla24_and3002_y0, h_u_cla24_and3001_y0, h_u_cla24_and3003_y0);
  and_gate and_gate_h_u_cla24_and3004_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3004_y0);
  and_gate and_gate_h_u_cla24_and3005_y0(h_u_cla24_and3004_y0, h_u_cla24_and3003_y0, h_u_cla24_and3005_y0);
  and_gate and_gate_h_u_cla24_and3006_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3006_y0);
  and_gate and_gate_h_u_cla24_and3007_y0(h_u_cla24_and3006_y0, h_u_cla24_and3005_y0, h_u_cla24_and3007_y0);
  and_gate and_gate_h_u_cla24_and3008_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3008_y0);
  and_gate and_gate_h_u_cla24_and3009_y0(h_u_cla24_and3008_y0, h_u_cla24_and3007_y0, h_u_cla24_and3009_y0);
  and_gate and_gate_h_u_cla24_and3010_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3010_y0);
  and_gate and_gate_h_u_cla24_and3011_y0(h_u_cla24_and3010_y0, h_u_cla24_and3009_y0, h_u_cla24_and3011_y0);
  and_gate and_gate_h_u_cla24_and3012_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3012_y0);
  and_gate and_gate_h_u_cla24_and3013_y0(h_u_cla24_and3012_y0, h_u_cla24_and3011_y0, h_u_cla24_and3013_y0);
  and_gate and_gate_h_u_cla24_and3014_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3014_y0);
  and_gate and_gate_h_u_cla24_and3015_y0(h_u_cla24_and3014_y0, h_u_cla24_and3013_y0, h_u_cla24_and3015_y0);
  and_gate and_gate_h_u_cla24_and3016_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3016_y0);
  and_gate and_gate_h_u_cla24_and3017_y0(h_u_cla24_and3016_y0, h_u_cla24_and3015_y0, h_u_cla24_and3017_y0);
  and_gate and_gate_h_u_cla24_and3018_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3018_y0);
  and_gate and_gate_h_u_cla24_and3019_y0(h_u_cla24_and3018_y0, h_u_cla24_and3017_y0, h_u_cla24_and3019_y0);
  and_gate and_gate_h_u_cla24_and3020_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3020_y0);
  and_gate and_gate_h_u_cla24_and3021_y0(h_u_cla24_and3020_y0, h_u_cla24_and3019_y0, h_u_cla24_and3021_y0);
  and_gate and_gate_h_u_cla24_and3022_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3022_y0);
  and_gate and_gate_h_u_cla24_and3023_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3023_y0);
  and_gate and_gate_h_u_cla24_and3024_y0(h_u_cla24_and3023_y0, h_u_cla24_and3022_y0, h_u_cla24_and3024_y0);
  and_gate and_gate_h_u_cla24_and3025_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3025_y0);
  and_gate and_gate_h_u_cla24_and3026_y0(h_u_cla24_and3025_y0, h_u_cla24_and3024_y0, h_u_cla24_and3026_y0);
  and_gate and_gate_h_u_cla24_and3027_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3027_y0);
  and_gate and_gate_h_u_cla24_and3028_y0(h_u_cla24_and3027_y0, h_u_cla24_and3026_y0, h_u_cla24_and3028_y0);
  and_gate and_gate_h_u_cla24_and3029_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3029_y0);
  and_gate and_gate_h_u_cla24_and3030_y0(h_u_cla24_and3029_y0, h_u_cla24_and3028_y0, h_u_cla24_and3030_y0);
  and_gate and_gate_h_u_cla24_and3031_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3031_y0);
  and_gate and_gate_h_u_cla24_and3032_y0(h_u_cla24_and3031_y0, h_u_cla24_and3030_y0, h_u_cla24_and3032_y0);
  and_gate and_gate_h_u_cla24_and3033_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3033_y0);
  and_gate and_gate_h_u_cla24_and3034_y0(h_u_cla24_and3033_y0, h_u_cla24_and3032_y0, h_u_cla24_and3034_y0);
  and_gate and_gate_h_u_cla24_and3035_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3035_y0);
  and_gate and_gate_h_u_cla24_and3036_y0(h_u_cla24_and3035_y0, h_u_cla24_and3034_y0, h_u_cla24_and3036_y0);
  and_gate and_gate_h_u_cla24_and3037_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3037_y0);
  and_gate and_gate_h_u_cla24_and3038_y0(h_u_cla24_and3037_y0, h_u_cla24_and3036_y0, h_u_cla24_and3038_y0);
  and_gate and_gate_h_u_cla24_and3039_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3039_y0);
  and_gate and_gate_h_u_cla24_and3040_y0(h_u_cla24_and3039_y0, h_u_cla24_and3038_y0, h_u_cla24_and3040_y0);
  and_gate and_gate_h_u_cla24_and3041_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3041_y0);
  and_gate and_gate_h_u_cla24_and3042_y0(h_u_cla24_and3041_y0, h_u_cla24_and3040_y0, h_u_cla24_and3042_y0);
  and_gate and_gate_h_u_cla24_and3043_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3043_y0);
  and_gate and_gate_h_u_cla24_and3044_y0(h_u_cla24_and3043_y0, h_u_cla24_and3042_y0, h_u_cla24_and3044_y0);
  and_gate and_gate_h_u_cla24_and3045_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3045_y0);
  and_gate and_gate_h_u_cla24_and3046_y0(h_u_cla24_and3045_y0, h_u_cla24_and3044_y0, h_u_cla24_and3046_y0);
  and_gate and_gate_h_u_cla24_and3047_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3047_y0);
  and_gate and_gate_h_u_cla24_and3048_y0(h_u_cla24_and3047_y0, h_u_cla24_and3046_y0, h_u_cla24_and3048_y0);
  and_gate and_gate_h_u_cla24_and3049_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3049_y0);
  and_gate and_gate_h_u_cla24_and3050_y0(h_u_cla24_and3049_y0, h_u_cla24_and3048_y0, h_u_cla24_and3050_y0);
  and_gate and_gate_h_u_cla24_and3051_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3051_y0);
  and_gate and_gate_h_u_cla24_and3052_y0(h_u_cla24_and3051_y0, h_u_cla24_and3050_y0, h_u_cla24_and3052_y0);
  and_gate and_gate_h_u_cla24_and3053_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3053_y0);
  and_gate and_gate_h_u_cla24_and3054_y0(h_u_cla24_and3053_y0, h_u_cla24_and3052_y0, h_u_cla24_and3054_y0);
  and_gate and_gate_h_u_cla24_and3055_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3055_y0);
  and_gate and_gate_h_u_cla24_and3056_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3056_y0);
  and_gate and_gate_h_u_cla24_and3057_y0(h_u_cla24_and3056_y0, h_u_cla24_and3055_y0, h_u_cla24_and3057_y0);
  and_gate and_gate_h_u_cla24_and3058_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3058_y0);
  and_gate and_gate_h_u_cla24_and3059_y0(h_u_cla24_and3058_y0, h_u_cla24_and3057_y0, h_u_cla24_and3059_y0);
  and_gate and_gate_h_u_cla24_and3060_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3060_y0);
  and_gate and_gate_h_u_cla24_and3061_y0(h_u_cla24_and3060_y0, h_u_cla24_and3059_y0, h_u_cla24_and3061_y0);
  and_gate and_gate_h_u_cla24_and3062_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3062_y0);
  and_gate and_gate_h_u_cla24_and3063_y0(h_u_cla24_and3062_y0, h_u_cla24_and3061_y0, h_u_cla24_and3063_y0);
  and_gate and_gate_h_u_cla24_and3064_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3064_y0);
  and_gate and_gate_h_u_cla24_and3065_y0(h_u_cla24_and3064_y0, h_u_cla24_and3063_y0, h_u_cla24_and3065_y0);
  and_gate and_gate_h_u_cla24_and3066_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3066_y0);
  and_gate and_gate_h_u_cla24_and3067_y0(h_u_cla24_and3066_y0, h_u_cla24_and3065_y0, h_u_cla24_and3067_y0);
  and_gate and_gate_h_u_cla24_and3068_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3068_y0);
  and_gate and_gate_h_u_cla24_and3069_y0(h_u_cla24_and3068_y0, h_u_cla24_and3067_y0, h_u_cla24_and3069_y0);
  and_gate and_gate_h_u_cla24_and3070_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3070_y0);
  and_gate and_gate_h_u_cla24_and3071_y0(h_u_cla24_and3070_y0, h_u_cla24_and3069_y0, h_u_cla24_and3071_y0);
  and_gate and_gate_h_u_cla24_and3072_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3072_y0);
  and_gate and_gate_h_u_cla24_and3073_y0(h_u_cla24_and3072_y0, h_u_cla24_and3071_y0, h_u_cla24_and3073_y0);
  and_gate and_gate_h_u_cla24_and3074_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3074_y0);
  and_gate and_gate_h_u_cla24_and3075_y0(h_u_cla24_and3074_y0, h_u_cla24_and3073_y0, h_u_cla24_and3075_y0);
  and_gate and_gate_h_u_cla24_and3076_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3076_y0);
  and_gate and_gate_h_u_cla24_and3077_y0(h_u_cla24_and3076_y0, h_u_cla24_and3075_y0, h_u_cla24_and3077_y0);
  and_gate and_gate_h_u_cla24_and3078_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3078_y0);
  and_gate and_gate_h_u_cla24_and3079_y0(h_u_cla24_and3078_y0, h_u_cla24_and3077_y0, h_u_cla24_and3079_y0);
  and_gate and_gate_h_u_cla24_and3080_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3080_y0);
  and_gate and_gate_h_u_cla24_and3081_y0(h_u_cla24_and3080_y0, h_u_cla24_and3079_y0, h_u_cla24_and3081_y0);
  and_gate and_gate_h_u_cla24_and3082_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3082_y0);
  and_gate and_gate_h_u_cla24_and3083_y0(h_u_cla24_and3082_y0, h_u_cla24_and3081_y0, h_u_cla24_and3083_y0);
  and_gate and_gate_h_u_cla24_and3084_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3084_y0);
  and_gate and_gate_h_u_cla24_and3085_y0(h_u_cla24_and3084_y0, h_u_cla24_and3083_y0, h_u_cla24_and3085_y0);
  and_gate and_gate_h_u_cla24_and3086_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3086_y0);
  and_gate and_gate_h_u_cla24_and3087_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3087_y0);
  and_gate and_gate_h_u_cla24_and3088_y0(h_u_cla24_and3087_y0, h_u_cla24_and3086_y0, h_u_cla24_and3088_y0);
  and_gate and_gate_h_u_cla24_and3089_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3089_y0);
  and_gate and_gate_h_u_cla24_and3090_y0(h_u_cla24_and3089_y0, h_u_cla24_and3088_y0, h_u_cla24_and3090_y0);
  and_gate and_gate_h_u_cla24_and3091_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3091_y0);
  and_gate and_gate_h_u_cla24_and3092_y0(h_u_cla24_and3091_y0, h_u_cla24_and3090_y0, h_u_cla24_and3092_y0);
  and_gate and_gate_h_u_cla24_and3093_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3093_y0);
  and_gate and_gate_h_u_cla24_and3094_y0(h_u_cla24_and3093_y0, h_u_cla24_and3092_y0, h_u_cla24_and3094_y0);
  and_gate and_gate_h_u_cla24_and3095_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3095_y0);
  and_gate and_gate_h_u_cla24_and3096_y0(h_u_cla24_and3095_y0, h_u_cla24_and3094_y0, h_u_cla24_and3096_y0);
  and_gate and_gate_h_u_cla24_and3097_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3097_y0);
  and_gate and_gate_h_u_cla24_and3098_y0(h_u_cla24_and3097_y0, h_u_cla24_and3096_y0, h_u_cla24_and3098_y0);
  and_gate and_gate_h_u_cla24_and3099_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3099_y0);
  and_gate and_gate_h_u_cla24_and3100_y0(h_u_cla24_and3099_y0, h_u_cla24_and3098_y0, h_u_cla24_and3100_y0);
  and_gate and_gate_h_u_cla24_and3101_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3101_y0);
  and_gate and_gate_h_u_cla24_and3102_y0(h_u_cla24_and3101_y0, h_u_cla24_and3100_y0, h_u_cla24_and3102_y0);
  and_gate and_gate_h_u_cla24_and3103_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3103_y0);
  and_gate and_gate_h_u_cla24_and3104_y0(h_u_cla24_and3103_y0, h_u_cla24_and3102_y0, h_u_cla24_and3104_y0);
  and_gate and_gate_h_u_cla24_and3105_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3105_y0);
  and_gate and_gate_h_u_cla24_and3106_y0(h_u_cla24_and3105_y0, h_u_cla24_and3104_y0, h_u_cla24_and3106_y0);
  and_gate and_gate_h_u_cla24_and3107_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3107_y0);
  and_gate and_gate_h_u_cla24_and3108_y0(h_u_cla24_and3107_y0, h_u_cla24_and3106_y0, h_u_cla24_and3108_y0);
  and_gate and_gate_h_u_cla24_and3109_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3109_y0);
  and_gate and_gate_h_u_cla24_and3110_y0(h_u_cla24_and3109_y0, h_u_cla24_and3108_y0, h_u_cla24_and3110_y0);
  and_gate and_gate_h_u_cla24_and3111_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3111_y0);
  and_gate and_gate_h_u_cla24_and3112_y0(h_u_cla24_and3111_y0, h_u_cla24_and3110_y0, h_u_cla24_and3112_y0);
  and_gate and_gate_h_u_cla24_and3113_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3113_y0);
  and_gate and_gate_h_u_cla24_and3114_y0(h_u_cla24_and3113_y0, h_u_cla24_and3112_y0, h_u_cla24_and3114_y0);
  and_gate and_gate_h_u_cla24_and3115_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3115_y0);
  and_gate and_gate_h_u_cla24_and3116_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3116_y0);
  and_gate and_gate_h_u_cla24_and3117_y0(h_u_cla24_and3116_y0, h_u_cla24_and3115_y0, h_u_cla24_and3117_y0);
  and_gate and_gate_h_u_cla24_and3118_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3118_y0);
  and_gate and_gate_h_u_cla24_and3119_y0(h_u_cla24_and3118_y0, h_u_cla24_and3117_y0, h_u_cla24_and3119_y0);
  and_gate and_gate_h_u_cla24_and3120_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3120_y0);
  and_gate and_gate_h_u_cla24_and3121_y0(h_u_cla24_and3120_y0, h_u_cla24_and3119_y0, h_u_cla24_and3121_y0);
  and_gate and_gate_h_u_cla24_and3122_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3122_y0);
  and_gate and_gate_h_u_cla24_and3123_y0(h_u_cla24_and3122_y0, h_u_cla24_and3121_y0, h_u_cla24_and3123_y0);
  and_gate and_gate_h_u_cla24_and3124_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3124_y0);
  and_gate and_gate_h_u_cla24_and3125_y0(h_u_cla24_and3124_y0, h_u_cla24_and3123_y0, h_u_cla24_and3125_y0);
  and_gate and_gate_h_u_cla24_and3126_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3126_y0);
  and_gate and_gate_h_u_cla24_and3127_y0(h_u_cla24_and3126_y0, h_u_cla24_and3125_y0, h_u_cla24_and3127_y0);
  and_gate and_gate_h_u_cla24_and3128_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3128_y0);
  and_gate and_gate_h_u_cla24_and3129_y0(h_u_cla24_and3128_y0, h_u_cla24_and3127_y0, h_u_cla24_and3129_y0);
  and_gate and_gate_h_u_cla24_and3130_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3130_y0);
  and_gate and_gate_h_u_cla24_and3131_y0(h_u_cla24_and3130_y0, h_u_cla24_and3129_y0, h_u_cla24_and3131_y0);
  and_gate and_gate_h_u_cla24_and3132_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3132_y0);
  and_gate and_gate_h_u_cla24_and3133_y0(h_u_cla24_and3132_y0, h_u_cla24_and3131_y0, h_u_cla24_and3133_y0);
  and_gate and_gate_h_u_cla24_and3134_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3134_y0);
  and_gate and_gate_h_u_cla24_and3135_y0(h_u_cla24_and3134_y0, h_u_cla24_and3133_y0, h_u_cla24_and3135_y0);
  and_gate and_gate_h_u_cla24_and3136_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3136_y0);
  and_gate and_gate_h_u_cla24_and3137_y0(h_u_cla24_and3136_y0, h_u_cla24_and3135_y0, h_u_cla24_and3137_y0);
  and_gate and_gate_h_u_cla24_and3138_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3138_y0);
  and_gate and_gate_h_u_cla24_and3139_y0(h_u_cla24_and3138_y0, h_u_cla24_and3137_y0, h_u_cla24_and3139_y0);
  and_gate and_gate_h_u_cla24_and3140_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3140_y0);
  and_gate and_gate_h_u_cla24_and3141_y0(h_u_cla24_and3140_y0, h_u_cla24_and3139_y0, h_u_cla24_and3141_y0);
  and_gate and_gate_h_u_cla24_and3142_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3142_y0);
  and_gate and_gate_h_u_cla24_and3143_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3143_y0);
  and_gate and_gate_h_u_cla24_and3144_y0(h_u_cla24_and3143_y0, h_u_cla24_and3142_y0, h_u_cla24_and3144_y0);
  and_gate and_gate_h_u_cla24_and3145_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3145_y0);
  and_gate and_gate_h_u_cla24_and3146_y0(h_u_cla24_and3145_y0, h_u_cla24_and3144_y0, h_u_cla24_and3146_y0);
  and_gate and_gate_h_u_cla24_and3147_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3147_y0);
  and_gate and_gate_h_u_cla24_and3148_y0(h_u_cla24_and3147_y0, h_u_cla24_and3146_y0, h_u_cla24_and3148_y0);
  and_gate and_gate_h_u_cla24_and3149_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3149_y0);
  and_gate and_gate_h_u_cla24_and3150_y0(h_u_cla24_and3149_y0, h_u_cla24_and3148_y0, h_u_cla24_and3150_y0);
  and_gate and_gate_h_u_cla24_and3151_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3151_y0);
  and_gate and_gate_h_u_cla24_and3152_y0(h_u_cla24_and3151_y0, h_u_cla24_and3150_y0, h_u_cla24_and3152_y0);
  and_gate and_gate_h_u_cla24_and3153_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3153_y0);
  and_gate and_gate_h_u_cla24_and3154_y0(h_u_cla24_and3153_y0, h_u_cla24_and3152_y0, h_u_cla24_and3154_y0);
  and_gate and_gate_h_u_cla24_and3155_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3155_y0);
  and_gate and_gate_h_u_cla24_and3156_y0(h_u_cla24_and3155_y0, h_u_cla24_and3154_y0, h_u_cla24_and3156_y0);
  and_gate and_gate_h_u_cla24_and3157_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3157_y0);
  and_gate and_gate_h_u_cla24_and3158_y0(h_u_cla24_and3157_y0, h_u_cla24_and3156_y0, h_u_cla24_and3158_y0);
  and_gate and_gate_h_u_cla24_and3159_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3159_y0);
  and_gate and_gate_h_u_cla24_and3160_y0(h_u_cla24_and3159_y0, h_u_cla24_and3158_y0, h_u_cla24_and3160_y0);
  and_gate and_gate_h_u_cla24_and3161_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3161_y0);
  and_gate and_gate_h_u_cla24_and3162_y0(h_u_cla24_and3161_y0, h_u_cla24_and3160_y0, h_u_cla24_and3162_y0);
  and_gate and_gate_h_u_cla24_and3163_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3163_y0);
  and_gate and_gate_h_u_cla24_and3164_y0(h_u_cla24_and3163_y0, h_u_cla24_and3162_y0, h_u_cla24_and3164_y0);
  and_gate and_gate_h_u_cla24_and3165_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3165_y0);
  and_gate and_gate_h_u_cla24_and3166_y0(h_u_cla24_and3165_y0, h_u_cla24_and3164_y0, h_u_cla24_and3166_y0);
  and_gate and_gate_h_u_cla24_and3167_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3167_y0);
  and_gate and_gate_h_u_cla24_and3168_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3168_y0);
  and_gate and_gate_h_u_cla24_and3169_y0(h_u_cla24_and3168_y0, h_u_cla24_and3167_y0, h_u_cla24_and3169_y0);
  and_gate and_gate_h_u_cla24_and3170_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3170_y0);
  and_gate and_gate_h_u_cla24_and3171_y0(h_u_cla24_and3170_y0, h_u_cla24_and3169_y0, h_u_cla24_and3171_y0);
  and_gate and_gate_h_u_cla24_and3172_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3172_y0);
  and_gate and_gate_h_u_cla24_and3173_y0(h_u_cla24_and3172_y0, h_u_cla24_and3171_y0, h_u_cla24_and3173_y0);
  and_gate and_gate_h_u_cla24_and3174_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3174_y0);
  and_gate and_gate_h_u_cla24_and3175_y0(h_u_cla24_and3174_y0, h_u_cla24_and3173_y0, h_u_cla24_and3175_y0);
  and_gate and_gate_h_u_cla24_and3176_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3176_y0);
  and_gate and_gate_h_u_cla24_and3177_y0(h_u_cla24_and3176_y0, h_u_cla24_and3175_y0, h_u_cla24_and3177_y0);
  and_gate and_gate_h_u_cla24_and3178_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3178_y0);
  and_gate and_gate_h_u_cla24_and3179_y0(h_u_cla24_and3178_y0, h_u_cla24_and3177_y0, h_u_cla24_and3179_y0);
  and_gate and_gate_h_u_cla24_and3180_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3180_y0);
  and_gate and_gate_h_u_cla24_and3181_y0(h_u_cla24_and3180_y0, h_u_cla24_and3179_y0, h_u_cla24_and3181_y0);
  and_gate and_gate_h_u_cla24_and3182_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3182_y0);
  and_gate and_gate_h_u_cla24_and3183_y0(h_u_cla24_and3182_y0, h_u_cla24_and3181_y0, h_u_cla24_and3183_y0);
  and_gate and_gate_h_u_cla24_and3184_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3184_y0);
  and_gate and_gate_h_u_cla24_and3185_y0(h_u_cla24_and3184_y0, h_u_cla24_and3183_y0, h_u_cla24_and3185_y0);
  and_gate and_gate_h_u_cla24_and3186_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3186_y0);
  and_gate and_gate_h_u_cla24_and3187_y0(h_u_cla24_and3186_y0, h_u_cla24_and3185_y0, h_u_cla24_and3187_y0);
  and_gate and_gate_h_u_cla24_and3188_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3188_y0);
  and_gate and_gate_h_u_cla24_and3189_y0(h_u_cla24_and3188_y0, h_u_cla24_and3187_y0, h_u_cla24_and3189_y0);
  and_gate and_gate_h_u_cla24_and3190_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3190_y0);
  and_gate and_gate_h_u_cla24_and3191_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3191_y0);
  and_gate and_gate_h_u_cla24_and3192_y0(h_u_cla24_and3191_y0, h_u_cla24_and3190_y0, h_u_cla24_and3192_y0);
  and_gate and_gate_h_u_cla24_and3193_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3193_y0);
  and_gate and_gate_h_u_cla24_and3194_y0(h_u_cla24_and3193_y0, h_u_cla24_and3192_y0, h_u_cla24_and3194_y0);
  and_gate and_gate_h_u_cla24_and3195_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3195_y0);
  and_gate and_gate_h_u_cla24_and3196_y0(h_u_cla24_and3195_y0, h_u_cla24_and3194_y0, h_u_cla24_and3196_y0);
  and_gate and_gate_h_u_cla24_and3197_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3197_y0);
  and_gate and_gate_h_u_cla24_and3198_y0(h_u_cla24_and3197_y0, h_u_cla24_and3196_y0, h_u_cla24_and3198_y0);
  and_gate and_gate_h_u_cla24_and3199_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3199_y0);
  and_gate and_gate_h_u_cla24_and3200_y0(h_u_cla24_and3199_y0, h_u_cla24_and3198_y0, h_u_cla24_and3200_y0);
  and_gate and_gate_h_u_cla24_and3201_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3201_y0);
  and_gate and_gate_h_u_cla24_and3202_y0(h_u_cla24_and3201_y0, h_u_cla24_and3200_y0, h_u_cla24_and3202_y0);
  and_gate and_gate_h_u_cla24_and3203_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3203_y0);
  and_gate and_gate_h_u_cla24_and3204_y0(h_u_cla24_and3203_y0, h_u_cla24_and3202_y0, h_u_cla24_and3204_y0);
  and_gate and_gate_h_u_cla24_and3205_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3205_y0);
  and_gate and_gate_h_u_cla24_and3206_y0(h_u_cla24_and3205_y0, h_u_cla24_and3204_y0, h_u_cla24_and3206_y0);
  and_gate and_gate_h_u_cla24_and3207_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3207_y0);
  and_gate and_gate_h_u_cla24_and3208_y0(h_u_cla24_and3207_y0, h_u_cla24_and3206_y0, h_u_cla24_and3208_y0);
  and_gate and_gate_h_u_cla24_and3209_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3209_y0);
  and_gate and_gate_h_u_cla24_and3210_y0(h_u_cla24_and3209_y0, h_u_cla24_and3208_y0, h_u_cla24_and3210_y0);
  and_gate and_gate_h_u_cla24_and3211_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3211_y0);
  and_gate and_gate_h_u_cla24_and3212_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3212_y0);
  and_gate and_gate_h_u_cla24_and3213_y0(h_u_cla24_and3212_y0, h_u_cla24_and3211_y0, h_u_cla24_and3213_y0);
  and_gate and_gate_h_u_cla24_and3214_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3214_y0);
  and_gate and_gate_h_u_cla24_and3215_y0(h_u_cla24_and3214_y0, h_u_cla24_and3213_y0, h_u_cla24_and3215_y0);
  and_gate and_gate_h_u_cla24_and3216_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3216_y0);
  and_gate and_gate_h_u_cla24_and3217_y0(h_u_cla24_and3216_y0, h_u_cla24_and3215_y0, h_u_cla24_and3217_y0);
  and_gate and_gate_h_u_cla24_and3218_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3218_y0);
  and_gate and_gate_h_u_cla24_and3219_y0(h_u_cla24_and3218_y0, h_u_cla24_and3217_y0, h_u_cla24_and3219_y0);
  and_gate and_gate_h_u_cla24_and3220_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3220_y0);
  and_gate and_gate_h_u_cla24_and3221_y0(h_u_cla24_and3220_y0, h_u_cla24_and3219_y0, h_u_cla24_and3221_y0);
  and_gate and_gate_h_u_cla24_and3222_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3222_y0);
  and_gate and_gate_h_u_cla24_and3223_y0(h_u_cla24_and3222_y0, h_u_cla24_and3221_y0, h_u_cla24_and3223_y0);
  and_gate and_gate_h_u_cla24_and3224_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3224_y0);
  and_gate and_gate_h_u_cla24_and3225_y0(h_u_cla24_and3224_y0, h_u_cla24_and3223_y0, h_u_cla24_and3225_y0);
  and_gate and_gate_h_u_cla24_and3226_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3226_y0);
  and_gate and_gate_h_u_cla24_and3227_y0(h_u_cla24_and3226_y0, h_u_cla24_and3225_y0, h_u_cla24_and3227_y0);
  and_gate and_gate_h_u_cla24_and3228_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3228_y0);
  and_gate and_gate_h_u_cla24_and3229_y0(h_u_cla24_and3228_y0, h_u_cla24_and3227_y0, h_u_cla24_and3229_y0);
  and_gate and_gate_h_u_cla24_and3230_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3230_y0);
  and_gate and_gate_h_u_cla24_and3231_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3231_y0);
  and_gate and_gate_h_u_cla24_and3232_y0(h_u_cla24_and3231_y0, h_u_cla24_and3230_y0, h_u_cla24_and3232_y0);
  and_gate and_gate_h_u_cla24_and3233_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3233_y0);
  and_gate and_gate_h_u_cla24_and3234_y0(h_u_cla24_and3233_y0, h_u_cla24_and3232_y0, h_u_cla24_and3234_y0);
  and_gate and_gate_h_u_cla24_and3235_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3235_y0);
  and_gate and_gate_h_u_cla24_and3236_y0(h_u_cla24_and3235_y0, h_u_cla24_and3234_y0, h_u_cla24_and3236_y0);
  and_gate and_gate_h_u_cla24_and3237_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3237_y0);
  and_gate and_gate_h_u_cla24_and3238_y0(h_u_cla24_and3237_y0, h_u_cla24_and3236_y0, h_u_cla24_and3238_y0);
  and_gate and_gate_h_u_cla24_and3239_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3239_y0);
  and_gate and_gate_h_u_cla24_and3240_y0(h_u_cla24_and3239_y0, h_u_cla24_and3238_y0, h_u_cla24_and3240_y0);
  and_gate and_gate_h_u_cla24_and3241_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3241_y0);
  and_gate and_gate_h_u_cla24_and3242_y0(h_u_cla24_and3241_y0, h_u_cla24_and3240_y0, h_u_cla24_and3242_y0);
  and_gate and_gate_h_u_cla24_and3243_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3243_y0);
  and_gate and_gate_h_u_cla24_and3244_y0(h_u_cla24_and3243_y0, h_u_cla24_and3242_y0, h_u_cla24_and3244_y0);
  and_gate and_gate_h_u_cla24_and3245_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3245_y0);
  and_gate and_gate_h_u_cla24_and3246_y0(h_u_cla24_and3245_y0, h_u_cla24_and3244_y0, h_u_cla24_and3246_y0);
  and_gate and_gate_h_u_cla24_and3247_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3247_y0);
  and_gate and_gate_h_u_cla24_and3248_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3248_y0);
  and_gate and_gate_h_u_cla24_and3249_y0(h_u_cla24_and3248_y0, h_u_cla24_and3247_y0, h_u_cla24_and3249_y0);
  and_gate and_gate_h_u_cla24_and3250_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3250_y0);
  and_gate and_gate_h_u_cla24_and3251_y0(h_u_cla24_and3250_y0, h_u_cla24_and3249_y0, h_u_cla24_and3251_y0);
  and_gate and_gate_h_u_cla24_and3252_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3252_y0);
  and_gate and_gate_h_u_cla24_and3253_y0(h_u_cla24_and3252_y0, h_u_cla24_and3251_y0, h_u_cla24_and3253_y0);
  and_gate and_gate_h_u_cla24_and3254_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3254_y0);
  and_gate and_gate_h_u_cla24_and3255_y0(h_u_cla24_and3254_y0, h_u_cla24_and3253_y0, h_u_cla24_and3255_y0);
  and_gate and_gate_h_u_cla24_and3256_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3256_y0);
  and_gate and_gate_h_u_cla24_and3257_y0(h_u_cla24_and3256_y0, h_u_cla24_and3255_y0, h_u_cla24_and3257_y0);
  and_gate and_gate_h_u_cla24_and3258_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3258_y0);
  and_gate and_gate_h_u_cla24_and3259_y0(h_u_cla24_and3258_y0, h_u_cla24_and3257_y0, h_u_cla24_and3259_y0);
  and_gate and_gate_h_u_cla24_and3260_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3260_y0);
  and_gate and_gate_h_u_cla24_and3261_y0(h_u_cla24_and3260_y0, h_u_cla24_and3259_y0, h_u_cla24_and3261_y0);
  and_gate and_gate_h_u_cla24_and3262_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3262_y0);
  and_gate and_gate_h_u_cla24_and3263_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3263_y0);
  and_gate and_gate_h_u_cla24_and3264_y0(h_u_cla24_and3263_y0, h_u_cla24_and3262_y0, h_u_cla24_and3264_y0);
  and_gate and_gate_h_u_cla24_and3265_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3265_y0);
  and_gate and_gate_h_u_cla24_and3266_y0(h_u_cla24_and3265_y0, h_u_cla24_and3264_y0, h_u_cla24_and3266_y0);
  and_gate and_gate_h_u_cla24_and3267_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3267_y0);
  and_gate and_gate_h_u_cla24_and3268_y0(h_u_cla24_and3267_y0, h_u_cla24_and3266_y0, h_u_cla24_and3268_y0);
  and_gate and_gate_h_u_cla24_and3269_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3269_y0);
  and_gate and_gate_h_u_cla24_and3270_y0(h_u_cla24_and3269_y0, h_u_cla24_and3268_y0, h_u_cla24_and3270_y0);
  and_gate and_gate_h_u_cla24_and3271_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3271_y0);
  and_gate and_gate_h_u_cla24_and3272_y0(h_u_cla24_and3271_y0, h_u_cla24_and3270_y0, h_u_cla24_and3272_y0);
  and_gate and_gate_h_u_cla24_and3273_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3273_y0);
  and_gate and_gate_h_u_cla24_and3274_y0(h_u_cla24_and3273_y0, h_u_cla24_and3272_y0, h_u_cla24_and3274_y0);
  and_gate and_gate_h_u_cla24_and3275_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3275_y0);
  and_gate and_gate_h_u_cla24_and3276_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3276_y0);
  and_gate and_gate_h_u_cla24_and3277_y0(h_u_cla24_and3276_y0, h_u_cla24_and3275_y0, h_u_cla24_and3277_y0);
  and_gate and_gate_h_u_cla24_and3278_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3278_y0);
  and_gate and_gate_h_u_cla24_and3279_y0(h_u_cla24_and3278_y0, h_u_cla24_and3277_y0, h_u_cla24_and3279_y0);
  and_gate and_gate_h_u_cla24_and3280_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3280_y0);
  and_gate and_gate_h_u_cla24_and3281_y0(h_u_cla24_and3280_y0, h_u_cla24_and3279_y0, h_u_cla24_and3281_y0);
  and_gate and_gate_h_u_cla24_and3282_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3282_y0);
  and_gate and_gate_h_u_cla24_and3283_y0(h_u_cla24_and3282_y0, h_u_cla24_and3281_y0, h_u_cla24_and3283_y0);
  and_gate and_gate_h_u_cla24_and3284_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3284_y0);
  and_gate and_gate_h_u_cla24_and3285_y0(h_u_cla24_and3284_y0, h_u_cla24_and3283_y0, h_u_cla24_and3285_y0);
  and_gate and_gate_h_u_cla24_and3286_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3286_y0);
  and_gate and_gate_h_u_cla24_and3287_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3287_y0);
  and_gate and_gate_h_u_cla24_and3288_y0(h_u_cla24_and3287_y0, h_u_cla24_and3286_y0, h_u_cla24_and3288_y0);
  and_gate and_gate_h_u_cla24_and3289_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3289_y0);
  and_gate and_gate_h_u_cla24_and3290_y0(h_u_cla24_and3289_y0, h_u_cla24_and3288_y0, h_u_cla24_and3290_y0);
  and_gate and_gate_h_u_cla24_and3291_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3291_y0);
  and_gate and_gate_h_u_cla24_and3292_y0(h_u_cla24_and3291_y0, h_u_cla24_and3290_y0, h_u_cla24_and3292_y0);
  and_gate and_gate_h_u_cla24_and3293_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3293_y0);
  and_gate and_gate_h_u_cla24_and3294_y0(h_u_cla24_and3293_y0, h_u_cla24_and3292_y0, h_u_cla24_and3294_y0);
  and_gate and_gate_h_u_cla24_and3295_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and3295_y0);
  and_gate and_gate_h_u_cla24_and3296_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and3296_y0);
  and_gate and_gate_h_u_cla24_and3297_y0(h_u_cla24_and3296_y0, h_u_cla24_and3295_y0, h_u_cla24_and3297_y0);
  and_gate and_gate_h_u_cla24_and3298_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and3298_y0);
  and_gate and_gate_h_u_cla24_and3299_y0(h_u_cla24_and3298_y0, h_u_cla24_and3297_y0, h_u_cla24_and3299_y0);
  and_gate and_gate_h_u_cla24_and3300_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and3300_y0);
  and_gate and_gate_h_u_cla24_and3301_y0(h_u_cla24_and3300_y0, h_u_cla24_and3299_y0, h_u_cla24_and3301_y0);
  and_gate and_gate_h_u_cla24_and3302_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and3302_y0);
  and_gate and_gate_h_u_cla24_and3303_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and3303_y0);
  and_gate and_gate_h_u_cla24_and3304_y0(h_u_cla24_and3303_y0, h_u_cla24_and3302_y0, h_u_cla24_and3304_y0);
  and_gate and_gate_h_u_cla24_and3305_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and3305_y0);
  and_gate and_gate_h_u_cla24_and3306_y0(h_u_cla24_and3305_y0, h_u_cla24_and3304_y0, h_u_cla24_and3306_y0);
  and_gate and_gate_h_u_cla24_and3307_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and3307_y0);
  and_gate and_gate_h_u_cla24_and3308_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and3308_y0);
  and_gate and_gate_h_u_cla24_and3309_y0(h_u_cla24_and3308_y0, h_u_cla24_and3307_y0, h_u_cla24_and3309_y0);
  and_gate and_gate_h_u_cla24_and3310_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and3310_y0);
  or_gate or_gate_h_u_cla24_or210_y0(h_u_cla24_and3310_y0, h_u_cla24_and2910_y0, h_u_cla24_or210_y0);
  or_gate or_gate_h_u_cla24_or211_y0(h_u_cla24_or210_y0, h_u_cla24_and2949_y0, h_u_cla24_or211_y0);
  or_gate or_gate_h_u_cla24_or212_y0(h_u_cla24_or211_y0, h_u_cla24_and2986_y0, h_u_cla24_or212_y0);
  or_gate or_gate_h_u_cla24_or213_y0(h_u_cla24_or212_y0, h_u_cla24_and3021_y0, h_u_cla24_or213_y0);
  or_gate or_gate_h_u_cla24_or214_y0(h_u_cla24_or213_y0, h_u_cla24_and3054_y0, h_u_cla24_or214_y0);
  or_gate or_gate_h_u_cla24_or215_y0(h_u_cla24_or214_y0, h_u_cla24_and3085_y0, h_u_cla24_or215_y0);
  or_gate or_gate_h_u_cla24_or216_y0(h_u_cla24_or215_y0, h_u_cla24_and3114_y0, h_u_cla24_or216_y0);
  or_gate or_gate_h_u_cla24_or217_y0(h_u_cla24_or216_y0, h_u_cla24_and3141_y0, h_u_cla24_or217_y0);
  or_gate or_gate_h_u_cla24_or218_y0(h_u_cla24_or217_y0, h_u_cla24_and3166_y0, h_u_cla24_or218_y0);
  or_gate or_gate_h_u_cla24_or219_y0(h_u_cla24_or218_y0, h_u_cla24_and3189_y0, h_u_cla24_or219_y0);
  or_gate or_gate_h_u_cla24_or220_y0(h_u_cla24_or219_y0, h_u_cla24_and3210_y0, h_u_cla24_or220_y0);
  or_gate or_gate_h_u_cla24_or221_y0(h_u_cla24_or220_y0, h_u_cla24_and3229_y0, h_u_cla24_or221_y0);
  or_gate or_gate_h_u_cla24_or222_y0(h_u_cla24_or221_y0, h_u_cla24_and3246_y0, h_u_cla24_or222_y0);
  or_gate or_gate_h_u_cla24_or223_y0(h_u_cla24_or222_y0, h_u_cla24_and3261_y0, h_u_cla24_or223_y0);
  or_gate or_gate_h_u_cla24_or224_y0(h_u_cla24_or223_y0, h_u_cla24_and3274_y0, h_u_cla24_or224_y0);
  or_gate or_gate_h_u_cla24_or225_y0(h_u_cla24_or224_y0, h_u_cla24_and3285_y0, h_u_cla24_or225_y0);
  or_gate or_gate_h_u_cla24_or226_y0(h_u_cla24_or225_y0, h_u_cla24_and3294_y0, h_u_cla24_or226_y0);
  or_gate or_gate_h_u_cla24_or227_y0(h_u_cla24_or226_y0, h_u_cla24_and3301_y0, h_u_cla24_or227_y0);
  or_gate or_gate_h_u_cla24_or228_y0(h_u_cla24_or227_y0, h_u_cla24_and3306_y0, h_u_cla24_or228_y0);
  or_gate or_gate_h_u_cla24_or229_y0(h_u_cla24_or228_y0, h_u_cla24_and3309_y0, h_u_cla24_or229_y0);
  or_gate or_gate_h_u_cla24_or230_y0(h_u_cla24_pg_logic20_y1, h_u_cla24_or229_y0, h_u_cla24_or230_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic21_y0(a_21, b_21, h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic21_y1, h_u_cla24_pg_logic21_y2);
  xor_gate xor_gate_h_u_cla24_xor21_y0(h_u_cla24_pg_logic21_y2, h_u_cla24_or230_y0, h_u_cla24_xor21_y0);
  and_gate and_gate_h_u_cla24_and3311_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and3311_y0);
  and_gate and_gate_h_u_cla24_and3312_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and3312_y0);
  and_gate and_gate_h_u_cla24_and3313_y0(h_u_cla24_and3312_y0, h_u_cla24_and3311_y0, h_u_cla24_and3313_y0);
  and_gate and_gate_h_u_cla24_and3314_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and3314_y0);
  and_gate and_gate_h_u_cla24_and3315_y0(h_u_cla24_and3314_y0, h_u_cla24_and3313_y0, h_u_cla24_and3315_y0);
  and_gate and_gate_h_u_cla24_and3316_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and3316_y0);
  and_gate and_gate_h_u_cla24_and3317_y0(h_u_cla24_and3316_y0, h_u_cla24_and3315_y0, h_u_cla24_and3317_y0);
  and_gate and_gate_h_u_cla24_and3318_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and3318_y0);
  and_gate and_gate_h_u_cla24_and3319_y0(h_u_cla24_and3318_y0, h_u_cla24_and3317_y0, h_u_cla24_and3319_y0);
  and_gate and_gate_h_u_cla24_and3320_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and3320_y0);
  and_gate and_gate_h_u_cla24_and3321_y0(h_u_cla24_and3320_y0, h_u_cla24_and3319_y0, h_u_cla24_and3321_y0);
  and_gate and_gate_h_u_cla24_and3322_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and3322_y0);
  and_gate and_gate_h_u_cla24_and3323_y0(h_u_cla24_and3322_y0, h_u_cla24_and3321_y0, h_u_cla24_and3323_y0);
  and_gate and_gate_h_u_cla24_and3324_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and3324_y0);
  and_gate and_gate_h_u_cla24_and3325_y0(h_u_cla24_and3324_y0, h_u_cla24_and3323_y0, h_u_cla24_and3325_y0);
  and_gate and_gate_h_u_cla24_and3326_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and3326_y0);
  and_gate and_gate_h_u_cla24_and3327_y0(h_u_cla24_and3326_y0, h_u_cla24_and3325_y0, h_u_cla24_and3327_y0);
  and_gate and_gate_h_u_cla24_and3328_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and3328_y0);
  and_gate and_gate_h_u_cla24_and3329_y0(h_u_cla24_and3328_y0, h_u_cla24_and3327_y0, h_u_cla24_and3329_y0);
  and_gate and_gate_h_u_cla24_and3330_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and3330_y0);
  and_gate and_gate_h_u_cla24_and3331_y0(h_u_cla24_and3330_y0, h_u_cla24_and3329_y0, h_u_cla24_and3331_y0);
  and_gate and_gate_h_u_cla24_and3332_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and3332_y0);
  and_gate and_gate_h_u_cla24_and3333_y0(h_u_cla24_and3332_y0, h_u_cla24_and3331_y0, h_u_cla24_and3333_y0);
  and_gate and_gate_h_u_cla24_and3334_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and3334_y0);
  and_gate and_gate_h_u_cla24_and3335_y0(h_u_cla24_and3334_y0, h_u_cla24_and3333_y0, h_u_cla24_and3335_y0);
  and_gate and_gate_h_u_cla24_and3336_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and3336_y0);
  and_gate and_gate_h_u_cla24_and3337_y0(h_u_cla24_and3336_y0, h_u_cla24_and3335_y0, h_u_cla24_and3337_y0);
  and_gate and_gate_h_u_cla24_and3338_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and3338_y0);
  and_gate and_gate_h_u_cla24_and3339_y0(h_u_cla24_and3338_y0, h_u_cla24_and3337_y0, h_u_cla24_and3339_y0);
  and_gate and_gate_h_u_cla24_and3340_y0(h_u_cla24_pg_logic15_y0, constant_wire_0, h_u_cla24_and3340_y0);
  and_gate and_gate_h_u_cla24_and3341_y0(h_u_cla24_and3340_y0, h_u_cla24_and3339_y0, h_u_cla24_and3341_y0);
  and_gate and_gate_h_u_cla24_and3342_y0(h_u_cla24_pg_logic16_y0, constant_wire_0, h_u_cla24_and3342_y0);
  and_gate and_gate_h_u_cla24_and3343_y0(h_u_cla24_and3342_y0, h_u_cla24_and3341_y0, h_u_cla24_and3343_y0);
  and_gate and_gate_h_u_cla24_and3344_y0(h_u_cla24_pg_logic17_y0, constant_wire_0, h_u_cla24_and3344_y0);
  and_gate and_gate_h_u_cla24_and3345_y0(h_u_cla24_and3344_y0, h_u_cla24_and3343_y0, h_u_cla24_and3345_y0);
  and_gate and_gate_h_u_cla24_and3346_y0(h_u_cla24_pg_logic18_y0, constant_wire_0, h_u_cla24_and3346_y0);
  and_gate and_gate_h_u_cla24_and3347_y0(h_u_cla24_and3346_y0, h_u_cla24_and3345_y0, h_u_cla24_and3347_y0);
  and_gate and_gate_h_u_cla24_and3348_y0(h_u_cla24_pg_logic19_y0, constant_wire_0, h_u_cla24_and3348_y0);
  and_gate and_gate_h_u_cla24_and3349_y0(h_u_cla24_and3348_y0, h_u_cla24_and3347_y0, h_u_cla24_and3349_y0);
  and_gate and_gate_h_u_cla24_and3350_y0(h_u_cla24_pg_logic20_y0, constant_wire_0, h_u_cla24_and3350_y0);
  and_gate and_gate_h_u_cla24_and3351_y0(h_u_cla24_and3350_y0, h_u_cla24_and3349_y0, h_u_cla24_and3351_y0);
  and_gate and_gate_h_u_cla24_and3352_y0(h_u_cla24_pg_logic21_y0, constant_wire_0, h_u_cla24_and3352_y0);
  and_gate and_gate_h_u_cla24_and3353_y0(h_u_cla24_and3352_y0, h_u_cla24_and3351_y0, h_u_cla24_and3353_y0);
  and_gate and_gate_h_u_cla24_and3354_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3354_y0);
  and_gate and_gate_h_u_cla24_and3355_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3355_y0);
  and_gate and_gate_h_u_cla24_and3356_y0(h_u_cla24_and3355_y0, h_u_cla24_and3354_y0, h_u_cla24_and3356_y0);
  and_gate and_gate_h_u_cla24_and3357_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3357_y0);
  and_gate and_gate_h_u_cla24_and3358_y0(h_u_cla24_and3357_y0, h_u_cla24_and3356_y0, h_u_cla24_and3358_y0);
  and_gate and_gate_h_u_cla24_and3359_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3359_y0);
  and_gate and_gate_h_u_cla24_and3360_y0(h_u_cla24_and3359_y0, h_u_cla24_and3358_y0, h_u_cla24_and3360_y0);
  and_gate and_gate_h_u_cla24_and3361_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3361_y0);
  and_gate and_gate_h_u_cla24_and3362_y0(h_u_cla24_and3361_y0, h_u_cla24_and3360_y0, h_u_cla24_and3362_y0);
  and_gate and_gate_h_u_cla24_and3363_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3363_y0);
  and_gate and_gate_h_u_cla24_and3364_y0(h_u_cla24_and3363_y0, h_u_cla24_and3362_y0, h_u_cla24_and3364_y0);
  and_gate and_gate_h_u_cla24_and3365_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3365_y0);
  and_gate and_gate_h_u_cla24_and3366_y0(h_u_cla24_and3365_y0, h_u_cla24_and3364_y0, h_u_cla24_and3366_y0);
  and_gate and_gate_h_u_cla24_and3367_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3367_y0);
  and_gate and_gate_h_u_cla24_and3368_y0(h_u_cla24_and3367_y0, h_u_cla24_and3366_y0, h_u_cla24_and3368_y0);
  and_gate and_gate_h_u_cla24_and3369_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3369_y0);
  and_gate and_gate_h_u_cla24_and3370_y0(h_u_cla24_and3369_y0, h_u_cla24_and3368_y0, h_u_cla24_and3370_y0);
  and_gate and_gate_h_u_cla24_and3371_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3371_y0);
  and_gate and_gate_h_u_cla24_and3372_y0(h_u_cla24_and3371_y0, h_u_cla24_and3370_y0, h_u_cla24_and3372_y0);
  and_gate and_gate_h_u_cla24_and3373_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3373_y0);
  and_gate and_gate_h_u_cla24_and3374_y0(h_u_cla24_and3373_y0, h_u_cla24_and3372_y0, h_u_cla24_and3374_y0);
  and_gate and_gate_h_u_cla24_and3375_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3375_y0);
  and_gate and_gate_h_u_cla24_and3376_y0(h_u_cla24_and3375_y0, h_u_cla24_and3374_y0, h_u_cla24_and3376_y0);
  and_gate and_gate_h_u_cla24_and3377_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3377_y0);
  and_gate and_gate_h_u_cla24_and3378_y0(h_u_cla24_and3377_y0, h_u_cla24_and3376_y0, h_u_cla24_and3378_y0);
  and_gate and_gate_h_u_cla24_and3379_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3379_y0);
  and_gate and_gate_h_u_cla24_and3380_y0(h_u_cla24_and3379_y0, h_u_cla24_and3378_y0, h_u_cla24_and3380_y0);
  and_gate and_gate_h_u_cla24_and3381_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3381_y0);
  and_gate and_gate_h_u_cla24_and3382_y0(h_u_cla24_and3381_y0, h_u_cla24_and3380_y0, h_u_cla24_and3382_y0);
  and_gate and_gate_h_u_cla24_and3383_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3383_y0);
  and_gate and_gate_h_u_cla24_and3384_y0(h_u_cla24_and3383_y0, h_u_cla24_and3382_y0, h_u_cla24_and3384_y0);
  and_gate and_gate_h_u_cla24_and3385_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3385_y0);
  and_gate and_gate_h_u_cla24_and3386_y0(h_u_cla24_and3385_y0, h_u_cla24_and3384_y0, h_u_cla24_and3386_y0);
  and_gate and_gate_h_u_cla24_and3387_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3387_y0);
  and_gate and_gate_h_u_cla24_and3388_y0(h_u_cla24_and3387_y0, h_u_cla24_and3386_y0, h_u_cla24_and3388_y0);
  and_gate and_gate_h_u_cla24_and3389_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3389_y0);
  and_gate and_gate_h_u_cla24_and3390_y0(h_u_cla24_and3389_y0, h_u_cla24_and3388_y0, h_u_cla24_and3390_y0);
  and_gate and_gate_h_u_cla24_and3391_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3391_y0);
  and_gate and_gate_h_u_cla24_and3392_y0(h_u_cla24_and3391_y0, h_u_cla24_and3390_y0, h_u_cla24_and3392_y0);
  and_gate and_gate_h_u_cla24_and3393_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3393_y0);
  and_gate and_gate_h_u_cla24_and3394_y0(h_u_cla24_and3393_y0, h_u_cla24_and3392_y0, h_u_cla24_and3394_y0);
  and_gate and_gate_h_u_cla24_and3395_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3395_y0);
  and_gate and_gate_h_u_cla24_and3396_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3396_y0);
  and_gate and_gate_h_u_cla24_and3397_y0(h_u_cla24_and3396_y0, h_u_cla24_and3395_y0, h_u_cla24_and3397_y0);
  and_gate and_gate_h_u_cla24_and3398_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3398_y0);
  and_gate and_gate_h_u_cla24_and3399_y0(h_u_cla24_and3398_y0, h_u_cla24_and3397_y0, h_u_cla24_and3399_y0);
  and_gate and_gate_h_u_cla24_and3400_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3400_y0);
  and_gate and_gate_h_u_cla24_and3401_y0(h_u_cla24_and3400_y0, h_u_cla24_and3399_y0, h_u_cla24_and3401_y0);
  and_gate and_gate_h_u_cla24_and3402_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3402_y0);
  and_gate and_gate_h_u_cla24_and3403_y0(h_u_cla24_and3402_y0, h_u_cla24_and3401_y0, h_u_cla24_and3403_y0);
  and_gate and_gate_h_u_cla24_and3404_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3404_y0);
  and_gate and_gate_h_u_cla24_and3405_y0(h_u_cla24_and3404_y0, h_u_cla24_and3403_y0, h_u_cla24_and3405_y0);
  and_gate and_gate_h_u_cla24_and3406_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3406_y0);
  and_gate and_gate_h_u_cla24_and3407_y0(h_u_cla24_and3406_y0, h_u_cla24_and3405_y0, h_u_cla24_and3407_y0);
  and_gate and_gate_h_u_cla24_and3408_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3408_y0);
  and_gate and_gate_h_u_cla24_and3409_y0(h_u_cla24_and3408_y0, h_u_cla24_and3407_y0, h_u_cla24_and3409_y0);
  and_gate and_gate_h_u_cla24_and3410_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3410_y0);
  and_gate and_gate_h_u_cla24_and3411_y0(h_u_cla24_and3410_y0, h_u_cla24_and3409_y0, h_u_cla24_and3411_y0);
  and_gate and_gate_h_u_cla24_and3412_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3412_y0);
  and_gate and_gate_h_u_cla24_and3413_y0(h_u_cla24_and3412_y0, h_u_cla24_and3411_y0, h_u_cla24_and3413_y0);
  and_gate and_gate_h_u_cla24_and3414_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3414_y0);
  and_gate and_gate_h_u_cla24_and3415_y0(h_u_cla24_and3414_y0, h_u_cla24_and3413_y0, h_u_cla24_and3415_y0);
  and_gate and_gate_h_u_cla24_and3416_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3416_y0);
  and_gate and_gate_h_u_cla24_and3417_y0(h_u_cla24_and3416_y0, h_u_cla24_and3415_y0, h_u_cla24_and3417_y0);
  and_gate and_gate_h_u_cla24_and3418_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3418_y0);
  and_gate and_gate_h_u_cla24_and3419_y0(h_u_cla24_and3418_y0, h_u_cla24_and3417_y0, h_u_cla24_and3419_y0);
  and_gate and_gate_h_u_cla24_and3420_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3420_y0);
  and_gate and_gate_h_u_cla24_and3421_y0(h_u_cla24_and3420_y0, h_u_cla24_and3419_y0, h_u_cla24_and3421_y0);
  and_gate and_gate_h_u_cla24_and3422_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3422_y0);
  and_gate and_gate_h_u_cla24_and3423_y0(h_u_cla24_and3422_y0, h_u_cla24_and3421_y0, h_u_cla24_and3423_y0);
  and_gate and_gate_h_u_cla24_and3424_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3424_y0);
  and_gate and_gate_h_u_cla24_and3425_y0(h_u_cla24_and3424_y0, h_u_cla24_and3423_y0, h_u_cla24_and3425_y0);
  and_gate and_gate_h_u_cla24_and3426_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3426_y0);
  and_gate and_gate_h_u_cla24_and3427_y0(h_u_cla24_and3426_y0, h_u_cla24_and3425_y0, h_u_cla24_and3427_y0);
  and_gate and_gate_h_u_cla24_and3428_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3428_y0);
  and_gate and_gate_h_u_cla24_and3429_y0(h_u_cla24_and3428_y0, h_u_cla24_and3427_y0, h_u_cla24_and3429_y0);
  and_gate and_gate_h_u_cla24_and3430_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3430_y0);
  and_gate and_gate_h_u_cla24_and3431_y0(h_u_cla24_and3430_y0, h_u_cla24_and3429_y0, h_u_cla24_and3431_y0);
  and_gate and_gate_h_u_cla24_and3432_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3432_y0);
  and_gate and_gate_h_u_cla24_and3433_y0(h_u_cla24_and3432_y0, h_u_cla24_and3431_y0, h_u_cla24_and3433_y0);
  and_gate and_gate_h_u_cla24_and3434_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3434_y0);
  and_gate and_gate_h_u_cla24_and3435_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3435_y0);
  and_gate and_gate_h_u_cla24_and3436_y0(h_u_cla24_and3435_y0, h_u_cla24_and3434_y0, h_u_cla24_and3436_y0);
  and_gate and_gate_h_u_cla24_and3437_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3437_y0);
  and_gate and_gate_h_u_cla24_and3438_y0(h_u_cla24_and3437_y0, h_u_cla24_and3436_y0, h_u_cla24_and3438_y0);
  and_gate and_gate_h_u_cla24_and3439_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3439_y0);
  and_gate and_gate_h_u_cla24_and3440_y0(h_u_cla24_and3439_y0, h_u_cla24_and3438_y0, h_u_cla24_and3440_y0);
  and_gate and_gate_h_u_cla24_and3441_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3441_y0);
  and_gate and_gate_h_u_cla24_and3442_y0(h_u_cla24_and3441_y0, h_u_cla24_and3440_y0, h_u_cla24_and3442_y0);
  and_gate and_gate_h_u_cla24_and3443_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3443_y0);
  and_gate and_gate_h_u_cla24_and3444_y0(h_u_cla24_and3443_y0, h_u_cla24_and3442_y0, h_u_cla24_and3444_y0);
  and_gate and_gate_h_u_cla24_and3445_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3445_y0);
  and_gate and_gate_h_u_cla24_and3446_y0(h_u_cla24_and3445_y0, h_u_cla24_and3444_y0, h_u_cla24_and3446_y0);
  and_gate and_gate_h_u_cla24_and3447_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3447_y0);
  and_gate and_gate_h_u_cla24_and3448_y0(h_u_cla24_and3447_y0, h_u_cla24_and3446_y0, h_u_cla24_and3448_y0);
  and_gate and_gate_h_u_cla24_and3449_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3449_y0);
  and_gate and_gate_h_u_cla24_and3450_y0(h_u_cla24_and3449_y0, h_u_cla24_and3448_y0, h_u_cla24_and3450_y0);
  and_gate and_gate_h_u_cla24_and3451_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3451_y0);
  and_gate and_gate_h_u_cla24_and3452_y0(h_u_cla24_and3451_y0, h_u_cla24_and3450_y0, h_u_cla24_and3452_y0);
  and_gate and_gate_h_u_cla24_and3453_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3453_y0);
  and_gate and_gate_h_u_cla24_and3454_y0(h_u_cla24_and3453_y0, h_u_cla24_and3452_y0, h_u_cla24_and3454_y0);
  and_gate and_gate_h_u_cla24_and3455_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3455_y0);
  and_gate and_gate_h_u_cla24_and3456_y0(h_u_cla24_and3455_y0, h_u_cla24_and3454_y0, h_u_cla24_and3456_y0);
  and_gate and_gate_h_u_cla24_and3457_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3457_y0);
  and_gate and_gate_h_u_cla24_and3458_y0(h_u_cla24_and3457_y0, h_u_cla24_and3456_y0, h_u_cla24_and3458_y0);
  and_gate and_gate_h_u_cla24_and3459_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3459_y0);
  and_gate and_gate_h_u_cla24_and3460_y0(h_u_cla24_and3459_y0, h_u_cla24_and3458_y0, h_u_cla24_and3460_y0);
  and_gate and_gate_h_u_cla24_and3461_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3461_y0);
  and_gate and_gate_h_u_cla24_and3462_y0(h_u_cla24_and3461_y0, h_u_cla24_and3460_y0, h_u_cla24_and3462_y0);
  and_gate and_gate_h_u_cla24_and3463_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3463_y0);
  and_gate and_gate_h_u_cla24_and3464_y0(h_u_cla24_and3463_y0, h_u_cla24_and3462_y0, h_u_cla24_and3464_y0);
  and_gate and_gate_h_u_cla24_and3465_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3465_y0);
  and_gate and_gate_h_u_cla24_and3466_y0(h_u_cla24_and3465_y0, h_u_cla24_and3464_y0, h_u_cla24_and3466_y0);
  and_gate and_gate_h_u_cla24_and3467_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3467_y0);
  and_gate and_gate_h_u_cla24_and3468_y0(h_u_cla24_and3467_y0, h_u_cla24_and3466_y0, h_u_cla24_and3468_y0);
  and_gate and_gate_h_u_cla24_and3469_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3469_y0);
  and_gate and_gate_h_u_cla24_and3470_y0(h_u_cla24_and3469_y0, h_u_cla24_and3468_y0, h_u_cla24_and3470_y0);
  and_gate and_gate_h_u_cla24_and3471_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3471_y0);
  and_gate and_gate_h_u_cla24_and3472_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3472_y0);
  and_gate and_gate_h_u_cla24_and3473_y0(h_u_cla24_and3472_y0, h_u_cla24_and3471_y0, h_u_cla24_and3473_y0);
  and_gate and_gate_h_u_cla24_and3474_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3474_y0);
  and_gate and_gate_h_u_cla24_and3475_y0(h_u_cla24_and3474_y0, h_u_cla24_and3473_y0, h_u_cla24_and3475_y0);
  and_gate and_gate_h_u_cla24_and3476_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3476_y0);
  and_gate and_gate_h_u_cla24_and3477_y0(h_u_cla24_and3476_y0, h_u_cla24_and3475_y0, h_u_cla24_and3477_y0);
  and_gate and_gate_h_u_cla24_and3478_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3478_y0);
  and_gate and_gate_h_u_cla24_and3479_y0(h_u_cla24_and3478_y0, h_u_cla24_and3477_y0, h_u_cla24_and3479_y0);
  and_gate and_gate_h_u_cla24_and3480_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3480_y0);
  and_gate and_gate_h_u_cla24_and3481_y0(h_u_cla24_and3480_y0, h_u_cla24_and3479_y0, h_u_cla24_and3481_y0);
  and_gate and_gate_h_u_cla24_and3482_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3482_y0);
  and_gate and_gate_h_u_cla24_and3483_y0(h_u_cla24_and3482_y0, h_u_cla24_and3481_y0, h_u_cla24_and3483_y0);
  and_gate and_gate_h_u_cla24_and3484_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3484_y0);
  and_gate and_gate_h_u_cla24_and3485_y0(h_u_cla24_and3484_y0, h_u_cla24_and3483_y0, h_u_cla24_and3485_y0);
  and_gate and_gate_h_u_cla24_and3486_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3486_y0);
  and_gate and_gate_h_u_cla24_and3487_y0(h_u_cla24_and3486_y0, h_u_cla24_and3485_y0, h_u_cla24_and3487_y0);
  and_gate and_gate_h_u_cla24_and3488_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3488_y0);
  and_gate and_gate_h_u_cla24_and3489_y0(h_u_cla24_and3488_y0, h_u_cla24_and3487_y0, h_u_cla24_and3489_y0);
  and_gate and_gate_h_u_cla24_and3490_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3490_y0);
  and_gate and_gate_h_u_cla24_and3491_y0(h_u_cla24_and3490_y0, h_u_cla24_and3489_y0, h_u_cla24_and3491_y0);
  and_gate and_gate_h_u_cla24_and3492_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3492_y0);
  and_gate and_gate_h_u_cla24_and3493_y0(h_u_cla24_and3492_y0, h_u_cla24_and3491_y0, h_u_cla24_and3493_y0);
  and_gate and_gate_h_u_cla24_and3494_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3494_y0);
  and_gate and_gate_h_u_cla24_and3495_y0(h_u_cla24_and3494_y0, h_u_cla24_and3493_y0, h_u_cla24_and3495_y0);
  and_gate and_gate_h_u_cla24_and3496_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3496_y0);
  and_gate and_gate_h_u_cla24_and3497_y0(h_u_cla24_and3496_y0, h_u_cla24_and3495_y0, h_u_cla24_and3497_y0);
  and_gate and_gate_h_u_cla24_and3498_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3498_y0);
  and_gate and_gate_h_u_cla24_and3499_y0(h_u_cla24_and3498_y0, h_u_cla24_and3497_y0, h_u_cla24_and3499_y0);
  and_gate and_gate_h_u_cla24_and3500_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3500_y0);
  and_gate and_gate_h_u_cla24_and3501_y0(h_u_cla24_and3500_y0, h_u_cla24_and3499_y0, h_u_cla24_and3501_y0);
  and_gate and_gate_h_u_cla24_and3502_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3502_y0);
  and_gate and_gate_h_u_cla24_and3503_y0(h_u_cla24_and3502_y0, h_u_cla24_and3501_y0, h_u_cla24_and3503_y0);
  and_gate and_gate_h_u_cla24_and3504_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3504_y0);
  and_gate and_gate_h_u_cla24_and3505_y0(h_u_cla24_and3504_y0, h_u_cla24_and3503_y0, h_u_cla24_and3505_y0);
  and_gate and_gate_h_u_cla24_and3506_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3506_y0);
  and_gate and_gate_h_u_cla24_and3507_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3507_y0);
  and_gate and_gate_h_u_cla24_and3508_y0(h_u_cla24_and3507_y0, h_u_cla24_and3506_y0, h_u_cla24_and3508_y0);
  and_gate and_gate_h_u_cla24_and3509_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3509_y0);
  and_gate and_gate_h_u_cla24_and3510_y0(h_u_cla24_and3509_y0, h_u_cla24_and3508_y0, h_u_cla24_and3510_y0);
  and_gate and_gate_h_u_cla24_and3511_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3511_y0);
  and_gate and_gate_h_u_cla24_and3512_y0(h_u_cla24_and3511_y0, h_u_cla24_and3510_y0, h_u_cla24_and3512_y0);
  and_gate and_gate_h_u_cla24_and3513_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3513_y0);
  and_gate and_gate_h_u_cla24_and3514_y0(h_u_cla24_and3513_y0, h_u_cla24_and3512_y0, h_u_cla24_and3514_y0);
  and_gate and_gate_h_u_cla24_and3515_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3515_y0);
  and_gate and_gate_h_u_cla24_and3516_y0(h_u_cla24_and3515_y0, h_u_cla24_and3514_y0, h_u_cla24_and3516_y0);
  and_gate and_gate_h_u_cla24_and3517_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3517_y0);
  and_gate and_gate_h_u_cla24_and3518_y0(h_u_cla24_and3517_y0, h_u_cla24_and3516_y0, h_u_cla24_and3518_y0);
  and_gate and_gate_h_u_cla24_and3519_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3519_y0);
  and_gate and_gate_h_u_cla24_and3520_y0(h_u_cla24_and3519_y0, h_u_cla24_and3518_y0, h_u_cla24_and3520_y0);
  and_gate and_gate_h_u_cla24_and3521_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3521_y0);
  and_gate and_gate_h_u_cla24_and3522_y0(h_u_cla24_and3521_y0, h_u_cla24_and3520_y0, h_u_cla24_and3522_y0);
  and_gate and_gate_h_u_cla24_and3523_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3523_y0);
  and_gate and_gate_h_u_cla24_and3524_y0(h_u_cla24_and3523_y0, h_u_cla24_and3522_y0, h_u_cla24_and3524_y0);
  and_gate and_gate_h_u_cla24_and3525_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3525_y0);
  and_gate and_gate_h_u_cla24_and3526_y0(h_u_cla24_and3525_y0, h_u_cla24_and3524_y0, h_u_cla24_and3526_y0);
  and_gate and_gate_h_u_cla24_and3527_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3527_y0);
  and_gate and_gate_h_u_cla24_and3528_y0(h_u_cla24_and3527_y0, h_u_cla24_and3526_y0, h_u_cla24_and3528_y0);
  and_gate and_gate_h_u_cla24_and3529_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3529_y0);
  and_gate and_gate_h_u_cla24_and3530_y0(h_u_cla24_and3529_y0, h_u_cla24_and3528_y0, h_u_cla24_and3530_y0);
  and_gate and_gate_h_u_cla24_and3531_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3531_y0);
  and_gate and_gate_h_u_cla24_and3532_y0(h_u_cla24_and3531_y0, h_u_cla24_and3530_y0, h_u_cla24_and3532_y0);
  and_gate and_gate_h_u_cla24_and3533_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3533_y0);
  and_gate and_gate_h_u_cla24_and3534_y0(h_u_cla24_and3533_y0, h_u_cla24_and3532_y0, h_u_cla24_and3534_y0);
  and_gate and_gate_h_u_cla24_and3535_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3535_y0);
  and_gate and_gate_h_u_cla24_and3536_y0(h_u_cla24_and3535_y0, h_u_cla24_and3534_y0, h_u_cla24_and3536_y0);
  and_gate and_gate_h_u_cla24_and3537_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and3537_y0);
  and_gate and_gate_h_u_cla24_and3538_y0(h_u_cla24_and3537_y0, h_u_cla24_and3536_y0, h_u_cla24_and3538_y0);
  and_gate and_gate_h_u_cla24_and3539_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3539_y0);
  and_gate and_gate_h_u_cla24_and3540_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3540_y0);
  and_gate and_gate_h_u_cla24_and3541_y0(h_u_cla24_and3540_y0, h_u_cla24_and3539_y0, h_u_cla24_and3541_y0);
  and_gate and_gate_h_u_cla24_and3542_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3542_y0);
  and_gate and_gate_h_u_cla24_and3543_y0(h_u_cla24_and3542_y0, h_u_cla24_and3541_y0, h_u_cla24_and3543_y0);
  and_gate and_gate_h_u_cla24_and3544_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3544_y0);
  and_gate and_gate_h_u_cla24_and3545_y0(h_u_cla24_and3544_y0, h_u_cla24_and3543_y0, h_u_cla24_and3545_y0);
  and_gate and_gate_h_u_cla24_and3546_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3546_y0);
  and_gate and_gate_h_u_cla24_and3547_y0(h_u_cla24_and3546_y0, h_u_cla24_and3545_y0, h_u_cla24_and3547_y0);
  and_gate and_gate_h_u_cla24_and3548_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3548_y0);
  and_gate and_gate_h_u_cla24_and3549_y0(h_u_cla24_and3548_y0, h_u_cla24_and3547_y0, h_u_cla24_and3549_y0);
  and_gate and_gate_h_u_cla24_and3550_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3550_y0);
  and_gate and_gate_h_u_cla24_and3551_y0(h_u_cla24_and3550_y0, h_u_cla24_and3549_y0, h_u_cla24_and3551_y0);
  and_gate and_gate_h_u_cla24_and3552_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3552_y0);
  and_gate and_gate_h_u_cla24_and3553_y0(h_u_cla24_and3552_y0, h_u_cla24_and3551_y0, h_u_cla24_and3553_y0);
  and_gate and_gate_h_u_cla24_and3554_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3554_y0);
  and_gate and_gate_h_u_cla24_and3555_y0(h_u_cla24_and3554_y0, h_u_cla24_and3553_y0, h_u_cla24_and3555_y0);
  and_gate and_gate_h_u_cla24_and3556_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3556_y0);
  and_gate and_gate_h_u_cla24_and3557_y0(h_u_cla24_and3556_y0, h_u_cla24_and3555_y0, h_u_cla24_and3557_y0);
  and_gate and_gate_h_u_cla24_and3558_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3558_y0);
  and_gate and_gate_h_u_cla24_and3559_y0(h_u_cla24_and3558_y0, h_u_cla24_and3557_y0, h_u_cla24_and3559_y0);
  and_gate and_gate_h_u_cla24_and3560_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3560_y0);
  and_gate and_gate_h_u_cla24_and3561_y0(h_u_cla24_and3560_y0, h_u_cla24_and3559_y0, h_u_cla24_and3561_y0);
  and_gate and_gate_h_u_cla24_and3562_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3562_y0);
  and_gate and_gate_h_u_cla24_and3563_y0(h_u_cla24_and3562_y0, h_u_cla24_and3561_y0, h_u_cla24_and3563_y0);
  and_gate and_gate_h_u_cla24_and3564_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3564_y0);
  and_gate and_gate_h_u_cla24_and3565_y0(h_u_cla24_and3564_y0, h_u_cla24_and3563_y0, h_u_cla24_and3565_y0);
  and_gate and_gate_h_u_cla24_and3566_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3566_y0);
  and_gate and_gate_h_u_cla24_and3567_y0(h_u_cla24_and3566_y0, h_u_cla24_and3565_y0, h_u_cla24_and3567_y0);
  and_gate and_gate_h_u_cla24_and3568_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and3568_y0);
  and_gate and_gate_h_u_cla24_and3569_y0(h_u_cla24_and3568_y0, h_u_cla24_and3567_y0, h_u_cla24_and3569_y0);
  and_gate and_gate_h_u_cla24_and3570_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3570_y0);
  and_gate and_gate_h_u_cla24_and3571_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3571_y0);
  and_gate and_gate_h_u_cla24_and3572_y0(h_u_cla24_and3571_y0, h_u_cla24_and3570_y0, h_u_cla24_and3572_y0);
  and_gate and_gate_h_u_cla24_and3573_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3573_y0);
  and_gate and_gate_h_u_cla24_and3574_y0(h_u_cla24_and3573_y0, h_u_cla24_and3572_y0, h_u_cla24_and3574_y0);
  and_gate and_gate_h_u_cla24_and3575_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3575_y0);
  and_gate and_gate_h_u_cla24_and3576_y0(h_u_cla24_and3575_y0, h_u_cla24_and3574_y0, h_u_cla24_and3576_y0);
  and_gate and_gate_h_u_cla24_and3577_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3577_y0);
  and_gate and_gate_h_u_cla24_and3578_y0(h_u_cla24_and3577_y0, h_u_cla24_and3576_y0, h_u_cla24_and3578_y0);
  and_gate and_gate_h_u_cla24_and3579_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3579_y0);
  and_gate and_gate_h_u_cla24_and3580_y0(h_u_cla24_and3579_y0, h_u_cla24_and3578_y0, h_u_cla24_and3580_y0);
  and_gate and_gate_h_u_cla24_and3581_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3581_y0);
  and_gate and_gate_h_u_cla24_and3582_y0(h_u_cla24_and3581_y0, h_u_cla24_and3580_y0, h_u_cla24_and3582_y0);
  and_gate and_gate_h_u_cla24_and3583_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3583_y0);
  and_gate and_gate_h_u_cla24_and3584_y0(h_u_cla24_and3583_y0, h_u_cla24_and3582_y0, h_u_cla24_and3584_y0);
  and_gate and_gate_h_u_cla24_and3585_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3585_y0);
  and_gate and_gate_h_u_cla24_and3586_y0(h_u_cla24_and3585_y0, h_u_cla24_and3584_y0, h_u_cla24_and3586_y0);
  and_gate and_gate_h_u_cla24_and3587_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3587_y0);
  and_gate and_gate_h_u_cla24_and3588_y0(h_u_cla24_and3587_y0, h_u_cla24_and3586_y0, h_u_cla24_and3588_y0);
  and_gate and_gate_h_u_cla24_and3589_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3589_y0);
  and_gate and_gate_h_u_cla24_and3590_y0(h_u_cla24_and3589_y0, h_u_cla24_and3588_y0, h_u_cla24_and3590_y0);
  and_gate and_gate_h_u_cla24_and3591_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3591_y0);
  and_gate and_gate_h_u_cla24_and3592_y0(h_u_cla24_and3591_y0, h_u_cla24_and3590_y0, h_u_cla24_and3592_y0);
  and_gate and_gate_h_u_cla24_and3593_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3593_y0);
  and_gate and_gate_h_u_cla24_and3594_y0(h_u_cla24_and3593_y0, h_u_cla24_and3592_y0, h_u_cla24_and3594_y0);
  and_gate and_gate_h_u_cla24_and3595_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3595_y0);
  and_gate and_gate_h_u_cla24_and3596_y0(h_u_cla24_and3595_y0, h_u_cla24_and3594_y0, h_u_cla24_and3596_y0);
  and_gate and_gate_h_u_cla24_and3597_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and3597_y0);
  and_gate and_gate_h_u_cla24_and3598_y0(h_u_cla24_and3597_y0, h_u_cla24_and3596_y0, h_u_cla24_and3598_y0);
  and_gate and_gate_h_u_cla24_and3599_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3599_y0);
  and_gate and_gate_h_u_cla24_and3600_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3600_y0);
  and_gate and_gate_h_u_cla24_and3601_y0(h_u_cla24_and3600_y0, h_u_cla24_and3599_y0, h_u_cla24_and3601_y0);
  and_gate and_gate_h_u_cla24_and3602_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3602_y0);
  and_gate and_gate_h_u_cla24_and3603_y0(h_u_cla24_and3602_y0, h_u_cla24_and3601_y0, h_u_cla24_and3603_y0);
  and_gate and_gate_h_u_cla24_and3604_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3604_y0);
  and_gate and_gate_h_u_cla24_and3605_y0(h_u_cla24_and3604_y0, h_u_cla24_and3603_y0, h_u_cla24_and3605_y0);
  and_gate and_gate_h_u_cla24_and3606_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3606_y0);
  and_gate and_gate_h_u_cla24_and3607_y0(h_u_cla24_and3606_y0, h_u_cla24_and3605_y0, h_u_cla24_and3607_y0);
  and_gate and_gate_h_u_cla24_and3608_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3608_y0);
  and_gate and_gate_h_u_cla24_and3609_y0(h_u_cla24_and3608_y0, h_u_cla24_and3607_y0, h_u_cla24_and3609_y0);
  and_gate and_gate_h_u_cla24_and3610_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3610_y0);
  and_gate and_gate_h_u_cla24_and3611_y0(h_u_cla24_and3610_y0, h_u_cla24_and3609_y0, h_u_cla24_and3611_y0);
  and_gate and_gate_h_u_cla24_and3612_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3612_y0);
  and_gate and_gate_h_u_cla24_and3613_y0(h_u_cla24_and3612_y0, h_u_cla24_and3611_y0, h_u_cla24_and3613_y0);
  and_gate and_gate_h_u_cla24_and3614_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3614_y0);
  and_gate and_gate_h_u_cla24_and3615_y0(h_u_cla24_and3614_y0, h_u_cla24_and3613_y0, h_u_cla24_and3615_y0);
  and_gate and_gate_h_u_cla24_and3616_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3616_y0);
  and_gate and_gate_h_u_cla24_and3617_y0(h_u_cla24_and3616_y0, h_u_cla24_and3615_y0, h_u_cla24_and3617_y0);
  and_gate and_gate_h_u_cla24_and3618_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3618_y0);
  and_gate and_gate_h_u_cla24_and3619_y0(h_u_cla24_and3618_y0, h_u_cla24_and3617_y0, h_u_cla24_and3619_y0);
  and_gate and_gate_h_u_cla24_and3620_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3620_y0);
  and_gate and_gate_h_u_cla24_and3621_y0(h_u_cla24_and3620_y0, h_u_cla24_and3619_y0, h_u_cla24_and3621_y0);
  and_gate and_gate_h_u_cla24_and3622_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3622_y0);
  and_gate and_gate_h_u_cla24_and3623_y0(h_u_cla24_and3622_y0, h_u_cla24_and3621_y0, h_u_cla24_and3623_y0);
  and_gate and_gate_h_u_cla24_and3624_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and3624_y0);
  and_gate and_gate_h_u_cla24_and3625_y0(h_u_cla24_and3624_y0, h_u_cla24_and3623_y0, h_u_cla24_and3625_y0);
  and_gate and_gate_h_u_cla24_and3626_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3626_y0);
  and_gate and_gate_h_u_cla24_and3627_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3627_y0);
  and_gate and_gate_h_u_cla24_and3628_y0(h_u_cla24_and3627_y0, h_u_cla24_and3626_y0, h_u_cla24_and3628_y0);
  and_gate and_gate_h_u_cla24_and3629_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3629_y0);
  and_gate and_gate_h_u_cla24_and3630_y0(h_u_cla24_and3629_y0, h_u_cla24_and3628_y0, h_u_cla24_and3630_y0);
  and_gate and_gate_h_u_cla24_and3631_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3631_y0);
  and_gate and_gate_h_u_cla24_and3632_y0(h_u_cla24_and3631_y0, h_u_cla24_and3630_y0, h_u_cla24_and3632_y0);
  and_gate and_gate_h_u_cla24_and3633_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3633_y0);
  and_gate and_gate_h_u_cla24_and3634_y0(h_u_cla24_and3633_y0, h_u_cla24_and3632_y0, h_u_cla24_and3634_y0);
  and_gate and_gate_h_u_cla24_and3635_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3635_y0);
  and_gate and_gate_h_u_cla24_and3636_y0(h_u_cla24_and3635_y0, h_u_cla24_and3634_y0, h_u_cla24_and3636_y0);
  and_gate and_gate_h_u_cla24_and3637_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3637_y0);
  and_gate and_gate_h_u_cla24_and3638_y0(h_u_cla24_and3637_y0, h_u_cla24_and3636_y0, h_u_cla24_and3638_y0);
  and_gate and_gate_h_u_cla24_and3639_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3639_y0);
  and_gate and_gate_h_u_cla24_and3640_y0(h_u_cla24_and3639_y0, h_u_cla24_and3638_y0, h_u_cla24_and3640_y0);
  and_gate and_gate_h_u_cla24_and3641_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3641_y0);
  and_gate and_gate_h_u_cla24_and3642_y0(h_u_cla24_and3641_y0, h_u_cla24_and3640_y0, h_u_cla24_and3642_y0);
  and_gate and_gate_h_u_cla24_and3643_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3643_y0);
  and_gate and_gate_h_u_cla24_and3644_y0(h_u_cla24_and3643_y0, h_u_cla24_and3642_y0, h_u_cla24_and3644_y0);
  and_gate and_gate_h_u_cla24_and3645_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3645_y0);
  and_gate and_gate_h_u_cla24_and3646_y0(h_u_cla24_and3645_y0, h_u_cla24_and3644_y0, h_u_cla24_and3646_y0);
  and_gate and_gate_h_u_cla24_and3647_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3647_y0);
  and_gate and_gate_h_u_cla24_and3648_y0(h_u_cla24_and3647_y0, h_u_cla24_and3646_y0, h_u_cla24_and3648_y0);
  and_gate and_gate_h_u_cla24_and3649_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and3649_y0);
  and_gate and_gate_h_u_cla24_and3650_y0(h_u_cla24_and3649_y0, h_u_cla24_and3648_y0, h_u_cla24_and3650_y0);
  and_gate and_gate_h_u_cla24_and3651_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3651_y0);
  and_gate and_gate_h_u_cla24_and3652_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3652_y0);
  and_gate and_gate_h_u_cla24_and3653_y0(h_u_cla24_and3652_y0, h_u_cla24_and3651_y0, h_u_cla24_and3653_y0);
  and_gate and_gate_h_u_cla24_and3654_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3654_y0);
  and_gate and_gate_h_u_cla24_and3655_y0(h_u_cla24_and3654_y0, h_u_cla24_and3653_y0, h_u_cla24_and3655_y0);
  and_gate and_gate_h_u_cla24_and3656_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3656_y0);
  and_gate and_gate_h_u_cla24_and3657_y0(h_u_cla24_and3656_y0, h_u_cla24_and3655_y0, h_u_cla24_and3657_y0);
  and_gate and_gate_h_u_cla24_and3658_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3658_y0);
  and_gate and_gate_h_u_cla24_and3659_y0(h_u_cla24_and3658_y0, h_u_cla24_and3657_y0, h_u_cla24_and3659_y0);
  and_gate and_gate_h_u_cla24_and3660_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3660_y0);
  and_gate and_gate_h_u_cla24_and3661_y0(h_u_cla24_and3660_y0, h_u_cla24_and3659_y0, h_u_cla24_and3661_y0);
  and_gate and_gate_h_u_cla24_and3662_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3662_y0);
  and_gate and_gate_h_u_cla24_and3663_y0(h_u_cla24_and3662_y0, h_u_cla24_and3661_y0, h_u_cla24_and3663_y0);
  and_gate and_gate_h_u_cla24_and3664_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3664_y0);
  and_gate and_gate_h_u_cla24_and3665_y0(h_u_cla24_and3664_y0, h_u_cla24_and3663_y0, h_u_cla24_and3665_y0);
  and_gate and_gate_h_u_cla24_and3666_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3666_y0);
  and_gate and_gate_h_u_cla24_and3667_y0(h_u_cla24_and3666_y0, h_u_cla24_and3665_y0, h_u_cla24_and3667_y0);
  and_gate and_gate_h_u_cla24_and3668_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3668_y0);
  and_gate and_gate_h_u_cla24_and3669_y0(h_u_cla24_and3668_y0, h_u_cla24_and3667_y0, h_u_cla24_and3669_y0);
  and_gate and_gate_h_u_cla24_and3670_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3670_y0);
  and_gate and_gate_h_u_cla24_and3671_y0(h_u_cla24_and3670_y0, h_u_cla24_and3669_y0, h_u_cla24_and3671_y0);
  and_gate and_gate_h_u_cla24_and3672_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and3672_y0);
  and_gate and_gate_h_u_cla24_and3673_y0(h_u_cla24_and3672_y0, h_u_cla24_and3671_y0, h_u_cla24_and3673_y0);
  and_gate and_gate_h_u_cla24_and3674_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3674_y0);
  and_gate and_gate_h_u_cla24_and3675_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3675_y0);
  and_gate and_gate_h_u_cla24_and3676_y0(h_u_cla24_and3675_y0, h_u_cla24_and3674_y0, h_u_cla24_and3676_y0);
  and_gate and_gate_h_u_cla24_and3677_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3677_y0);
  and_gate and_gate_h_u_cla24_and3678_y0(h_u_cla24_and3677_y0, h_u_cla24_and3676_y0, h_u_cla24_and3678_y0);
  and_gate and_gate_h_u_cla24_and3679_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3679_y0);
  and_gate and_gate_h_u_cla24_and3680_y0(h_u_cla24_and3679_y0, h_u_cla24_and3678_y0, h_u_cla24_and3680_y0);
  and_gate and_gate_h_u_cla24_and3681_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3681_y0);
  and_gate and_gate_h_u_cla24_and3682_y0(h_u_cla24_and3681_y0, h_u_cla24_and3680_y0, h_u_cla24_and3682_y0);
  and_gate and_gate_h_u_cla24_and3683_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3683_y0);
  and_gate and_gate_h_u_cla24_and3684_y0(h_u_cla24_and3683_y0, h_u_cla24_and3682_y0, h_u_cla24_and3684_y0);
  and_gate and_gate_h_u_cla24_and3685_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3685_y0);
  and_gate and_gate_h_u_cla24_and3686_y0(h_u_cla24_and3685_y0, h_u_cla24_and3684_y0, h_u_cla24_and3686_y0);
  and_gate and_gate_h_u_cla24_and3687_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3687_y0);
  and_gate and_gate_h_u_cla24_and3688_y0(h_u_cla24_and3687_y0, h_u_cla24_and3686_y0, h_u_cla24_and3688_y0);
  and_gate and_gate_h_u_cla24_and3689_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3689_y0);
  and_gate and_gate_h_u_cla24_and3690_y0(h_u_cla24_and3689_y0, h_u_cla24_and3688_y0, h_u_cla24_and3690_y0);
  and_gate and_gate_h_u_cla24_and3691_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3691_y0);
  and_gate and_gate_h_u_cla24_and3692_y0(h_u_cla24_and3691_y0, h_u_cla24_and3690_y0, h_u_cla24_and3692_y0);
  and_gate and_gate_h_u_cla24_and3693_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and3693_y0);
  and_gate and_gate_h_u_cla24_and3694_y0(h_u_cla24_and3693_y0, h_u_cla24_and3692_y0, h_u_cla24_and3694_y0);
  and_gate and_gate_h_u_cla24_and3695_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3695_y0);
  and_gate and_gate_h_u_cla24_and3696_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3696_y0);
  and_gate and_gate_h_u_cla24_and3697_y0(h_u_cla24_and3696_y0, h_u_cla24_and3695_y0, h_u_cla24_and3697_y0);
  and_gate and_gate_h_u_cla24_and3698_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3698_y0);
  and_gate and_gate_h_u_cla24_and3699_y0(h_u_cla24_and3698_y0, h_u_cla24_and3697_y0, h_u_cla24_and3699_y0);
  and_gate and_gate_h_u_cla24_and3700_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3700_y0);
  and_gate and_gate_h_u_cla24_and3701_y0(h_u_cla24_and3700_y0, h_u_cla24_and3699_y0, h_u_cla24_and3701_y0);
  and_gate and_gate_h_u_cla24_and3702_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3702_y0);
  and_gate and_gate_h_u_cla24_and3703_y0(h_u_cla24_and3702_y0, h_u_cla24_and3701_y0, h_u_cla24_and3703_y0);
  and_gate and_gate_h_u_cla24_and3704_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3704_y0);
  and_gate and_gate_h_u_cla24_and3705_y0(h_u_cla24_and3704_y0, h_u_cla24_and3703_y0, h_u_cla24_and3705_y0);
  and_gate and_gate_h_u_cla24_and3706_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3706_y0);
  and_gate and_gate_h_u_cla24_and3707_y0(h_u_cla24_and3706_y0, h_u_cla24_and3705_y0, h_u_cla24_and3707_y0);
  and_gate and_gate_h_u_cla24_and3708_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3708_y0);
  and_gate and_gate_h_u_cla24_and3709_y0(h_u_cla24_and3708_y0, h_u_cla24_and3707_y0, h_u_cla24_and3709_y0);
  and_gate and_gate_h_u_cla24_and3710_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3710_y0);
  and_gate and_gate_h_u_cla24_and3711_y0(h_u_cla24_and3710_y0, h_u_cla24_and3709_y0, h_u_cla24_and3711_y0);
  and_gate and_gate_h_u_cla24_and3712_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and3712_y0);
  and_gate and_gate_h_u_cla24_and3713_y0(h_u_cla24_and3712_y0, h_u_cla24_and3711_y0, h_u_cla24_and3713_y0);
  and_gate and_gate_h_u_cla24_and3714_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3714_y0);
  and_gate and_gate_h_u_cla24_and3715_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3715_y0);
  and_gate and_gate_h_u_cla24_and3716_y0(h_u_cla24_and3715_y0, h_u_cla24_and3714_y0, h_u_cla24_and3716_y0);
  and_gate and_gate_h_u_cla24_and3717_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3717_y0);
  and_gate and_gate_h_u_cla24_and3718_y0(h_u_cla24_and3717_y0, h_u_cla24_and3716_y0, h_u_cla24_and3718_y0);
  and_gate and_gate_h_u_cla24_and3719_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3719_y0);
  and_gate and_gate_h_u_cla24_and3720_y0(h_u_cla24_and3719_y0, h_u_cla24_and3718_y0, h_u_cla24_and3720_y0);
  and_gate and_gate_h_u_cla24_and3721_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3721_y0);
  and_gate and_gate_h_u_cla24_and3722_y0(h_u_cla24_and3721_y0, h_u_cla24_and3720_y0, h_u_cla24_and3722_y0);
  and_gate and_gate_h_u_cla24_and3723_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3723_y0);
  and_gate and_gate_h_u_cla24_and3724_y0(h_u_cla24_and3723_y0, h_u_cla24_and3722_y0, h_u_cla24_and3724_y0);
  and_gate and_gate_h_u_cla24_and3725_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3725_y0);
  and_gate and_gate_h_u_cla24_and3726_y0(h_u_cla24_and3725_y0, h_u_cla24_and3724_y0, h_u_cla24_and3726_y0);
  and_gate and_gate_h_u_cla24_and3727_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3727_y0);
  and_gate and_gate_h_u_cla24_and3728_y0(h_u_cla24_and3727_y0, h_u_cla24_and3726_y0, h_u_cla24_and3728_y0);
  and_gate and_gate_h_u_cla24_and3729_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and3729_y0);
  and_gate and_gate_h_u_cla24_and3730_y0(h_u_cla24_and3729_y0, h_u_cla24_and3728_y0, h_u_cla24_and3730_y0);
  and_gate and_gate_h_u_cla24_and3731_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3731_y0);
  and_gate and_gate_h_u_cla24_and3732_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3732_y0);
  and_gate and_gate_h_u_cla24_and3733_y0(h_u_cla24_and3732_y0, h_u_cla24_and3731_y0, h_u_cla24_and3733_y0);
  and_gate and_gate_h_u_cla24_and3734_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3734_y0);
  and_gate and_gate_h_u_cla24_and3735_y0(h_u_cla24_and3734_y0, h_u_cla24_and3733_y0, h_u_cla24_and3735_y0);
  and_gate and_gate_h_u_cla24_and3736_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3736_y0);
  and_gate and_gate_h_u_cla24_and3737_y0(h_u_cla24_and3736_y0, h_u_cla24_and3735_y0, h_u_cla24_and3737_y0);
  and_gate and_gate_h_u_cla24_and3738_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3738_y0);
  and_gate and_gate_h_u_cla24_and3739_y0(h_u_cla24_and3738_y0, h_u_cla24_and3737_y0, h_u_cla24_and3739_y0);
  and_gate and_gate_h_u_cla24_and3740_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3740_y0);
  and_gate and_gate_h_u_cla24_and3741_y0(h_u_cla24_and3740_y0, h_u_cla24_and3739_y0, h_u_cla24_and3741_y0);
  and_gate and_gate_h_u_cla24_and3742_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3742_y0);
  and_gate and_gate_h_u_cla24_and3743_y0(h_u_cla24_and3742_y0, h_u_cla24_and3741_y0, h_u_cla24_and3743_y0);
  and_gate and_gate_h_u_cla24_and3744_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and3744_y0);
  and_gate and_gate_h_u_cla24_and3745_y0(h_u_cla24_and3744_y0, h_u_cla24_and3743_y0, h_u_cla24_and3745_y0);
  and_gate and_gate_h_u_cla24_and3746_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3746_y0);
  and_gate and_gate_h_u_cla24_and3747_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3747_y0);
  and_gate and_gate_h_u_cla24_and3748_y0(h_u_cla24_and3747_y0, h_u_cla24_and3746_y0, h_u_cla24_and3748_y0);
  and_gate and_gate_h_u_cla24_and3749_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3749_y0);
  and_gate and_gate_h_u_cla24_and3750_y0(h_u_cla24_and3749_y0, h_u_cla24_and3748_y0, h_u_cla24_and3750_y0);
  and_gate and_gate_h_u_cla24_and3751_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3751_y0);
  and_gate and_gate_h_u_cla24_and3752_y0(h_u_cla24_and3751_y0, h_u_cla24_and3750_y0, h_u_cla24_and3752_y0);
  and_gate and_gate_h_u_cla24_and3753_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3753_y0);
  and_gate and_gate_h_u_cla24_and3754_y0(h_u_cla24_and3753_y0, h_u_cla24_and3752_y0, h_u_cla24_and3754_y0);
  and_gate and_gate_h_u_cla24_and3755_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3755_y0);
  and_gate and_gate_h_u_cla24_and3756_y0(h_u_cla24_and3755_y0, h_u_cla24_and3754_y0, h_u_cla24_and3756_y0);
  and_gate and_gate_h_u_cla24_and3757_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and3757_y0);
  and_gate and_gate_h_u_cla24_and3758_y0(h_u_cla24_and3757_y0, h_u_cla24_and3756_y0, h_u_cla24_and3758_y0);
  and_gate and_gate_h_u_cla24_and3759_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3759_y0);
  and_gate and_gate_h_u_cla24_and3760_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3760_y0);
  and_gate and_gate_h_u_cla24_and3761_y0(h_u_cla24_and3760_y0, h_u_cla24_and3759_y0, h_u_cla24_and3761_y0);
  and_gate and_gate_h_u_cla24_and3762_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3762_y0);
  and_gate and_gate_h_u_cla24_and3763_y0(h_u_cla24_and3762_y0, h_u_cla24_and3761_y0, h_u_cla24_and3763_y0);
  and_gate and_gate_h_u_cla24_and3764_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3764_y0);
  and_gate and_gate_h_u_cla24_and3765_y0(h_u_cla24_and3764_y0, h_u_cla24_and3763_y0, h_u_cla24_and3765_y0);
  and_gate and_gate_h_u_cla24_and3766_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3766_y0);
  and_gate and_gate_h_u_cla24_and3767_y0(h_u_cla24_and3766_y0, h_u_cla24_and3765_y0, h_u_cla24_and3767_y0);
  and_gate and_gate_h_u_cla24_and3768_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and3768_y0);
  and_gate and_gate_h_u_cla24_and3769_y0(h_u_cla24_and3768_y0, h_u_cla24_and3767_y0, h_u_cla24_and3769_y0);
  and_gate and_gate_h_u_cla24_and3770_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and3770_y0);
  and_gate and_gate_h_u_cla24_and3771_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and3771_y0);
  and_gate and_gate_h_u_cla24_and3772_y0(h_u_cla24_and3771_y0, h_u_cla24_and3770_y0, h_u_cla24_and3772_y0);
  and_gate and_gate_h_u_cla24_and3773_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and3773_y0);
  and_gate and_gate_h_u_cla24_and3774_y0(h_u_cla24_and3773_y0, h_u_cla24_and3772_y0, h_u_cla24_and3774_y0);
  and_gate and_gate_h_u_cla24_and3775_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and3775_y0);
  and_gate and_gate_h_u_cla24_and3776_y0(h_u_cla24_and3775_y0, h_u_cla24_and3774_y0, h_u_cla24_and3776_y0);
  and_gate and_gate_h_u_cla24_and3777_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and3777_y0);
  and_gate and_gate_h_u_cla24_and3778_y0(h_u_cla24_and3777_y0, h_u_cla24_and3776_y0, h_u_cla24_and3778_y0);
  and_gate and_gate_h_u_cla24_and3779_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and3779_y0);
  and_gate and_gate_h_u_cla24_and3780_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and3780_y0);
  and_gate and_gate_h_u_cla24_and3781_y0(h_u_cla24_and3780_y0, h_u_cla24_and3779_y0, h_u_cla24_and3781_y0);
  and_gate and_gate_h_u_cla24_and3782_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and3782_y0);
  and_gate and_gate_h_u_cla24_and3783_y0(h_u_cla24_and3782_y0, h_u_cla24_and3781_y0, h_u_cla24_and3783_y0);
  and_gate and_gate_h_u_cla24_and3784_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and3784_y0);
  and_gate and_gate_h_u_cla24_and3785_y0(h_u_cla24_and3784_y0, h_u_cla24_and3783_y0, h_u_cla24_and3785_y0);
  and_gate and_gate_h_u_cla24_and3786_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and3786_y0);
  and_gate and_gate_h_u_cla24_and3787_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and3787_y0);
  and_gate and_gate_h_u_cla24_and3788_y0(h_u_cla24_and3787_y0, h_u_cla24_and3786_y0, h_u_cla24_and3788_y0);
  and_gate and_gate_h_u_cla24_and3789_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and3789_y0);
  and_gate and_gate_h_u_cla24_and3790_y0(h_u_cla24_and3789_y0, h_u_cla24_and3788_y0, h_u_cla24_and3790_y0);
  and_gate and_gate_h_u_cla24_and3791_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and3791_y0);
  and_gate and_gate_h_u_cla24_and3792_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and3792_y0);
  and_gate and_gate_h_u_cla24_and3793_y0(h_u_cla24_and3792_y0, h_u_cla24_and3791_y0, h_u_cla24_and3793_y0);
  and_gate and_gate_h_u_cla24_and3794_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic20_y1, h_u_cla24_and3794_y0);
  or_gate or_gate_h_u_cla24_or231_y0(h_u_cla24_and3794_y0, h_u_cla24_and3353_y0, h_u_cla24_or231_y0);
  or_gate or_gate_h_u_cla24_or232_y0(h_u_cla24_or231_y0, h_u_cla24_and3394_y0, h_u_cla24_or232_y0);
  or_gate or_gate_h_u_cla24_or233_y0(h_u_cla24_or232_y0, h_u_cla24_and3433_y0, h_u_cla24_or233_y0);
  or_gate or_gate_h_u_cla24_or234_y0(h_u_cla24_or233_y0, h_u_cla24_and3470_y0, h_u_cla24_or234_y0);
  or_gate or_gate_h_u_cla24_or235_y0(h_u_cla24_or234_y0, h_u_cla24_and3505_y0, h_u_cla24_or235_y0);
  or_gate or_gate_h_u_cla24_or236_y0(h_u_cla24_or235_y0, h_u_cla24_and3538_y0, h_u_cla24_or236_y0);
  or_gate or_gate_h_u_cla24_or237_y0(h_u_cla24_or236_y0, h_u_cla24_and3569_y0, h_u_cla24_or237_y0);
  or_gate or_gate_h_u_cla24_or238_y0(h_u_cla24_or237_y0, h_u_cla24_and3598_y0, h_u_cla24_or238_y0);
  or_gate or_gate_h_u_cla24_or239_y0(h_u_cla24_or238_y0, h_u_cla24_and3625_y0, h_u_cla24_or239_y0);
  or_gate or_gate_h_u_cla24_or240_y0(h_u_cla24_or239_y0, h_u_cla24_and3650_y0, h_u_cla24_or240_y0);
  or_gate or_gate_h_u_cla24_or241_y0(h_u_cla24_or240_y0, h_u_cla24_and3673_y0, h_u_cla24_or241_y0);
  or_gate or_gate_h_u_cla24_or242_y0(h_u_cla24_or241_y0, h_u_cla24_and3694_y0, h_u_cla24_or242_y0);
  or_gate or_gate_h_u_cla24_or243_y0(h_u_cla24_or242_y0, h_u_cla24_and3713_y0, h_u_cla24_or243_y0);
  or_gate or_gate_h_u_cla24_or244_y0(h_u_cla24_or243_y0, h_u_cla24_and3730_y0, h_u_cla24_or244_y0);
  or_gate or_gate_h_u_cla24_or245_y0(h_u_cla24_or244_y0, h_u_cla24_and3745_y0, h_u_cla24_or245_y0);
  or_gate or_gate_h_u_cla24_or246_y0(h_u_cla24_or245_y0, h_u_cla24_and3758_y0, h_u_cla24_or246_y0);
  or_gate or_gate_h_u_cla24_or247_y0(h_u_cla24_or246_y0, h_u_cla24_and3769_y0, h_u_cla24_or247_y0);
  or_gate or_gate_h_u_cla24_or248_y0(h_u_cla24_or247_y0, h_u_cla24_and3778_y0, h_u_cla24_or248_y0);
  or_gate or_gate_h_u_cla24_or249_y0(h_u_cla24_or248_y0, h_u_cla24_and3785_y0, h_u_cla24_or249_y0);
  or_gate or_gate_h_u_cla24_or250_y0(h_u_cla24_or249_y0, h_u_cla24_and3790_y0, h_u_cla24_or250_y0);
  or_gate or_gate_h_u_cla24_or251_y0(h_u_cla24_or250_y0, h_u_cla24_and3793_y0, h_u_cla24_or251_y0);
  or_gate or_gate_h_u_cla24_or252_y0(h_u_cla24_pg_logic21_y1, h_u_cla24_or251_y0, h_u_cla24_or252_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic22_y0(a_22, b_22, h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic22_y1, h_u_cla24_pg_logic22_y2);
  xor_gate xor_gate_h_u_cla24_xor22_y0(h_u_cla24_pg_logic22_y2, h_u_cla24_or252_y0, h_u_cla24_xor22_y0);
  and_gate and_gate_h_u_cla24_and3795_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and3795_y0);
  and_gate and_gate_h_u_cla24_and3796_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and3796_y0);
  and_gate and_gate_h_u_cla24_and3797_y0(h_u_cla24_and3796_y0, h_u_cla24_and3795_y0, h_u_cla24_and3797_y0);
  and_gate and_gate_h_u_cla24_and3798_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and3798_y0);
  and_gate and_gate_h_u_cla24_and3799_y0(h_u_cla24_and3798_y0, h_u_cla24_and3797_y0, h_u_cla24_and3799_y0);
  and_gate and_gate_h_u_cla24_and3800_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and3800_y0);
  and_gate and_gate_h_u_cla24_and3801_y0(h_u_cla24_and3800_y0, h_u_cla24_and3799_y0, h_u_cla24_and3801_y0);
  and_gate and_gate_h_u_cla24_and3802_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and3802_y0);
  and_gate and_gate_h_u_cla24_and3803_y0(h_u_cla24_and3802_y0, h_u_cla24_and3801_y0, h_u_cla24_and3803_y0);
  and_gate and_gate_h_u_cla24_and3804_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and3804_y0);
  and_gate and_gate_h_u_cla24_and3805_y0(h_u_cla24_and3804_y0, h_u_cla24_and3803_y0, h_u_cla24_and3805_y0);
  and_gate and_gate_h_u_cla24_and3806_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and3806_y0);
  and_gate and_gate_h_u_cla24_and3807_y0(h_u_cla24_and3806_y0, h_u_cla24_and3805_y0, h_u_cla24_and3807_y0);
  and_gate and_gate_h_u_cla24_and3808_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and3808_y0);
  and_gate and_gate_h_u_cla24_and3809_y0(h_u_cla24_and3808_y0, h_u_cla24_and3807_y0, h_u_cla24_and3809_y0);
  and_gate and_gate_h_u_cla24_and3810_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and3810_y0);
  and_gate and_gate_h_u_cla24_and3811_y0(h_u_cla24_and3810_y0, h_u_cla24_and3809_y0, h_u_cla24_and3811_y0);
  and_gate and_gate_h_u_cla24_and3812_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and3812_y0);
  and_gate and_gate_h_u_cla24_and3813_y0(h_u_cla24_and3812_y0, h_u_cla24_and3811_y0, h_u_cla24_and3813_y0);
  and_gate and_gate_h_u_cla24_and3814_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and3814_y0);
  and_gate and_gate_h_u_cla24_and3815_y0(h_u_cla24_and3814_y0, h_u_cla24_and3813_y0, h_u_cla24_and3815_y0);
  and_gate and_gate_h_u_cla24_and3816_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and3816_y0);
  and_gate and_gate_h_u_cla24_and3817_y0(h_u_cla24_and3816_y0, h_u_cla24_and3815_y0, h_u_cla24_and3817_y0);
  and_gate and_gate_h_u_cla24_and3818_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and3818_y0);
  and_gate and_gate_h_u_cla24_and3819_y0(h_u_cla24_and3818_y0, h_u_cla24_and3817_y0, h_u_cla24_and3819_y0);
  and_gate and_gate_h_u_cla24_and3820_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and3820_y0);
  and_gate and_gate_h_u_cla24_and3821_y0(h_u_cla24_and3820_y0, h_u_cla24_and3819_y0, h_u_cla24_and3821_y0);
  and_gate and_gate_h_u_cla24_and3822_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and3822_y0);
  and_gate and_gate_h_u_cla24_and3823_y0(h_u_cla24_and3822_y0, h_u_cla24_and3821_y0, h_u_cla24_and3823_y0);
  and_gate and_gate_h_u_cla24_and3824_y0(h_u_cla24_pg_logic15_y0, constant_wire_0, h_u_cla24_and3824_y0);
  and_gate and_gate_h_u_cla24_and3825_y0(h_u_cla24_and3824_y0, h_u_cla24_and3823_y0, h_u_cla24_and3825_y0);
  and_gate and_gate_h_u_cla24_and3826_y0(h_u_cla24_pg_logic16_y0, constant_wire_0, h_u_cla24_and3826_y0);
  and_gate and_gate_h_u_cla24_and3827_y0(h_u_cla24_and3826_y0, h_u_cla24_and3825_y0, h_u_cla24_and3827_y0);
  and_gate and_gate_h_u_cla24_and3828_y0(h_u_cla24_pg_logic17_y0, constant_wire_0, h_u_cla24_and3828_y0);
  and_gate and_gate_h_u_cla24_and3829_y0(h_u_cla24_and3828_y0, h_u_cla24_and3827_y0, h_u_cla24_and3829_y0);
  and_gate and_gate_h_u_cla24_and3830_y0(h_u_cla24_pg_logic18_y0, constant_wire_0, h_u_cla24_and3830_y0);
  and_gate and_gate_h_u_cla24_and3831_y0(h_u_cla24_and3830_y0, h_u_cla24_and3829_y0, h_u_cla24_and3831_y0);
  and_gate and_gate_h_u_cla24_and3832_y0(h_u_cla24_pg_logic19_y0, constant_wire_0, h_u_cla24_and3832_y0);
  and_gate and_gate_h_u_cla24_and3833_y0(h_u_cla24_and3832_y0, h_u_cla24_and3831_y0, h_u_cla24_and3833_y0);
  and_gate and_gate_h_u_cla24_and3834_y0(h_u_cla24_pg_logic20_y0, constant_wire_0, h_u_cla24_and3834_y0);
  and_gate and_gate_h_u_cla24_and3835_y0(h_u_cla24_and3834_y0, h_u_cla24_and3833_y0, h_u_cla24_and3835_y0);
  and_gate and_gate_h_u_cla24_and3836_y0(h_u_cla24_pg_logic21_y0, constant_wire_0, h_u_cla24_and3836_y0);
  and_gate and_gate_h_u_cla24_and3837_y0(h_u_cla24_and3836_y0, h_u_cla24_and3835_y0, h_u_cla24_and3837_y0);
  and_gate and_gate_h_u_cla24_and3838_y0(h_u_cla24_pg_logic22_y0, constant_wire_0, h_u_cla24_and3838_y0);
  and_gate and_gate_h_u_cla24_and3839_y0(h_u_cla24_and3838_y0, h_u_cla24_and3837_y0, h_u_cla24_and3839_y0);
  and_gate and_gate_h_u_cla24_and3840_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3840_y0);
  and_gate and_gate_h_u_cla24_and3841_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3841_y0);
  and_gate and_gate_h_u_cla24_and3842_y0(h_u_cla24_and3841_y0, h_u_cla24_and3840_y0, h_u_cla24_and3842_y0);
  and_gate and_gate_h_u_cla24_and3843_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3843_y0);
  and_gate and_gate_h_u_cla24_and3844_y0(h_u_cla24_and3843_y0, h_u_cla24_and3842_y0, h_u_cla24_and3844_y0);
  and_gate and_gate_h_u_cla24_and3845_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3845_y0);
  and_gate and_gate_h_u_cla24_and3846_y0(h_u_cla24_and3845_y0, h_u_cla24_and3844_y0, h_u_cla24_and3846_y0);
  and_gate and_gate_h_u_cla24_and3847_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3847_y0);
  and_gate and_gate_h_u_cla24_and3848_y0(h_u_cla24_and3847_y0, h_u_cla24_and3846_y0, h_u_cla24_and3848_y0);
  and_gate and_gate_h_u_cla24_and3849_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3849_y0);
  and_gate and_gate_h_u_cla24_and3850_y0(h_u_cla24_and3849_y0, h_u_cla24_and3848_y0, h_u_cla24_and3850_y0);
  and_gate and_gate_h_u_cla24_and3851_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3851_y0);
  and_gate and_gate_h_u_cla24_and3852_y0(h_u_cla24_and3851_y0, h_u_cla24_and3850_y0, h_u_cla24_and3852_y0);
  and_gate and_gate_h_u_cla24_and3853_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3853_y0);
  and_gate and_gate_h_u_cla24_and3854_y0(h_u_cla24_and3853_y0, h_u_cla24_and3852_y0, h_u_cla24_and3854_y0);
  and_gate and_gate_h_u_cla24_and3855_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3855_y0);
  and_gate and_gate_h_u_cla24_and3856_y0(h_u_cla24_and3855_y0, h_u_cla24_and3854_y0, h_u_cla24_and3856_y0);
  and_gate and_gate_h_u_cla24_and3857_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3857_y0);
  and_gate and_gate_h_u_cla24_and3858_y0(h_u_cla24_and3857_y0, h_u_cla24_and3856_y0, h_u_cla24_and3858_y0);
  and_gate and_gate_h_u_cla24_and3859_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3859_y0);
  and_gate and_gate_h_u_cla24_and3860_y0(h_u_cla24_and3859_y0, h_u_cla24_and3858_y0, h_u_cla24_and3860_y0);
  and_gate and_gate_h_u_cla24_and3861_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3861_y0);
  and_gate and_gate_h_u_cla24_and3862_y0(h_u_cla24_and3861_y0, h_u_cla24_and3860_y0, h_u_cla24_and3862_y0);
  and_gate and_gate_h_u_cla24_and3863_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3863_y0);
  and_gate and_gate_h_u_cla24_and3864_y0(h_u_cla24_and3863_y0, h_u_cla24_and3862_y0, h_u_cla24_and3864_y0);
  and_gate and_gate_h_u_cla24_and3865_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3865_y0);
  and_gate and_gate_h_u_cla24_and3866_y0(h_u_cla24_and3865_y0, h_u_cla24_and3864_y0, h_u_cla24_and3866_y0);
  and_gate and_gate_h_u_cla24_and3867_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3867_y0);
  and_gate and_gate_h_u_cla24_and3868_y0(h_u_cla24_and3867_y0, h_u_cla24_and3866_y0, h_u_cla24_and3868_y0);
  and_gate and_gate_h_u_cla24_and3869_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3869_y0);
  and_gate and_gate_h_u_cla24_and3870_y0(h_u_cla24_and3869_y0, h_u_cla24_and3868_y0, h_u_cla24_and3870_y0);
  and_gate and_gate_h_u_cla24_and3871_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3871_y0);
  and_gate and_gate_h_u_cla24_and3872_y0(h_u_cla24_and3871_y0, h_u_cla24_and3870_y0, h_u_cla24_and3872_y0);
  and_gate and_gate_h_u_cla24_and3873_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3873_y0);
  and_gate and_gate_h_u_cla24_and3874_y0(h_u_cla24_and3873_y0, h_u_cla24_and3872_y0, h_u_cla24_and3874_y0);
  and_gate and_gate_h_u_cla24_and3875_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3875_y0);
  and_gate and_gate_h_u_cla24_and3876_y0(h_u_cla24_and3875_y0, h_u_cla24_and3874_y0, h_u_cla24_and3876_y0);
  and_gate and_gate_h_u_cla24_and3877_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3877_y0);
  and_gate and_gate_h_u_cla24_and3878_y0(h_u_cla24_and3877_y0, h_u_cla24_and3876_y0, h_u_cla24_and3878_y0);
  and_gate and_gate_h_u_cla24_and3879_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3879_y0);
  and_gate and_gate_h_u_cla24_and3880_y0(h_u_cla24_and3879_y0, h_u_cla24_and3878_y0, h_u_cla24_and3880_y0);
  and_gate and_gate_h_u_cla24_and3881_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and3881_y0);
  and_gate and_gate_h_u_cla24_and3882_y0(h_u_cla24_and3881_y0, h_u_cla24_and3880_y0, h_u_cla24_and3882_y0);
  and_gate and_gate_h_u_cla24_and3883_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3883_y0);
  and_gate and_gate_h_u_cla24_and3884_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3884_y0);
  and_gate and_gate_h_u_cla24_and3885_y0(h_u_cla24_and3884_y0, h_u_cla24_and3883_y0, h_u_cla24_and3885_y0);
  and_gate and_gate_h_u_cla24_and3886_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3886_y0);
  and_gate and_gate_h_u_cla24_and3887_y0(h_u_cla24_and3886_y0, h_u_cla24_and3885_y0, h_u_cla24_and3887_y0);
  and_gate and_gate_h_u_cla24_and3888_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3888_y0);
  and_gate and_gate_h_u_cla24_and3889_y0(h_u_cla24_and3888_y0, h_u_cla24_and3887_y0, h_u_cla24_and3889_y0);
  and_gate and_gate_h_u_cla24_and3890_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3890_y0);
  and_gate and_gate_h_u_cla24_and3891_y0(h_u_cla24_and3890_y0, h_u_cla24_and3889_y0, h_u_cla24_and3891_y0);
  and_gate and_gate_h_u_cla24_and3892_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3892_y0);
  and_gate and_gate_h_u_cla24_and3893_y0(h_u_cla24_and3892_y0, h_u_cla24_and3891_y0, h_u_cla24_and3893_y0);
  and_gate and_gate_h_u_cla24_and3894_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3894_y0);
  and_gate and_gate_h_u_cla24_and3895_y0(h_u_cla24_and3894_y0, h_u_cla24_and3893_y0, h_u_cla24_and3895_y0);
  and_gate and_gate_h_u_cla24_and3896_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3896_y0);
  and_gate and_gate_h_u_cla24_and3897_y0(h_u_cla24_and3896_y0, h_u_cla24_and3895_y0, h_u_cla24_and3897_y0);
  and_gate and_gate_h_u_cla24_and3898_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3898_y0);
  and_gate and_gate_h_u_cla24_and3899_y0(h_u_cla24_and3898_y0, h_u_cla24_and3897_y0, h_u_cla24_and3899_y0);
  and_gate and_gate_h_u_cla24_and3900_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3900_y0);
  and_gate and_gate_h_u_cla24_and3901_y0(h_u_cla24_and3900_y0, h_u_cla24_and3899_y0, h_u_cla24_and3901_y0);
  and_gate and_gate_h_u_cla24_and3902_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3902_y0);
  and_gate and_gate_h_u_cla24_and3903_y0(h_u_cla24_and3902_y0, h_u_cla24_and3901_y0, h_u_cla24_and3903_y0);
  and_gate and_gate_h_u_cla24_and3904_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3904_y0);
  and_gate and_gate_h_u_cla24_and3905_y0(h_u_cla24_and3904_y0, h_u_cla24_and3903_y0, h_u_cla24_and3905_y0);
  and_gate and_gate_h_u_cla24_and3906_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3906_y0);
  and_gate and_gate_h_u_cla24_and3907_y0(h_u_cla24_and3906_y0, h_u_cla24_and3905_y0, h_u_cla24_and3907_y0);
  and_gate and_gate_h_u_cla24_and3908_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3908_y0);
  and_gate and_gate_h_u_cla24_and3909_y0(h_u_cla24_and3908_y0, h_u_cla24_and3907_y0, h_u_cla24_and3909_y0);
  and_gate and_gate_h_u_cla24_and3910_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3910_y0);
  and_gate and_gate_h_u_cla24_and3911_y0(h_u_cla24_and3910_y0, h_u_cla24_and3909_y0, h_u_cla24_and3911_y0);
  and_gate and_gate_h_u_cla24_and3912_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3912_y0);
  and_gate and_gate_h_u_cla24_and3913_y0(h_u_cla24_and3912_y0, h_u_cla24_and3911_y0, h_u_cla24_and3913_y0);
  and_gate and_gate_h_u_cla24_and3914_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3914_y0);
  and_gate and_gate_h_u_cla24_and3915_y0(h_u_cla24_and3914_y0, h_u_cla24_and3913_y0, h_u_cla24_and3915_y0);
  and_gate and_gate_h_u_cla24_and3916_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3916_y0);
  and_gate and_gate_h_u_cla24_and3917_y0(h_u_cla24_and3916_y0, h_u_cla24_and3915_y0, h_u_cla24_and3917_y0);
  and_gate and_gate_h_u_cla24_and3918_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3918_y0);
  and_gate and_gate_h_u_cla24_and3919_y0(h_u_cla24_and3918_y0, h_u_cla24_and3917_y0, h_u_cla24_and3919_y0);
  and_gate and_gate_h_u_cla24_and3920_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3920_y0);
  and_gate and_gate_h_u_cla24_and3921_y0(h_u_cla24_and3920_y0, h_u_cla24_and3919_y0, h_u_cla24_and3921_y0);
  and_gate and_gate_h_u_cla24_and3922_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and3922_y0);
  and_gate and_gate_h_u_cla24_and3923_y0(h_u_cla24_and3922_y0, h_u_cla24_and3921_y0, h_u_cla24_and3923_y0);
  and_gate and_gate_h_u_cla24_and3924_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3924_y0);
  and_gate and_gate_h_u_cla24_and3925_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3925_y0);
  and_gate and_gate_h_u_cla24_and3926_y0(h_u_cla24_and3925_y0, h_u_cla24_and3924_y0, h_u_cla24_and3926_y0);
  and_gate and_gate_h_u_cla24_and3927_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3927_y0);
  and_gate and_gate_h_u_cla24_and3928_y0(h_u_cla24_and3927_y0, h_u_cla24_and3926_y0, h_u_cla24_and3928_y0);
  and_gate and_gate_h_u_cla24_and3929_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3929_y0);
  and_gate and_gate_h_u_cla24_and3930_y0(h_u_cla24_and3929_y0, h_u_cla24_and3928_y0, h_u_cla24_and3930_y0);
  and_gate and_gate_h_u_cla24_and3931_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3931_y0);
  and_gate and_gate_h_u_cla24_and3932_y0(h_u_cla24_and3931_y0, h_u_cla24_and3930_y0, h_u_cla24_and3932_y0);
  and_gate and_gate_h_u_cla24_and3933_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3933_y0);
  and_gate and_gate_h_u_cla24_and3934_y0(h_u_cla24_and3933_y0, h_u_cla24_and3932_y0, h_u_cla24_and3934_y0);
  and_gate and_gate_h_u_cla24_and3935_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3935_y0);
  and_gate and_gate_h_u_cla24_and3936_y0(h_u_cla24_and3935_y0, h_u_cla24_and3934_y0, h_u_cla24_and3936_y0);
  and_gate and_gate_h_u_cla24_and3937_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3937_y0);
  and_gate and_gate_h_u_cla24_and3938_y0(h_u_cla24_and3937_y0, h_u_cla24_and3936_y0, h_u_cla24_and3938_y0);
  and_gate and_gate_h_u_cla24_and3939_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3939_y0);
  and_gate and_gate_h_u_cla24_and3940_y0(h_u_cla24_and3939_y0, h_u_cla24_and3938_y0, h_u_cla24_and3940_y0);
  and_gate and_gate_h_u_cla24_and3941_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3941_y0);
  and_gate and_gate_h_u_cla24_and3942_y0(h_u_cla24_and3941_y0, h_u_cla24_and3940_y0, h_u_cla24_and3942_y0);
  and_gate and_gate_h_u_cla24_and3943_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3943_y0);
  and_gate and_gate_h_u_cla24_and3944_y0(h_u_cla24_and3943_y0, h_u_cla24_and3942_y0, h_u_cla24_and3944_y0);
  and_gate and_gate_h_u_cla24_and3945_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3945_y0);
  and_gate and_gate_h_u_cla24_and3946_y0(h_u_cla24_and3945_y0, h_u_cla24_and3944_y0, h_u_cla24_and3946_y0);
  and_gate and_gate_h_u_cla24_and3947_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3947_y0);
  and_gate and_gate_h_u_cla24_and3948_y0(h_u_cla24_and3947_y0, h_u_cla24_and3946_y0, h_u_cla24_and3948_y0);
  and_gate and_gate_h_u_cla24_and3949_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3949_y0);
  and_gate and_gate_h_u_cla24_and3950_y0(h_u_cla24_and3949_y0, h_u_cla24_and3948_y0, h_u_cla24_and3950_y0);
  and_gate and_gate_h_u_cla24_and3951_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3951_y0);
  and_gate and_gate_h_u_cla24_and3952_y0(h_u_cla24_and3951_y0, h_u_cla24_and3950_y0, h_u_cla24_and3952_y0);
  and_gate and_gate_h_u_cla24_and3953_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3953_y0);
  and_gate and_gate_h_u_cla24_and3954_y0(h_u_cla24_and3953_y0, h_u_cla24_and3952_y0, h_u_cla24_and3954_y0);
  and_gate and_gate_h_u_cla24_and3955_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3955_y0);
  and_gate and_gate_h_u_cla24_and3956_y0(h_u_cla24_and3955_y0, h_u_cla24_and3954_y0, h_u_cla24_and3956_y0);
  and_gate and_gate_h_u_cla24_and3957_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3957_y0);
  and_gate and_gate_h_u_cla24_and3958_y0(h_u_cla24_and3957_y0, h_u_cla24_and3956_y0, h_u_cla24_and3958_y0);
  and_gate and_gate_h_u_cla24_and3959_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3959_y0);
  and_gate and_gate_h_u_cla24_and3960_y0(h_u_cla24_and3959_y0, h_u_cla24_and3958_y0, h_u_cla24_and3960_y0);
  and_gate and_gate_h_u_cla24_and3961_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and3961_y0);
  and_gate and_gate_h_u_cla24_and3962_y0(h_u_cla24_and3961_y0, h_u_cla24_and3960_y0, h_u_cla24_and3962_y0);
  and_gate and_gate_h_u_cla24_and3963_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3963_y0);
  and_gate and_gate_h_u_cla24_and3964_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3964_y0);
  and_gate and_gate_h_u_cla24_and3965_y0(h_u_cla24_and3964_y0, h_u_cla24_and3963_y0, h_u_cla24_and3965_y0);
  and_gate and_gate_h_u_cla24_and3966_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3966_y0);
  and_gate and_gate_h_u_cla24_and3967_y0(h_u_cla24_and3966_y0, h_u_cla24_and3965_y0, h_u_cla24_and3967_y0);
  and_gate and_gate_h_u_cla24_and3968_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3968_y0);
  and_gate and_gate_h_u_cla24_and3969_y0(h_u_cla24_and3968_y0, h_u_cla24_and3967_y0, h_u_cla24_and3969_y0);
  and_gate and_gate_h_u_cla24_and3970_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3970_y0);
  and_gate and_gate_h_u_cla24_and3971_y0(h_u_cla24_and3970_y0, h_u_cla24_and3969_y0, h_u_cla24_and3971_y0);
  and_gate and_gate_h_u_cla24_and3972_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3972_y0);
  and_gate and_gate_h_u_cla24_and3973_y0(h_u_cla24_and3972_y0, h_u_cla24_and3971_y0, h_u_cla24_and3973_y0);
  and_gate and_gate_h_u_cla24_and3974_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3974_y0);
  and_gate and_gate_h_u_cla24_and3975_y0(h_u_cla24_and3974_y0, h_u_cla24_and3973_y0, h_u_cla24_and3975_y0);
  and_gate and_gate_h_u_cla24_and3976_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3976_y0);
  and_gate and_gate_h_u_cla24_and3977_y0(h_u_cla24_and3976_y0, h_u_cla24_and3975_y0, h_u_cla24_and3977_y0);
  and_gate and_gate_h_u_cla24_and3978_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3978_y0);
  and_gate and_gate_h_u_cla24_and3979_y0(h_u_cla24_and3978_y0, h_u_cla24_and3977_y0, h_u_cla24_and3979_y0);
  and_gate and_gate_h_u_cla24_and3980_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3980_y0);
  and_gate and_gate_h_u_cla24_and3981_y0(h_u_cla24_and3980_y0, h_u_cla24_and3979_y0, h_u_cla24_and3981_y0);
  and_gate and_gate_h_u_cla24_and3982_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3982_y0);
  and_gate and_gate_h_u_cla24_and3983_y0(h_u_cla24_and3982_y0, h_u_cla24_and3981_y0, h_u_cla24_and3983_y0);
  and_gate and_gate_h_u_cla24_and3984_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3984_y0);
  and_gate and_gate_h_u_cla24_and3985_y0(h_u_cla24_and3984_y0, h_u_cla24_and3983_y0, h_u_cla24_and3985_y0);
  and_gate and_gate_h_u_cla24_and3986_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3986_y0);
  and_gate and_gate_h_u_cla24_and3987_y0(h_u_cla24_and3986_y0, h_u_cla24_and3985_y0, h_u_cla24_and3987_y0);
  and_gate and_gate_h_u_cla24_and3988_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3988_y0);
  and_gate and_gate_h_u_cla24_and3989_y0(h_u_cla24_and3988_y0, h_u_cla24_and3987_y0, h_u_cla24_and3989_y0);
  and_gate and_gate_h_u_cla24_and3990_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3990_y0);
  and_gate and_gate_h_u_cla24_and3991_y0(h_u_cla24_and3990_y0, h_u_cla24_and3989_y0, h_u_cla24_and3991_y0);
  and_gate and_gate_h_u_cla24_and3992_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3992_y0);
  and_gate and_gate_h_u_cla24_and3993_y0(h_u_cla24_and3992_y0, h_u_cla24_and3991_y0, h_u_cla24_and3993_y0);
  and_gate and_gate_h_u_cla24_and3994_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3994_y0);
  and_gate and_gate_h_u_cla24_and3995_y0(h_u_cla24_and3994_y0, h_u_cla24_and3993_y0, h_u_cla24_and3995_y0);
  and_gate and_gate_h_u_cla24_and3996_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3996_y0);
  and_gate and_gate_h_u_cla24_and3997_y0(h_u_cla24_and3996_y0, h_u_cla24_and3995_y0, h_u_cla24_and3997_y0);
  and_gate and_gate_h_u_cla24_and3998_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and3998_y0);
  and_gate and_gate_h_u_cla24_and3999_y0(h_u_cla24_and3998_y0, h_u_cla24_and3997_y0, h_u_cla24_and3999_y0);
  and_gate and_gate_h_u_cla24_and4000_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4000_y0);
  and_gate and_gate_h_u_cla24_and4001_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4001_y0);
  and_gate and_gate_h_u_cla24_and4002_y0(h_u_cla24_and4001_y0, h_u_cla24_and4000_y0, h_u_cla24_and4002_y0);
  and_gate and_gate_h_u_cla24_and4003_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4003_y0);
  and_gate and_gate_h_u_cla24_and4004_y0(h_u_cla24_and4003_y0, h_u_cla24_and4002_y0, h_u_cla24_and4004_y0);
  and_gate and_gate_h_u_cla24_and4005_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4005_y0);
  and_gate and_gate_h_u_cla24_and4006_y0(h_u_cla24_and4005_y0, h_u_cla24_and4004_y0, h_u_cla24_and4006_y0);
  and_gate and_gate_h_u_cla24_and4007_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4007_y0);
  and_gate and_gate_h_u_cla24_and4008_y0(h_u_cla24_and4007_y0, h_u_cla24_and4006_y0, h_u_cla24_and4008_y0);
  and_gate and_gate_h_u_cla24_and4009_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4009_y0);
  and_gate and_gate_h_u_cla24_and4010_y0(h_u_cla24_and4009_y0, h_u_cla24_and4008_y0, h_u_cla24_and4010_y0);
  and_gate and_gate_h_u_cla24_and4011_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4011_y0);
  and_gate and_gate_h_u_cla24_and4012_y0(h_u_cla24_and4011_y0, h_u_cla24_and4010_y0, h_u_cla24_and4012_y0);
  and_gate and_gate_h_u_cla24_and4013_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4013_y0);
  and_gate and_gate_h_u_cla24_and4014_y0(h_u_cla24_and4013_y0, h_u_cla24_and4012_y0, h_u_cla24_and4014_y0);
  and_gate and_gate_h_u_cla24_and4015_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4015_y0);
  and_gate and_gate_h_u_cla24_and4016_y0(h_u_cla24_and4015_y0, h_u_cla24_and4014_y0, h_u_cla24_and4016_y0);
  and_gate and_gate_h_u_cla24_and4017_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4017_y0);
  and_gate and_gate_h_u_cla24_and4018_y0(h_u_cla24_and4017_y0, h_u_cla24_and4016_y0, h_u_cla24_and4018_y0);
  and_gate and_gate_h_u_cla24_and4019_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4019_y0);
  and_gate and_gate_h_u_cla24_and4020_y0(h_u_cla24_and4019_y0, h_u_cla24_and4018_y0, h_u_cla24_and4020_y0);
  and_gate and_gate_h_u_cla24_and4021_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4021_y0);
  and_gate and_gate_h_u_cla24_and4022_y0(h_u_cla24_and4021_y0, h_u_cla24_and4020_y0, h_u_cla24_and4022_y0);
  and_gate and_gate_h_u_cla24_and4023_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4023_y0);
  and_gate and_gate_h_u_cla24_and4024_y0(h_u_cla24_and4023_y0, h_u_cla24_and4022_y0, h_u_cla24_and4024_y0);
  and_gate and_gate_h_u_cla24_and4025_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4025_y0);
  and_gate and_gate_h_u_cla24_and4026_y0(h_u_cla24_and4025_y0, h_u_cla24_and4024_y0, h_u_cla24_and4026_y0);
  and_gate and_gate_h_u_cla24_and4027_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4027_y0);
  and_gate and_gate_h_u_cla24_and4028_y0(h_u_cla24_and4027_y0, h_u_cla24_and4026_y0, h_u_cla24_and4028_y0);
  and_gate and_gate_h_u_cla24_and4029_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4029_y0);
  and_gate and_gate_h_u_cla24_and4030_y0(h_u_cla24_and4029_y0, h_u_cla24_and4028_y0, h_u_cla24_and4030_y0);
  and_gate and_gate_h_u_cla24_and4031_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4031_y0);
  and_gate and_gate_h_u_cla24_and4032_y0(h_u_cla24_and4031_y0, h_u_cla24_and4030_y0, h_u_cla24_and4032_y0);
  and_gate and_gate_h_u_cla24_and4033_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4033_y0);
  and_gate and_gate_h_u_cla24_and4034_y0(h_u_cla24_and4033_y0, h_u_cla24_and4032_y0, h_u_cla24_and4034_y0);
  and_gate and_gate_h_u_cla24_and4035_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4035_y0);
  and_gate and_gate_h_u_cla24_and4036_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4036_y0);
  and_gate and_gate_h_u_cla24_and4037_y0(h_u_cla24_and4036_y0, h_u_cla24_and4035_y0, h_u_cla24_and4037_y0);
  and_gate and_gate_h_u_cla24_and4038_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4038_y0);
  and_gate and_gate_h_u_cla24_and4039_y0(h_u_cla24_and4038_y0, h_u_cla24_and4037_y0, h_u_cla24_and4039_y0);
  and_gate and_gate_h_u_cla24_and4040_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4040_y0);
  and_gate and_gate_h_u_cla24_and4041_y0(h_u_cla24_and4040_y0, h_u_cla24_and4039_y0, h_u_cla24_and4041_y0);
  and_gate and_gate_h_u_cla24_and4042_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4042_y0);
  and_gate and_gate_h_u_cla24_and4043_y0(h_u_cla24_and4042_y0, h_u_cla24_and4041_y0, h_u_cla24_and4043_y0);
  and_gate and_gate_h_u_cla24_and4044_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4044_y0);
  and_gate and_gate_h_u_cla24_and4045_y0(h_u_cla24_and4044_y0, h_u_cla24_and4043_y0, h_u_cla24_and4045_y0);
  and_gate and_gate_h_u_cla24_and4046_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4046_y0);
  and_gate and_gate_h_u_cla24_and4047_y0(h_u_cla24_and4046_y0, h_u_cla24_and4045_y0, h_u_cla24_and4047_y0);
  and_gate and_gate_h_u_cla24_and4048_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4048_y0);
  and_gate and_gate_h_u_cla24_and4049_y0(h_u_cla24_and4048_y0, h_u_cla24_and4047_y0, h_u_cla24_and4049_y0);
  and_gate and_gate_h_u_cla24_and4050_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4050_y0);
  and_gate and_gate_h_u_cla24_and4051_y0(h_u_cla24_and4050_y0, h_u_cla24_and4049_y0, h_u_cla24_and4051_y0);
  and_gate and_gate_h_u_cla24_and4052_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4052_y0);
  and_gate and_gate_h_u_cla24_and4053_y0(h_u_cla24_and4052_y0, h_u_cla24_and4051_y0, h_u_cla24_and4053_y0);
  and_gate and_gate_h_u_cla24_and4054_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4054_y0);
  and_gate and_gate_h_u_cla24_and4055_y0(h_u_cla24_and4054_y0, h_u_cla24_and4053_y0, h_u_cla24_and4055_y0);
  and_gate and_gate_h_u_cla24_and4056_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4056_y0);
  and_gate and_gate_h_u_cla24_and4057_y0(h_u_cla24_and4056_y0, h_u_cla24_and4055_y0, h_u_cla24_and4057_y0);
  and_gate and_gate_h_u_cla24_and4058_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4058_y0);
  and_gate and_gate_h_u_cla24_and4059_y0(h_u_cla24_and4058_y0, h_u_cla24_and4057_y0, h_u_cla24_and4059_y0);
  and_gate and_gate_h_u_cla24_and4060_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4060_y0);
  and_gate and_gate_h_u_cla24_and4061_y0(h_u_cla24_and4060_y0, h_u_cla24_and4059_y0, h_u_cla24_and4061_y0);
  and_gate and_gate_h_u_cla24_and4062_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4062_y0);
  and_gate and_gate_h_u_cla24_and4063_y0(h_u_cla24_and4062_y0, h_u_cla24_and4061_y0, h_u_cla24_and4063_y0);
  and_gate and_gate_h_u_cla24_and4064_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4064_y0);
  and_gate and_gate_h_u_cla24_and4065_y0(h_u_cla24_and4064_y0, h_u_cla24_and4063_y0, h_u_cla24_and4065_y0);
  and_gate and_gate_h_u_cla24_and4066_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4066_y0);
  and_gate and_gate_h_u_cla24_and4067_y0(h_u_cla24_and4066_y0, h_u_cla24_and4065_y0, h_u_cla24_and4067_y0);
  and_gate and_gate_h_u_cla24_and4068_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4068_y0);
  and_gate and_gate_h_u_cla24_and4069_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4069_y0);
  and_gate and_gate_h_u_cla24_and4070_y0(h_u_cla24_and4069_y0, h_u_cla24_and4068_y0, h_u_cla24_and4070_y0);
  and_gate and_gate_h_u_cla24_and4071_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4071_y0);
  and_gate and_gate_h_u_cla24_and4072_y0(h_u_cla24_and4071_y0, h_u_cla24_and4070_y0, h_u_cla24_and4072_y0);
  and_gate and_gate_h_u_cla24_and4073_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4073_y0);
  and_gate and_gate_h_u_cla24_and4074_y0(h_u_cla24_and4073_y0, h_u_cla24_and4072_y0, h_u_cla24_and4074_y0);
  and_gate and_gate_h_u_cla24_and4075_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4075_y0);
  and_gate and_gate_h_u_cla24_and4076_y0(h_u_cla24_and4075_y0, h_u_cla24_and4074_y0, h_u_cla24_and4076_y0);
  and_gate and_gate_h_u_cla24_and4077_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4077_y0);
  and_gate and_gate_h_u_cla24_and4078_y0(h_u_cla24_and4077_y0, h_u_cla24_and4076_y0, h_u_cla24_and4078_y0);
  and_gate and_gate_h_u_cla24_and4079_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4079_y0);
  and_gate and_gate_h_u_cla24_and4080_y0(h_u_cla24_and4079_y0, h_u_cla24_and4078_y0, h_u_cla24_and4080_y0);
  and_gate and_gate_h_u_cla24_and4081_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4081_y0);
  and_gate and_gate_h_u_cla24_and4082_y0(h_u_cla24_and4081_y0, h_u_cla24_and4080_y0, h_u_cla24_and4082_y0);
  and_gate and_gate_h_u_cla24_and4083_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4083_y0);
  and_gate and_gate_h_u_cla24_and4084_y0(h_u_cla24_and4083_y0, h_u_cla24_and4082_y0, h_u_cla24_and4084_y0);
  and_gate and_gate_h_u_cla24_and4085_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4085_y0);
  and_gate and_gate_h_u_cla24_and4086_y0(h_u_cla24_and4085_y0, h_u_cla24_and4084_y0, h_u_cla24_and4086_y0);
  and_gate and_gate_h_u_cla24_and4087_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4087_y0);
  and_gate and_gate_h_u_cla24_and4088_y0(h_u_cla24_and4087_y0, h_u_cla24_and4086_y0, h_u_cla24_and4088_y0);
  and_gate and_gate_h_u_cla24_and4089_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4089_y0);
  and_gate and_gate_h_u_cla24_and4090_y0(h_u_cla24_and4089_y0, h_u_cla24_and4088_y0, h_u_cla24_and4090_y0);
  and_gate and_gate_h_u_cla24_and4091_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4091_y0);
  and_gate and_gate_h_u_cla24_and4092_y0(h_u_cla24_and4091_y0, h_u_cla24_and4090_y0, h_u_cla24_and4092_y0);
  and_gate and_gate_h_u_cla24_and4093_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4093_y0);
  and_gate and_gate_h_u_cla24_and4094_y0(h_u_cla24_and4093_y0, h_u_cla24_and4092_y0, h_u_cla24_and4094_y0);
  and_gate and_gate_h_u_cla24_and4095_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4095_y0);
  and_gate and_gate_h_u_cla24_and4096_y0(h_u_cla24_and4095_y0, h_u_cla24_and4094_y0, h_u_cla24_and4096_y0);
  and_gate and_gate_h_u_cla24_and4097_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4097_y0);
  and_gate and_gate_h_u_cla24_and4098_y0(h_u_cla24_and4097_y0, h_u_cla24_and4096_y0, h_u_cla24_and4098_y0);
  and_gate and_gate_h_u_cla24_and4099_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4099_y0);
  and_gate and_gate_h_u_cla24_and4100_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4100_y0);
  and_gate and_gate_h_u_cla24_and4101_y0(h_u_cla24_and4100_y0, h_u_cla24_and4099_y0, h_u_cla24_and4101_y0);
  and_gate and_gate_h_u_cla24_and4102_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4102_y0);
  and_gate and_gate_h_u_cla24_and4103_y0(h_u_cla24_and4102_y0, h_u_cla24_and4101_y0, h_u_cla24_and4103_y0);
  and_gate and_gate_h_u_cla24_and4104_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4104_y0);
  and_gate and_gate_h_u_cla24_and4105_y0(h_u_cla24_and4104_y0, h_u_cla24_and4103_y0, h_u_cla24_and4105_y0);
  and_gate and_gate_h_u_cla24_and4106_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4106_y0);
  and_gate and_gate_h_u_cla24_and4107_y0(h_u_cla24_and4106_y0, h_u_cla24_and4105_y0, h_u_cla24_and4107_y0);
  and_gate and_gate_h_u_cla24_and4108_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4108_y0);
  and_gate and_gate_h_u_cla24_and4109_y0(h_u_cla24_and4108_y0, h_u_cla24_and4107_y0, h_u_cla24_and4109_y0);
  and_gate and_gate_h_u_cla24_and4110_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4110_y0);
  and_gate and_gate_h_u_cla24_and4111_y0(h_u_cla24_and4110_y0, h_u_cla24_and4109_y0, h_u_cla24_and4111_y0);
  and_gate and_gate_h_u_cla24_and4112_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4112_y0);
  and_gate and_gate_h_u_cla24_and4113_y0(h_u_cla24_and4112_y0, h_u_cla24_and4111_y0, h_u_cla24_and4113_y0);
  and_gate and_gate_h_u_cla24_and4114_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4114_y0);
  and_gate and_gate_h_u_cla24_and4115_y0(h_u_cla24_and4114_y0, h_u_cla24_and4113_y0, h_u_cla24_and4115_y0);
  and_gate and_gate_h_u_cla24_and4116_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4116_y0);
  and_gate and_gate_h_u_cla24_and4117_y0(h_u_cla24_and4116_y0, h_u_cla24_and4115_y0, h_u_cla24_and4117_y0);
  and_gate and_gate_h_u_cla24_and4118_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4118_y0);
  and_gate and_gate_h_u_cla24_and4119_y0(h_u_cla24_and4118_y0, h_u_cla24_and4117_y0, h_u_cla24_and4119_y0);
  and_gate and_gate_h_u_cla24_and4120_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4120_y0);
  and_gate and_gate_h_u_cla24_and4121_y0(h_u_cla24_and4120_y0, h_u_cla24_and4119_y0, h_u_cla24_and4121_y0);
  and_gate and_gate_h_u_cla24_and4122_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4122_y0);
  and_gate and_gate_h_u_cla24_and4123_y0(h_u_cla24_and4122_y0, h_u_cla24_and4121_y0, h_u_cla24_and4123_y0);
  and_gate and_gate_h_u_cla24_and4124_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4124_y0);
  and_gate and_gate_h_u_cla24_and4125_y0(h_u_cla24_and4124_y0, h_u_cla24_and4123_y0, h_u_cla24_and4125_y0);
  and_gate and_gate_h_u_cla24_and4126_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4126_y0);
  and_gate and_gate_h_u_cla24_and4127_y0(h_u_cla24_and4126_y0, h_u_cla24_and4125_y0, h_u_cla24_and4127_y0);
  and_gate and_gate_h_u_cla24_and4128_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4128_y0);
  and_gate and_gate_h_u_cla24_and4129_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4129_y0);
  and_gate and_gate_h_u_cla24_and4130_y0(h_u_cla24_and4129_y0, h_u_cla24_and4128_y0, h_u_cla24_and4130_y0);
  and_gate and_gate_h_u_cla24_and4131_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4131_y0);
  and_gate and_gate_h_u_cla24_and4132_y0(h_u_cla24_and4131_y0, h_u_cla24_and4130_y0, h_u_cla24_and4132_y0);
  and_gate and_gate_h_u_cla24_and4133_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4133_y0);
  and_gate and_gate_h_u_cla24_and4134_y0(h_u_cla24_and4133_y0, h_u_cla24_and4132_y0, h_u_cla24_and4134_y0);
  and_gate and_gate_h_u_cla24_and4135_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4135_y0);
  and_gate and_gate_h_u_cla24_and4136_y0(h_u_cla24_and4135_y0, h_u_cla24_and4134_y0, h_u_cla24_and4136_y0);
  and_gate and_gate_h_u_cla24_and4137_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4137_y0);
  and_gate and_gate_h_u_cla24_and4138_y0(h_u_cla24_and4137_y0, h_u_cla24_and4136_y0, h_u_cla24_and4138_y0);
  and_gate and_gate_h_u_cla24_and4139_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4139_y0);
  and_gate and_gate_h_u_cla24_and4140_y0(h_u_cla24_and4139_y0, h_u_cla24_and4138_y0, h_u_cla24_and4140_y0);
  and_gate and_gate_h_u_cla24_and4141_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4141_y0);
  and_gate and_gate_h_u_cla24_and4142_y0(h_u_cla24_and4141_y0, h_u_cla24_and4140_y0, h_u_cla24_and4142_y0);
  and_gate and_gate_h_u_cla24_and4143_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4143_y0);
  and_gate and_gate_h_u_cla24_and4144_y0(h_u_cla24_and4143_y0, h_u_cla24_and4142_y0, h_u_cla24_and4144_y0);
  and_gate and_gate_h_u_cla24_and4145_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4145_y0);
  and_gate and_gate_h_u_cla24_and4146_y0(h_u_cla24_and4145_y0, h_u_cla24_and4144_y0, h_u_cla24_and4146_y0);
  and_gate and_gate_h_u_cla24_and4147_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4147_y0);
  and_gate and_gate_h_u_cla24_and4148_y0(h_u_cla24_and4147_y0, h_u_cla24_and4146_y0, h_u_cla24_and4148_y0);
  and_gate and_gate_h_u_cla24_and4149_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4149_y0);
  and_gate and_gate_h_u_cla24_and4150_y0(h_u_cla24_and4149_y0, h_u_cla24_and4148_y0, h_u_cla24_and4150_y0);
  and_gate and_gate_h_u_cla24_and4151_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4151_y0);
  and_gate and_gate_h_u_cla24_and4152_y0(h_u_cla24_and4151_y0, h_u_cla24_and4150_y0, h_u_cla24_and4152_y0);
  and_gate and_gate_h_u_cla24_and4153_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4153_y0);
  and_gate and_gate_h_u_cla24_and4154_y0(h_u_cla24_and4153_y0, h_u_cla24_and4152_y0, h_u_cla24_and4154_y0);
  and_gate and_gate_h_u_cla24_and4155_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4155_y0);
  and_gate and_gate_h_u_cla24_and4156_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4156_y0);
  and_gate and_gate_h_u_cla24_and4157_y0(h_u_cla24_and4156_y0, h_u_cla24_and4155_y0, h_u_cla24_and4157_y0);
  and_gate and_gate_h_u_cla24_and4158_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4158_y0);
  and_gate and_gate_h_u_cla24_and4159_y0(h_u_cla24_and4158_y0, h_u_cla24_and4157_y0, h_u_cla24_and4159_y0);
  and_gate and_gate_h_u_cla24_and4160_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4160_y0);
  and_gate and_gate_h_u_cla24_and4161_y0(h_u_cla24_and4160_y0, h_u_cla24_and4159_y0, h_u_cla24_and4161_y0);
  and_gate and_gate_h_u_cla24_and4162_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4162_y0);
  and_gate and_gate_h_u_cla24_and4163_y0(h_u_cla24_and4162_y0, h_u_cla24_and4161_y0, h_u_cla24_and4163_y0);
  and_gate and_gate_h_u_cla24_and4164_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4164_y0);
  and_gate and_gate_h_u_cla24_and4165_y0(h_u_cla24_and4164_y0, h_u_cla24_and4163_y0, h_u_cla24_and4165_y0);
  and_gate and_gate_h_u_cla24_and4166_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4166_y0);
  and_gate and_gate_h_u_cla24_and4167_y0(h_u_cla24_and4166_y0, h_u_cla24_and4165_y0, h_u_cla24_and4167_y0);
  and_gate and_gate_h_u_cla24_and4168_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4168_y0);
  and_gate and_gate_h_u_cla24_and4169_y0(h_u_cla24_and4168_y0, h_u_cla24_and4167_y0, h_u_cla24_and4169_y0);
  and_gate and_gate_h_u_cla24_and4170_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4170_y0);
  and_gate and_gate_h_u_cla24_and4171_y0(h_u_cla24_and4170_y0, h_u_cla24_and4169_y0, h_u_cla24_and4171_y0);
  and_gate and_gate_h_u_cla24_and4172_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4172_y0);
  and_gate and_gate_h_u_cla24_and4173_y0(h_u_cla24_and4172_y0, h_u_cla24_and4171_y0, h_u_cla24_and4173_y0);
  and_gate and_gate_h_u_cla24_and4174_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4174_y0);
  and_gate and_gate_h_u_cla24_and4175_y0(h_u_cla24_and4174_y0, h_u_cla24_and4173_y0, h_u_cla24_and4175_y0);
  and_gate and_gate_h_u_cla24_and4176_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4176_y0);
  and_gate and_gate_h_u_cla24_and4177_y0(h_u_cla24_and4176_y0, h_u_cla24_and4175_y0, h_u_cla24_and4177_y0);
  and_gate and_gate_h_u_cla24_and4178_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4178_y0);
  and_gate and_gate_h_u_cla24_and4179_y0(h_u_cla24_and4178_y0, h_u_cla24_and4177_y0, h_u_cla24_and4179_y0);
  and_gate and_gate_h_u_cla24_and4180_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4180_y0);
  and_gate and_gate_h_u_cla24_and4181_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4181_y0);
  and_gate and_gate_h_u_cla24_and4182_y0(h_u_cla24_and4181_y0, h_u_cla24_and4180_y0, h_u_cla24_and4182_y0);
  and_gate and_gate_h_u_cla24_and4183_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4183_y0);
  and_gate and_gate_h_u_cla24_and4184_y0(h_u_cla24_and4183_y0, h_u_cla24_and4182_y0, h_u_cla24_and4184_y0);
  and_gate and_gate_h_u_cla24_and4185_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4185_y0);
  and_gate and_gate_h_u_cla24_and4186_y0(h_u_cla24_and4185_y0, h_u_cla24_and4184_y0, h_u_cla24_and4186_y0);
  and_gate and_gate_h_u_cla24_and4187_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4187_y0);
  and_gate and_gate_h_u_cla24_and4188_y0(h_u_cla24_and4187_y0, h_u_cla24_and4186_y0, h_u_cla24_and4188_y0);
  and_gate and_gate_h_u_cla24_and4189_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4189_y0);
  and_gate and_gate_h_u_cla24_and4190_y0(h_u_cla24_and4189_y0, h_u_cla24_and4188_y0, h_u_cla24_and4190_y0);
  and_gate and_gate_h_u_cla24_and4191_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4191_y0);
  and_gate and_gate_h_u_cla24_and4192_y0(h_u_cla24_and4191_y0, h_u_cla24_and4190_y0, h_u_cla24_and4192_y0);
  and_gate and_gate_h_u_cla24_and4193_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4193_y0);
  and_gate and_gate_h_u_cla24_and4194_y0(h_u_cla24_and4193_y0, h_u_cla24_and4192_y0, h_u_cla24_and4194_y0);
  and_gate and_gate_h_u_cla24_and4195_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4195_y0);
  and_gate and_gate_h_u_cla24_and4196_y0(h_u_cla24_and4195_y0, h_u_cla24_and4194_y0, h_u_cla24_and4196_y0);
  and_gate and_gate_h_u_cla24_and4197_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4197_y0);
  and_gate and_gate_h_u_cla24_and4198_y0(h_u_cla24_and4197_y0, h_u_cla24_and4196_y0, h_u_cla24_and4198_y0);
  and_gate and_gate_h_u_cla24_and4199_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4199_y0);
  and_gate and_gate_h_u_cla24_and4200_y0(h_u_cla24_and4199_y0, h_u_cla24_and4198_y0, h_u_cla24_and4200_y0);
  and_gate and_gate_h_u_cla24_and4201_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4201_y0);
  and_gate and_gate_h_u_cla24_and4202_y0(h_u_cla24_and4201_y0, h_u_cla24_and4200_y0, h_u_cla24_and4202_y0);
  and_gate and_gate_h_u_cla24_and4203_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4203_y0);
  and_gate and_gate_h_u_cla24_and4204_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4204_y0);
  and_gate and_gate_h_u_cla24_and4205_y0(h_u_cla24_and4204_y0, h_u_cla24_and4203_y0, h_u_cla24_and4205_y0);
  and_gate and_gate_h_u_cla24_and4206_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4206_y0);
  and_gate and_gate_h_u_cla24_and4207_y0(h_u_cla24_and4206_y0, h_u_cla24_and4205_y0, h_u_cla24_and4207_y0);
  and_gate and_gate_h_u_cla24_and4208_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4208_y0);
  and_gate and_gate_h_u_cla24_and4209_y0(h_u_cla24_and4208_y0, h_u_cla24_and4207_y0, h_u_cla24_and4209_y0);
  and_gate and_gate_h_u_cla24_and4210_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4210_y0);
  and_gate and_gate_h_u_cla24_and4211_y0(h_u_cla24_and4210_y0, h_u_cla24_and4209_y0, h_u_cla24_and4211_y0);
  and_gate and_gate_h_u_cla24_and4212_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4212_y0);
  and_gate and_gate_h_u_cla24_and4213_y0(h_u_cla24_and4212_y0, h_u_cla24_and4211_y0, h_u_cla24_and4213_y0);
  and_gate and_gate_h_u_cla24_and4214_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4214_y0);
  and_gate and_gate_h_u_cla24_and4215_y0(h_u_cla24_and4214_y0, h_u_cla24_and4213_y0, h_u_cla24_and4215_y0);
  and_gate and_gate_h_u_cla24_and4216_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4216_y0);
  and_gate and_gate_h_u_cla24_and4217_y0(h_u_cla24_and4216_y0, h_u_cla24_and4215_y0, h_u_cla24_and4217_y0);
  and_gate and_gate_h_u_cla24_and4218_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4218_y0);
  and_gate and_gate_h_u_cla24_and4219_y0(h_u_cla24_and4218_y0, h_u_cla24_and4217_y0, h_u_cla24_and4219_y0);
  and_gate and_gate_h_u_cla24_and4220_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4220_y0);
  and_gate and_gate_h_u_cla24_and4221_y0(h_u_cla24_and4220_y0, h_u_cla24_and4219_y0, h_u_cla24_and4221_y0);
  and_gate and_gate_h_u_cla24_and4222_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4222_y0);
  and_gate and_gate_h_u_cla24_and4223_y0(h_u_cla24_and4222_y0, h_u_cla24_and4221_y0, h_u_cla24_and4223_y0);
  and_gate and_gate_h_u_cla24_and4224_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4224_y0);
  and_gate and_gate_h_u_cla24_and4225_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4225_y0);
  and_gate and_gate_h_u_cla24_and4226_y0(h_u_cla24_and4225_y0, h_u_cla24_and4224_y0, h_u_cla24_and4226_y0);
  and_gate and_gate_h_u_cla24_and4227_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4227_y0);
  and_gate and_gate_h_u_cla24_and4228_y0(h_u_cla24_and4227_y0, h_u_cla24_and4226_y0, h_u_cla24_and4228_y0);
  and_gate and_gate_h_u_cla24_and4229_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4229_y0);
  and_gate and_gate_h_u_cla24_and4230_y0(h_u_cla24_and4229_y0, h_u_cla24_and4228_y0, h_u_cla24_and4230_y0);
  and_gate and_gate_h_u_cla24_and4231_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4231_y0);
  and_gate and_gate_h_u_cla24_and4232_y0(h_u_cla24_and4231_y0, h_u_cla24_and4230_y0, h_u_cla24_and4232_y0);
  and_gate and_gate_h_u_cla24_and4233_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4233_y0);
  and_gate and_gate_h_u_cla24_and4234_y0(h_u_cla24_and4233_y0, h_u_cla24_and4232_y0, h_u_cla24_and4234_y0);
  and_gate and_gate_h_u_cla24_and4235_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4235_y0);
  and_gate and_gate_h_u_cla24_and4236_y0(h_u_cla24_and4235_y0, h_u_cla24_and4234_y0, h_u_cla24_and4236_y0);
  and_gate and_gate_h_u_cla24_and4237_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4237_y0);
  and_gate and_gate_h_u_cla24_and4238_y0(h_u_cla24_and4237_y0, h_u_cla24_and4236_y0, h_u_cla24_and4238_y0);
  and_gate and_gate_h_u_cla24_and4239_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4239_y0);
  and_gate and_gate_h_u_cla24_and4240_y0(h_u_cla24_and4239_y0, h_u_cla24_and4238_y0, h_u_cla24_and4240_y0);
  and_gate and_gate_h_u_cla24_and4241_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4241_y0);
  and_gate and_gate_h_u_cla24_and4242_y0(h_u_cla24_and4241_y0, h_u_cla24_and4240_y0, h_u_cla24_and4242_y0);
  and_gate and_gate_h_u_cla24_and4243_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4243_y0);
  and_gate and_gate_h_u_cla24_and4244_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4244_y0);
  and_gate and_gate_h_u_cla24_and4245_y0(h_u_cla24_and4244_y0, h_u_cla24_and4243_y0, h_u_cla24_and4245_y0);
  and_gate and_gate_h_u_cla24_and4246_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4246_y0);
  and_gate and_gate_h_u_cla24_and4247_y0(h_u_cla24_and4246_y0, h_u_cla24_and4245_y0, h_u_cla24_and4247_y0);
  and_gate and_gate_h_u_cla24_and4248_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4248_y0);
  and_gate and_gate_h_u_cla24_and4249_y0(h_u_cla24_and4248_y0, h_u_cla24_and4247_y0, h_u_cla24_and4249_y0);
  and_gate and_gate_h_u_cla24_and4250_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4250_y0);
  and_gate and_gate_h_u_cla24_and4251_y0(h_u_cla24_and4250_y0, h_u_cla24_and4249_y0, h_u_cla24_and4251_y0);
  and_gate and_gate_h_u_cla24_and4252_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4252_y0);
  and_gate and_gate_h_u_cla24_and4253_y0(h_u_cla24_and4252_y0, h_u_cla24_and4251_y0, h_u_cla24_and4253_y0);
  and_gate and_gate_h_u_cla24_and4254_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4254_y0);
  and_gate and_gate_h_u_cla24_and4255_y0(h_u_cla24_and4254_y0, h_u_cla24_and4253_y0, h_u_cla24_and4255_y0);
  and_gate and_gate_h_u_cla24_and4256_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4256_y0);
  and_gate and_gate_h_u_cla24_and4257_y0(h_u_cla24_and4256_y0, h_u_cla24_and4255_y0, h_u_cla24_and4257_y0);
  and_gate and_gate_h_u_cla24_and4258_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4258_y0);
  and_gate and_gate_h_u_cla24_and4259_y0(h_u_cla24_and4258_y0, h_u_cla24_and4257_y0, h_u_cla24_and4259_y0);
  and_gate and_gate_h_u_cla24_and4260_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4260_y0);
  and_gate and_gate_h_u_cla24_and4261_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4261_y0);
  and_gate and_gate_h_u_cla24_and4262_y0(h_u_cla24_and4261_y0, h_u_cla24_and4260_y0, h_u_cla24_and4262_y0);
  and_gate and_gate_h_u_cla24_and4263_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4263_y0);
  and_gate and_gate_h_u_cla24_and4264_y0(h_u_cla24_and4263_y0, h_u_cla24_and4262_y0, h_u_cla24_and4264_y0);
  and_gate and_gate_h_u_cla24_and4265_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4265_y0);
  and_gate and_gate_h_u_cla24_and4266_y0(h_u_cla24_and4265_y0, h_u_cla24_and4264_y0, h_u_cla24_and4266_y0);
  and_gate and_gate_h_u_cla24_and4267_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4267_y0);
  and_gate and_gate_h_u_cla24_and4268_y0(h_u_cla24_and4267_y0, h_u_cla24_and4266_y0, h_u_cla24_and4268_y0);
  and_gate and_gate_h_u_cla24_and4269_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4269_y0);
  and_gate and_gate_h_u_cla24_and4270_y0(h_u_cla24_and4269_y0, h_u_cla24_and4268_y0, h_u_cla24_and4270_y0);
  and_gate and_gate_h_u_cla24_and4271_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4271_y0);
  and_gate and_gate_h_u_cla24_and4272_y0(h_u_cla24_and4271_y0, h_u_cla24_and4270_y0, h_u_cla24_and4272_y0);
  and_gate and_gate_h_u_cla24_and4273_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4273_y0);
  and_gate and_gate_h_u_cla24_and4274_y0(h_u_cla24_and4273_y0, h_u_cla24_and4272_y0, h_u_cla24_and4274_y0);
  and_gate and_gate_h_u_cla24_and4275_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4275_y0);
  and_gate and_gate_h_u_cla24_and4276_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4276_y0);
  and_gate and_gate_h_u_cla24_and4277_y0(h_u_cla24_and4276_y0, h_u_cla24_and4275_y0, h_u_cla24_and4277_y0);
  and_gate and_gate_h_u_cla24_and4278_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4278_y0);
  and_gate and_gate_h_u_cla24_and4279_y0(h_u_cla24_and4278_y0, h_u_cla24_and4277_y0, h_u_cla24_and4279_y0);
  and_gate and_gate_h_u_cla24_and4280_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4280_y0);
  and_gate and_gate_h_u_cla24_and4281_y0(h_u_cla24_and4280_y0, h_u_cla24_and4279_y0, h_u_cla24_and4281_y0);
  and_gate and_gate_h_u_cla24_and4282_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4282_y0);
  and_gate and_gate_h_u_cla24_and4283_y0(h_u_cla24_and4282_y0, h_u_cla24_and4281_y0, h_u_cla24_and4283_y0);
  and_gate and_gate_h_u_cla24_and4284_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4284_y0);
  and_gate and_gate_h_u_cla24_and4285_y0(h_u_cla24_and4284_y0, h_u_cla24_and4283_y0, h_u_cla24_and4285_y0);
  and_gate and_gate_h_u_cla24_and4286_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4286_y0);
  and_gate and_gate_h_u_cla24_and4287_y0(h_u_cla24_and4286_y0, h_u_cla24_and4285_y0, h_u_cla24_and4287_y0);
  and_gate and_gate_h_u_cla24_and4288_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4288_y0);
  and_gate and_gate_h_u_cla24_and4289_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4289_y0);
  and_gate and_gate_h_u_cla24_and4290_y0(h_u_cla24_and4289_y0, h_u_cla24_and4288_y0, h_u_cla24_and4290_y0);
  and_gate and_gate_h_u_cla24_and4291_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4291_y0);
  and_gate and_gate_h_u_cla24_and4292_y0(h_u_cla24_and4291_y0, h_u_cla24_and4290_y0, h_u_cla24_and4292_y0);
  and_gate and_gate_h_u_cla24_and4293_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4293_y0);
  and_gate and_gate_h_u_cla24_and4294_y0(h_u_cla24_and4293_y0, h_u_cla24_and4292_y0, h_u_cla24_and4294_y0);
  and_gate and_gate_h_u_cla24_and4295_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4295_y0);
  and_gate and_gate_h_u_cla24_and4296_y0(h_u_cla24_and4295_y0, h_u_cla24_and4294_y0, h_u_cla24_and4296_y0);
  and_gate and_gate_h_u_cla24_and4297_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4297_y0);
  and_gate and_gate_h_u_cla24_and4298_y0(h_u_cla24_and4297_y0, h_u_cla24_and4296_y0, h_u_cla24_and4298_y0);
  and_gate and_gate_h_u_cla24_and4299_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4299_y0);
  and_gate and_gate_h_u_cla24_and4300_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4300_y0);
  and_gate and_gate_h_u_cla24_and4301_y0(h_u_cla24_and4300_y0, h_u_cla24_and4299_y0, h_u_cla24_and4301_y0);
  and_gate and_gate_h_u_cla24_and4302_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4302_y0);
  and_gate and_gate_h_u_cla24_and4303_y0(h_u_cla24_and4302_y0, h_u_cla24_and4301_y0, h_u_cla24_and4303_y0);
  and_gate and_gate_h_u_cla24_and4304_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4304_y0);
  and_gate and_gate_h_u_cla24_and4305_y0(h_u_cla24_and4304_y0, h_u_cla24_and4303_y0, h_u_cla24_and4305_y0);
  and_gate and_gate_h_u_cla24_and4306_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4306_y0);
  and_gate and_gate_h_u_cla24_and4307_y0(h_u_cla24_and4306_y0, h_u_cla24_and4305_y0, h_u_cla24_and4307_y0);
  and_gate and_gate_h_u_cla24_and4308_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and4308_y0);
  and_gate and_gate_h_u_cla24_and4309_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and4309_y0);
  and_gate and_gate_h_u_cla24_and4310_y0(h_u_cla24_and4309_y0, h_u_cla24_and4308_y0, h_u_cla24_and4310_y0);
  and_gate and_gate_h_u_cla24_and4311_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and4311_y0);
  and_gate and_gate_h_u_cla24_and4312_y0(h_u_cla24_and4311_y0, h_u_cla24_and4310_y0, h_u_cla24_and4312_y0);
  and_gate and_gate_h_u_cla24_and4313_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and4313_y0);
  and_gate and_gate_h_u_cla24_and4314_y0(h_u_cla24_and4313_y0, h_u_cla24_and4312_y0, h_u_cla24_and4314_y0);
  and_gate and_gate_h_u_cla24_and4315_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and4315_y0);
  and_gate and_gate_h_u_cla24_and4316_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and4316_y0);
  and_gate and_gate_h_u_cla24_and4317_y0(h_u_cla24_and4316_y0, h_u_cla24_and4315_y0, h_u_cla24_and4317_y0);
  and_gate and_gate_h_u_cla24_and4318_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and4318_y0);
  and_gate and_gate_h_u_cla24_and4319_y0(h_u_cla24_and4318_y0, h_u_cla24_and4317_y0, h_u_cla24_and4319_y0);
  and_gate and_gate_h_u_cla24_and4320_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic20_y1, h_u_cla24_and4320_y0);
  and_gate and_gate_h_u_cla24_and4321_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic20_y1, h_u_cla24_and4321_y0);
  and_gate and_gate_h_u_cla24_and4322_y0(h_u_cla24_and4321_y0, h_u_cla24_and4320_y0, h_u_cla24_and4322_y0);
  and_gate and_gate_h_u_cla24_and4323_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic21_y1, h_u_cla24_and4323_y0);
  or_gate or_gate_h_u_cla24_or253_y0(h_u_cla24_and4323_y0, h_u_cla24_and3839_y0, h_u_cla24_or253_y0);
  or_gate or_gate_h_u_cla24_or254_y0(h_u_cla24_or253_y0, h_u_cla24_and3882_y0, h_u_cla24_or254_y0);
  or_gate or_gate_h_u_cla24_or255_y0(h_u_cla24_or254_y0, h_u_cla24_and3923_y0, h_u_cla24_or255_y0);
  or_gate or_gate_h_u_cla24_or256_y0(h_u_cla24_or255_y0, h_u_cla24_and3962_y0, h_u_cla24_or256_y0);
  or_gate or_gate_h_u_cla24_or257_y0(h_u_cla24_or256_y0, h_u_cla24_and3999_y0, h_u_cla24_or257_y0);
  or_gate or_gate_h_u_cla24_or258_y0(h_u_cla24_or257_y0, h_u_cla24_and4034_y0, h_u_cla24_or258_y0);
  or_gate or_gate_h_u_cla24_or259_y0(h_u_cla24_or258_y0, h_u_cla24_and4067_y0, h_u_cla24_or259_y0);
  or_gate or_gate_h_u_cla24_or260_y0(h_u_cla24_or259_y0, h_u_cla24_and4098_y0, h_u_cla24_or260_y0);
  or_gate or_gate_h_u_cla24_or261_y0(h_u_cla24_or260_y0, h_u_cla24_and4127_y0, h_u_cla24_or261_y0);
  or_gate or_gate_h_u_cla24_or262_y0(h_u_cla24_or261_y0, h_u_cla24_and4154_y0, h_u_cla24_or262_y0);
  or_gate or_gate_h_u_cla24_or263_y0(h_u_cla24_or262_y0, h_u_cla24_and4179_y0, h_u_cla24_or263_y0);
  or_gate or_gate_h_u_cla24_or264_y0(h_u_cla24_or263_y0, h_u_cla24_and4202_y0, h_u_cla24_or264_y0);
  or_gate or_gate_h_u_cla24_or265_y0(h_u_cla24_or264_y0, h_u_cla24_and4223_y0, h_u_cla24_or265_y0);
  or_gate or_gate_h_u_cla24_or266_y0(h_u_cla24_or265_y0, h_u_cla24_and4242_y0, h_u_cla24_or266_y0);
  or_gate or_gate_h_u_cla24_or267_y0(h_u_cla24_or266_y0, h_u_cla24_and4259_y0, h_u_cla24_or267_y0);
  or_gate or_gate_h_u_cla24_or268_y0(h_u_cla24_or267_y0, h_u_cla24_and4274_y0, h_u_cla24_or268_y0);
  or_gate or_gate_h_u_cla24_or269_y0(h_u_cla24_or268_y0, h_u_cla24_and4287_y0, h_u_cla24_or269_y0);
  or_gate or_gate_h_u_cla24_or270_y0(h_u_cla24_or269_y0, h_u_cla24_and4298_y0, h_u_cla24_or270_y0);
  or_gate or_gate_h_u_cla24_or271_y0(h_u_cla24_or270_y0, h_u_cla24_and4307_y0, h_u_cla24_or271_y0);
  or_gate or_gate_h_u_cla24_or272_y0(h_u_cla24_or271_y0, h_u_cla24_and4314_y0, h_u_cla24_or272_y0);
  or_gate or_gate_h_u_cla24_or273_y0(h_u_cla24_or272_y0, h_u_cla24_and4319_y0, h_u_cla24_or273_y0);
  or_gate or_gate_h_u_cla24_or274_y0(h_u_cla24_or273_y0, h_u_cla24_and4322_y0, h_u_cla24_or274_y0);
  or_gate or_gate_h_u_cla24_or275_y0(h_u_cla24_pg_logic22_y1, h_u_cla24_or274_y0, h_u_cla24_or275_y0);
  pg_logic pg_logic_h_u_cla24_pg_logic23_y0(a_23, b_23, h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic23_y1, h_u_cla24_pg_logic23_y2);
  xor_gate xor_gate_h_u_cla24_xor23_y0(h_u_cla24_pg_logic23_y2, h_u_cla24_or275_y0, h_u_cla24_xor23_y0);
  and_gate and_gate_h_u_cla24_and4324_y0(h_u_cla24_pg_logic0_y0, constant_wire_0, h_u_cla24_and4324_y0);
  and_gate and_gate_h_u_cla24_and4325_y0(h_u_cla24_pg_logic1_y0, constant_wire_0, h_u_cla24_and4325_y0);
  and_gate and_gate_h_u_cla24_and4326_y0(h_u_cla24_and4325_y0, h_u_cla24_and4324_y0, h_u_cla24_and4326_y0);
  and_gate and_gate_h_u_cla24_and4327_y0(h_u_cla24_pg_logic2_y0, constant_wire_0, h_u_cla24_and4327_y0);
  and_gate and_gate_h_u_cla24_and4328_y0(h_u_cla24_and4327_y0, h_u_cla24_and4326_y0, h_u_cla24_and4328_y0);
  and_gate and_gate_h_u_cla24_and4329_y0(h_u_cla24_pg_logic3_y0, constant_wire_0, h_u_cla24_and4329_y0);
  and_gate and_gate_h_u_cla24_and4330_y0(h_u_cla24_and4329_y0, h_u_cla24_and4328_y0, h_u_cla24_and4330_y0);
  and_gate and_gate_h_u_cla24_and4331_y0(h_u_cla24_pg_logic4_y0, constant_wire_0, h_u_cla24_and4331_y0);
  and_gate and_gate_h_u_cla24_and4332_y0(h_u_cla24_and4331_y0, h_u_cla24_and4330_y0, h_u_cla24_and4332_y0);
  and_gate and_gate_h_u_cla24_and4333_y0(h_u_cla24_pg_logic5_y0, constant_wire_0, h_u_cla24_and4333_y0);
  and_gate and_gate_h_u_cla24_and4334_y0(h_u_cla24_and4333_y0, h_u_cla24_and4332_y0, h_u_cla24_and4334_y0);
  and_gate and_gate_h_u_cla24_and4335_y0(h_u_cla24_pg_logic6_y0, constant_wire_0, h_u_cla24_and4335_y0);
  and_gate and_gate_h_u_cla24_and4336_y0(h_u_cla24_and4335_y0, h_u_cla24_and4334_y0, h_u_cla24_and4336_y0);
  and_gate and_gate_h_u_cla24_and4337_y0(h_u_cla24_pg_logic7_y0, constant_wire_0, h_u_cla24_and4337_y0);
  and_gate and_gate_h_u_cla24_and4338_y0(h_u_cla24_and4337_y0, h_u_cla24_and4336_y0, h_u_cla24_and4338_y0);
  and_gate and_gate_h_u_cla24_and4339_y0(h_u_cla24_pg_logic8_y0, constant_wire_0, h_u_cla24_and4339_y0);
  and_gate and_gate_h_u_cla24_and4340_y0(h_u_cla24_and4339_y0, h_u_cla24_and4338_y0, h_u_cla24_and4340_y0);
  and_gate and_gate_h_u_cla24_and4341_y0(h_u_cla24_pg_logic9_y0, constant_wire_0, h_u_cla24_and4341_y0);
  and_gate and_gate_h_u_cla24_and4342_y0(h_u_cla24_and4341_y0, h_u_cla24_and4340_y0, h_u_cla24_and4342_y0);
  and_gate and_gate_h_u_cla24_and4343_y0(h_u_cla24_pg_logic10_y0, constant_wire_0, h_u_cla24_and4343_y0);
  and_gate and_gate_h_u_cla24_and4344_y0(h_u_cla24_and4343_y0, h_u_cla24_and4342_y0, h_u_cla24_and4344_y0);
  and_gate and_gate_h_u_cla24_and4345_y0(h_u_cla24_pg_logic11_y0, constant_wire_0, h_u_cla24_and4345_y0);
  and_gate and_gate_h_u_cla24_and4346_y0(h_u_cla24_and4345_y0, h_u_cla24_and4344_y0, h_u_cla24_and4346_y0);
  and_gate and_gate_h_u_cla24_and4347_y0(h_u_cla24_pg_logic12_y0, constant_wire_0, h_u_cla24_and4347_y0);
  and_gate and_gate_h_u_cla24_and4348_y0(h_u_cla24_and4347_y0, h_u_cla24_and4346_y0, h_u_cla24_and4348_y0);
  and_gate and_gate_h_u_cla24_and4349_y0(h_u_cla24_pg_logic13_y0, constant_wire_0, h_u_cla24_and4349_y0);
  and_gate and_gate_h_u_cla24_and4350_y0(h_u_cla24_and4349_y0, h_u_cla24_and4348_y0, h_u_cla24_and4350_y0);
  and_gate and_gate_h_u_cla24_and4351_y0(h_u_cla24_pg_logic14_y0, constant_wire_0, h_u_cla24_and4351_y0);
  and_gate and_gate_h_u_cla24_and4352_y0(h_u_cla24_and4351_y0, h_u_cla24_and4350_y0, h_u_cla24_and4352_y0);
  and_gate and_gate_h_u_cla24_and4353_y0(h_u_cla24_pg_logic15_y0, constant_wire_0, h_u_cla24_and4353_y0);
  and_gate and_gate_h_u_cla24_and4354_y0(h_u_cla24_and4353_y0, h_u_cla24_and4352_y0, h_u_cla24_and4354_y0);
  and_gate and_gate_h_u_cla24_and4355_y0(h_u_cla24_pg_logic16_y0, constant_wire_0, h_u_cla24_and4355_y0);
  and_gate and_gate_h_u_cla24_and4356_y0(h_u_cla24_and4355_y0, h_u_cla24_and4354_y0, h_u_cla24_and4356_y0);
  and_gate and_gate_h_u_cla24_and4357_y0(h_u_cla24_pg_logic17_y0, constant_wire_0, h_u_cla24_and4357_y0);
  and_gate and_gate_h_u_cla24_and4358_y0(h_u_cla24_and4357_y0, h_u_cla24_and4356_y0, h_u_cla24_and4358_y0);
  and_gate and_gate_h_u_cla24_and4359_y0(h_u_cla24_pg_logic18_y0, constant_wire_0, h_u_cla24_and4359_y0);
  and_gate and_gate_h_u_cla24_and4360_y0(h_u_cla24_and4359_y0, h_u_cla24_and4358_y0, h_u_cla24_and4360_y0);
  and_gate and_gate_h_u_cla24_and4361_y0(h_u_cla24_pg_logic19_y0, constant_wire_0, h_u_cla24_and4361_y0);
  and_gate and_gate_h_u_cla24_and4362_y0(h_u_cla24_and4361_y0, h_u_cla24_and4360_y0, h_u_cla24_and4362_y0);
  and_gate and_gate_h_u_cla24_and4363_y0(h_u_cla24_pg_logic20_y0, constant_wire_0, h_u_cla24_and4363_y0);
  and_gate and_gate_h_u_cla24_and4364_y0(h_u_cla24_and4363_y0, h_u_cla24_and4362_y0, h_u_cla24_and4364_y0);
  and_gate and_gate_h_u_cla24_and4365_y0(h_u_cla24_pg_logic21_y0, constant_wire_0, h_u_cla24_and4365_y0);
  and_gate and_gate_h_u_cla24_and4366_y0(h_u_cla24_and4365_y0, h_u_cla24_and4364_y0, h_u_cla24_and4366_y0);
  and_gate and_gate_h_u_cla24_and4367_y0(h_u_cla24_pg_logic22_y0, constant_wire_0, h_u_cla24_and4367_y0);
  and_gate and_gate_h_u_cla24_and4368_y0(h_u_cla24_and4367_y0, h_u_cla24_and4366_y0, h_u_cla24_and4368_y0);
  and_gate and_gate_h_u_cla24_and4369_y0(h_u_cla24_pg_logic23_y0, constant_wire_0, h_u_cla24_and4369_y0);
  and_gate and_gate_h_u_cla24_and4370_y0(h_u_cla24_and4369_y0, h_u_cla24_and4368_y0, h_u_cla24_and4370_y0);
  and_gate and_gate_h_u_cla24_and4371_y0(h_u_cla24_pg_logic1_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4371_y0);
  and_gate and_gate_h_u_cla24_and4372_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4372_y0);
  and_gate and_gate_h_u_cla24_and4373_y0(h_u_cla24_and4372_y0, h_u_cla24_and4371_y0, h_u_cla24_and4373_y0);
  and_gate and_gate_h_u_cla24_and4374_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4374_y0);
  and_gate and_gate_h_u_cla24_and4375_y0(h_u_cla24_and4374_y0, h_u_cla24_and4373_y0, h_u_cla24_and4375_y0);
  and_gate and_gate_h_u_cla24_and4376_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4376_y0);
  and_gate and_gate_h_u_cla24_and4377_y0(h_u_cla24_and4376_y0, h_u_cla24_and4375_y0, h_u_cla24_and4377_y0);
  and_gate and_gate_h_u_cla24_and4378_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4378_y0);
  and_gate and_gate_h_u_cla24_and4379_y0(h_u_cla24_and4378_y0, h_u_cla24_and4377_y0, h_u_cla24_and4379_y0);
  and_gate and_gate_h_u_cla24_and4380_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4380_y0);
  and_gate and_gate_h_u_cla24_and4381_y0(h_u_cla24_and4380_y0, h_u_cla24_and4379_y0, h_u_cla24_and4381_y0);
  and_gate and_gate_h_u_cla24_and4382_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4382_y0);
  and_gate and_gate_h_u_cla24_and4383_y0(h_u_cla24_and4382_y0, h_u_cla24_and4381_y0, h_u_cla24_and4383_y0);
  and_gate and_gate_h_u_cla24_and4384_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4384_y0);
  and_gate and_gate_h_u_cla24_and4385_y0(h_u_cla24_and4384_y0, h_u_cla24_and4383_y0, h_u_cla24_and4385_y0);
  and_gate and_gate_h_u_cla24_and4386_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4386_y0);
  and_gate and_gate_h_u_cla24_and4387_y0(h_u_cla24_and4386_y0, h_u_cla24_and4385_y0, h_u_cla24_and4387_y0);
  and_gate and_gate_h_u_cla24_and4388_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4388_y0);
  and_gate and_gate_h_u_cla24_and4389_y0(h_u_cla24_and4388_y0, h_u_cla24_and4387_y0, h_u_cla24_and4389_y0);
  and_gate and_gate_h_u_cla24_and4390_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4390_y0);
  and_gate and_gate_h_u_cla24_and4391_y0(h_u_cla24_and4390_y0, h_u_cla24_and4389_y0, h_u_cla24_and4391_y0);
  and_gate and_gate_h_u_cla24_and4392_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4392_y0);
  and_gate and_gate_h_u_cla24_and4393_y0(h_u_cla24_and4392_y0, h_u_cla24_and4391_y0, h_u_cla24_and4393_y0);
  and_gate and_gate_h_u_cla24_and4394_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4394_y0);
  and_gate and_gate_h_u_cla24_and4395_y0(h_u_cla24_and4394_y0, h_u_cla24_and4393_y0, h_u_cla24_and4395_y0);
  and_gate and_gate_h_u_cla24_and4396_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4396_y0);
  and_gate and_gate_h_u_cla24_and4397_y0(h_u_cla24_and4396_y0, h_u_cla24_and4395_y0, h_u_cla24_and4397_y0);
  and_gate and_gate_h_u_cla24_and4398_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4398_y0);
  and_gate and_gate_h_u_cla24_and4399_y0(h_u_cla24_and4398_y0, h_u_cla24_and4397_y0, h_u_cla24_and4399_y0);
  and_gate and_gate_h_u_cla24_and4400_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4400_y0);
  and_gate and_gate_h_u_cla24_and4401_y0(h_u_cla24_and4400_y0, h_u_cla24_and4399_y0, h_u_cla24_and4401_y0);
  and_gate and_gate_h_u_cla24_and4402_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4402_y0);
  and_gate and_gate_h_u_cla24_and4403_y0(h_u_cla24_and4402_y0, h_u_cla24_and4401_y0, h_u_cla24_and4403_y0);
  and_gate and_gate_h_u_cla24_and4404_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4404_y0);
  and_gate and_gate_h_u_cla24_and4405_y0(h_u_cla24_and4404_y0, h_u_cla24_and4403_y0, h_u_cla24_and4405_y0);
  and_gate and_gate_h_u_cla24_and4406_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4406_y0);
  and_gate and_gate_h_u_cla24_and4407_y0(h_u_cla24_and4406_y0, h_u_cla24_and4405_y0, h_u_cla24_and4407_y0);
  and_gate and_gate_h_u_cla24_and4408_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4408_y0);
  and_gate and_gate_h_u_cla24_and4409_y0(h_u_cla24_and4408_y0, h_u_cla24_and4407_y0, h_u_cla24_and4409_y0);
  and_gate and_gate_h_u_cla24_and4410_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4410_y0);
  and_gate and_gate_h_u_cla24_and4411_y0(h_u_cla24_and4410_y0, h_u_cla24_and4409_y0, h_u_cla24_and4411_y0);
  and_gate and_gate_h_u_cla24_and4412_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4412_y0);
  and_gate and_gate_h_u_cla24_and4413_y0(h_u_cla24_and4412_y0, h_u_cla24_and4411_y0, h_u_cla24_and4413_y0);
  and_gate and_gate_h_u_cla24_and4414_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic0_y1, h_u_cla24_and4414_y0);
  and_gate and_gate_h_u_cla24_and4415_y0(h_u_cla24_and4414_y0, h_u_cla24_and4413_y0, h_u_cla24_and4415_y0);
  and_gate and_gate_h_u_cla24_and4416_y0(h_u_cla24_pg_logic2_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4416_y0);
  and_gate and_gate_h_u_cla24_and4417_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4417_y0);
  and_gate and_gate_h_u_cla24_and4418_y0(h_u_cla24_and4417_y0, h_u_cla24_and4416_y0, h_u_cla24_and4418_y0);
  and_gate and_gate_h_u_cla24_and4419_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4419_y0);
  and_gate and_gate_h_u_cla24_and4420_y0(h_u_cla24_and4419_y0, h_u_cla24_and4418_y0, h_u_cla24_and4420_y0);
  and_gate and_gate_h_u_cla24_and4421_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4421_y0);
  and_gate and_gate_h_u_cla24_and4422_y0(h_u_cla24_and4421_y0, h_u_cla24_and4420_y0, h_u_cla24_and4422_y0);
  and_gate and_gate_h_u_cla24_and4423_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4423_y0);
  and_gate and_gate_h_u_cla24_and4424_y0(h_u_cla24_and4423_y0, h_u_cla24_and4422_y0, h_u_cla24_and4424_y0);
  and_gate and_gate_h_u_cla24_and4425_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4425_y0);
  and_gate and_gate_h_u_cla24_and4426_y0(h_u_cla24_and4425_y0, h_u_cla24_and4424_y0, h_u_cla24_and4426_y0);
  and_gate and_gate_h_u_cla24_and4427_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4427_y0);
  and_gate and_gate_h_u_cla24_and4428_y0(h_u_cla24_and4427_y0, h_u_cla24_and4426_y0, h_u_cla24_and4428_y0);
  and_gate and_gate_h_u_cla24_and4429_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4429_y0);
  and_gate and_gate_h_u_cla24_and4430_y0(h_u_cla24_and4429_y0, h_u_cla24_and4428_y0, h_u_cla24_and4430_y0);
  and_gate and_gate_h_u_cla24_and4431_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4431_y0);
  and_gate and_gate_h_u_cla24_and4432_y0(h_u_cla24_and4431_y0, h_u_cla24_and4430_y0, h_u_cla24_and4432_y0);
  and_gate and_gate_h_u_cla24_and4433_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4433_y0);
  and_gate and_gate_h_u_cla24_and4434_y0(h_u_cla24_and4433_y0, h_u_cla24_and4432_y0, h_u_cla24_and4434_y0);
  and_gate and_gate_h_u_cla24_and4435_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4435_y0);
  and_gate and_gate_h_u_cla24_and4436_y0(h_u_cla24_and4435_y0, h_u_cla24_and4434_y0, h_u_cla24_and4436_y0);
  and_gate and_gate_h_u_cla24_and4437_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4437_y0);
  and_gate and_gate_h_u_cla24_and4438_y0(h_u_cla24_and4437_y0, h_u_cla24_and4436_y0, h_u_cla24_and4438_y0);
  and_gate and_gate_h_u_cla24_and4439_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4439_y0);
  and_gate and_gate_h_u_cla24_and4440_y0(h_u_cla24_and4439_y0, h_u_cla24_and4438_y0, h_u_cla24_and4440_y0);
  and_gate and_gate_h_u_cla24_and4441_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4441_y0);
  and_gate and_gate_h_u_cla24_and4442_y0(h_u_cla24_and4441_y0, h_u_cla24_and4440_y0, h_u_cla24_and4442_y0);
  and_gate and_gate_h_u_cla24_and4443_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4443_y0);
  and_gate and_gate_h_u_cla24_and4444_y0(h_u_cla24_and4443_y0, h_u_cla24_and4442_y0, h_u_cla24_and4444_y0);
  and_gate and_gate_h_u_cla24_and4445_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4445_y0);
  and_gate and_gate_h_u_cla24_and4446_y0(h_u_cla24_and4445_y0, h_u_cla24_and4444_y0, h_u_cla24_and4446_y0);
  and_gate and_gate_h_u_cla24_and4447_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4447_y0);
  and_gate and_gate_h_u_cla24_and4448_y0(h_u_cla24_and4447_y0, h_u_cla24_and4446_y0, h_u_cla24_and4448_y0);
  and_gate and_gate_h_u_cla24_and4449_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4449_y0);
  and_gate and_gate_h_u_cla24_and4450_y0(h_u_cla24_and4449_y0, h_u_cla24_and4448_y0, h_u_cla24_and4450_y0);
  and_gate and_gate_h_u_cla24_and4451_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4451_y0);
  and_gate and_gate_h_u_cla24_and4452_y0(h_u_cla24_and4451_y0, h_u_cla24_and4450_y0, h_u_cla24_and4452_y0);
  and_gate and_gate_h_u_cla24_and4453_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4453_y0);
  and_gate and_gate_h_u_cla24_and4454_y0(h_u_cla24_and4453_y0, h_u_cla24_and4452_y0, h_u_cla24_and4454_y0);
  and_gate and_gate_h_u_cla24_and4455_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4455_y0);
  and_gate and_gate_h_u_cla24_and4456_y0(h_u_cla24_and4455_y0, h_u_cla24_and4454_y0, h_u_cla24_and4456_y0);
  and_gate and_gate_h_u_cla24_and4457_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic1_y1, h_u_cla24_and4457_y0);
  and_gate and_gate_h_u_cla24_and4458_y0(h_u_cla24_and4457_y0, h_u_cla24_and4456_y0, h_u_cla24_and4458_y0);
  and_gate and_gate_h_u_cla24_and4459_y0(h_u_cla24_pg_logic3_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4459_y0);
  and_gate and_gate_h_u_cla24_and4460_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4460_y0);
  and_gate and_gate_h_u_cla24_and4461_y0(h_u_cla24_and4460_y0, h_u_cla24_and4459_y0, h_u_cla24_and4461_y0);
  and_gate and_gate_h_u_cla24_and4462_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4462_y0);
  and_gate and_gate_h_u_cla24_and4463_y0(h_u_cla24_and4462_y0, h_u_cla24_and4461_y0, h_u_cla24_and4463_y0);
  and_gate and_gate_h_u_cla24_and4464_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4464_y0);
  and_gate and_gate_h_u_cla24_and4465_y0(h_u_cla24_and4464_y0, h_u_cla24_and4463_y0, h_u_cla24_and4465_y0);
  and_gate and_gate_h_u_cla24_and4466_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4466_y0);
  and_gate and_gate_h_u_cla24_and4467_y0(h_u_cla24_and4466_y0, h_u_cla24_and4465_y0, h_u_cla24_and4467_y0);
  and_gate and_gate_h_u_cla24_and4468_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4468_y0);
  and_gate and_gate_h_u_cla24_and4469_y0(h_u_cla24_and4468_y0, h_u_cla24_and4467_y0, h_u_cla24_and4469_y0);
  and_gate and_gate_h_u_cla24_and4470_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4470_y0);
  and_gate and_gate_h_u_cla24_and4471_y0(h_u_cla24_and4470_y0, h_u_cla24_and4469_y0, h_u_cla24_and4471_y0);
  and_gate and_gate_h_u_cla24_and4472_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4472_y0);
  and_gate and_gate_h_u_cla24_and4473_y0(h_u_cla24_and4472_y0, h_u_cla24_and4471_y0, h_u_cla24_and4473_y0);
  and_gate and_gate_h_u_cla24_and4474_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4474_y0);
  and_gate and_gate_h_u_cla24_and4475_y0(h_u_cla24_and4474_y0, h_u_cla24_and4473_y0, h_u_cla24_and4475_y0);
  and_gate and_gate_h_u_cla24_and4476_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4476_y0);
  and_gate and_gate_h_u_cla24_and4477_y0(h_u_cla24_and4476_y0, h_u_cla24_and4475_y0, h_u_cla24_and4477_y0);
  and_gate and_gate_h_u_cla24_and4478_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4478_y0);
  and_gate and_gate_h_u_cla24_and4479_y0(h_u_cla24_and4478_y0, h_u_cla24_and4477_y0, h_u_cla24_and4479_y0);
  and_gate and_gate_h_u_cla24_and4480_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4480_y0);
  and_gate and_gate_h_u_cla24_and4481_y0(h_u_cla24_and4480_y0, h_u_cla24_and4479_y0, h_u_cla24_and4481_y0);
  and_gate and_gate_h_u_cla24_and4482_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4482_y0);
  and_gate and_gate_h_u_cla24_and4483_y0(h_u_cla24_and4482_y0, h_u_cla24_and4481_y0, h_u_cla24_and4483_y0);
  and_gate and_gate_h_u_cla24_and4484_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4484_y0);
  and_gate and_gate_h_u_cla24_and4485_y0(h_u_cla24_and4484_y0, h_u_cla24_and4483_y0, h_u_cla24_and4485_y0);
  and_gate and_gate_h_u_cla24_and4486_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4486_y0);
  and_gate and_gate_h_u_cla24_and4487_y0(h_u_cla24_and4486_y0, h_u_cla24_and4485_y0, h_u_cla24_and4487_y0);
  and_gate and_gate_h_u_cla24_and4488_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4488_y0);
  and_gate and_gate_h_u_cla24_and4489_y0(h_u_cla24_and4488_y0, h_u_cla24_and4487_y0, h_u_cla24_and4489_y0);
  and_gate and_gate_h_u_cla24_and4490_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4490_y0);
  and_gate and_gate_h_u_cla24_and4491_y0(h_u_cla24_and4490_y0, h_u_cla24_and4489_y0, h_u_cla24_and4491_y0);
  and_gate and_gate_h_u_cla24_and4492_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4492_y0);
  and_gate and_gate_h_u_cla24_and4493_y0(h_u_cla24_and4492_y0, h_u_cla24_and4491_y0, h_u_cla24_and4493_y0);
  and_gate and_gate_h_u_cla24_and4494_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4494_y0);
  and_gate and_gate_h_u_cla24_and4495_y0(h_u_cla24_and4494_y0, h_u_cla24_and4493_y0, h_u_cla24_and4495_y0);
  and_gate and_gate_h_u_cla24_and4496_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4496_y0);
  and_gate and_gate_h_u_cla24_and4497_y0(h_u_cla24_and4496_y0, h_u_cla24_and4495_y0, h_u_cla24_and4497_y0);
  and_gate and_gate_h_u_cla24_and4498_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic2_y1, h_u_cla24_and4498_y0);
  and_gate and_gate_h_u_cla24_and4499_y0(h_u_cla24_and4498_y0, h_u_cla24_and4497_y0, h_u_cla24_and4499_y0);
  and_gate and_gate_h_u_cla24_and4500_y0(h_u_cla24_pg_logic4_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4500_y0);
  and_gate and_gate_h_u_cla24_and4501_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4501_y0);
  and_gate and_gate_h_u_cla24_and4502_y0(h_u_cla24_and4501_y0, h_u_cla24_and4500_y0, h_u_cla24_and4502_y0);
  and_gate and_gate_h_u_cla24_and4503_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4503_y0);
  and_gate and_gate_h_u_cla24_and4504_y0(h_u_cla24_and4503_y0, h_u_cla24_and4502_y0, h_u_cla24_and4504_y0);
  and_gate and_gate_h_u_cla24_and4505_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4505_y0);
  and_gate and_gate_h_u_cla24_and4506_y0(h_u_cla24_and4505_y0, h_u_cla24_and4504_y0, h_u_cla24_and4506_y0);
  and_gate and_gate_h_u_cla24_and4507_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4507_y0);
  and_gate and_gate_h_u_cla24_and4508_y0(h_u_cla24_and4507_y0, h_u_cla24_and4506_y0, h_u_cla24_and4508_y0);
  and_gate and_gate_h_u_cla24_and4509_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4509_y0);
  and_gate and_gate_h_u_cla24_and4510_y0(h_u_cla24_and4509_y0, h_u_cla24_and4508_y0, h_u_cla24_and4510_y0);
  and_gate and_gate_h_u_cla24_and4511_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4511_y0);
  and_gate and_gate_h_u_cla24_and4512_y0(h_u_cla24_and4511_y0, h_u_cla24_and4510_y0, h_u_cla24_and4512_y0);
  and_gate and_gate_h_u_cla24_and4513_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4513_y0);
  and_gate and_gate_h_u_cla24_and4514_y0(h_u_cla24_and4513_y0, h_u_cla24_and4512_y0, h_u_cla24_and4514_y0);
  and_gate and_gate_h_u_cla24_and4515_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4515_y0);
  and_gate and_gate_h_u_cla24_and4516_y0(h_u_cla24_and4515_y0, h_u_cla24_and4514_y0, h_u_cla24_and4516_y0);
  and_gate and_gate_h_u_cla24_and4517_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4517_y0);
  and_gate and_gate_h_u_cla24_and4518_y0(h_u_cla24_and4517_y0, h_u_cla24_and4516_y0, h_u_cla24_and4518_y0);
  and_gate and_gate_h_u_cla24_and4519_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4519_y0);
  and_gate and_gate_h_u_cla24_and4520_y0(h_u_cla24_and4519_y0, h_u_cla24_and4518_y0, h_u_cla24_and4520_y0);
  and_gate and_gate_h_u_cla24_and4521_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4521_y0);
  and_gate and_gate_h_u_cla24_and4522_y0(h_u_cla24_and4521_y0, h_u_cla24_and4520_y0, h_u_cla24_and4522_y0);
  and_gate and_gate_h_u_cla24_and4523_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4523_y0);
  and_gate and_gate_h_u_cla24_and4524_y0(h_u_cla24_and4523_y0, h_u_cla24_and4522_y0, h_u_cla24_and4524_y0);
  and_gate and_gate_h_u_cla24_and4525_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4525_y0);
  and_gate and_gate_h_u_cla24_and4526_y0(h_u_cla24_and4525_y0, h_u_cla24_and4524_y0, h_u_cla24_and4526_y0);
  and_gate and_gate_h_u_cla24_and4527_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4527_y0);
  and_gate and_gate_h_u_cla24_and4528_y0(h_u_cla24_and4527_y0, h_u_cla24_and4526_y0, h_u_cla24_and4528_y0);
  and_gate and_gate_h_u_cla24_and4529_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4529_y0);
  and_gate and_gate_h_u_cla24_and4530_y0(h_u_cla24_and4529_y0, h_u_cla24_and4528_y0, h_u_cla24_and4530_y0);
  and_gate and_gate_h_u_cla24_and4531_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4531_y0);
  and_gate and_gate_h_u_cla24_and4532_y0(h_u_cla24_and4531_y0, h_u_cla24_and4530_y0, h_u_cla24_and4532_y0);
  and_gate and_gate_h_u_cla24_and4533_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4533_y0);
  and_gate and_gate_h_u_cla24_and4534_y0(h_u_cla24_and4533_y0, h_u_cla24_and4532_y0, h_u_cla24_and4534_y0);
  and_gate and_gate_h_u_cla24_and4535_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4535_y0);
  and_gate and_gate_h_u_cla24_and4536_y0(h_u_cla24_and4535_y0, h_u_cla24_and4534_y0, h_u_cla24_and4536_y0);
  and_gate and_gate_h_u_cla24_and4537_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic3_y1, h_u_cla24_and4537_y0);
  and_gate and_gate_h_u_cla24_and4538_y0(h_u_cla24_and4537_y0, h_u_cla24_and4536_y0, h_u_cla24_and4538_y0);
  and_gate and_gate_h_u_cla24_and4539_y0(h_u_cla24_pg_logic5_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4539_y0);
  and_gate and_gate_h_u_cla24_and4540_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4540_y0);
  and_gate and_gate_h_u_cla24_and4541_y0(h_u_cla24_and4540_y0, h_u_cla24_and4539_y0, h_u_cla24_and4541_y0);
  and_gate and_gate_h_u_cla24_and4542_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4542_y0);
  and_gate and_gate_h_u_cla24_and4543_y0(h_u_cla24_and4542_y0, h_u_cla24_and4541_y0, h_u_cla24_and4543_y0);
  and_gate and_gate_h_u_cla24_and4544_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4544_y0);
  and_gate and_gate_h_u_cla24_and4545_y0(h_u_cla24_and4544_y0, h_u_cla24_and4543_y0, h_u_cla24_and4545_y0);
  and_gate and_gate_h_u_cla24_and4546_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4546_y0);
  and_gate and_gate_h_u_cla24_and4547_y0(h_u_cla24_and4546_y0, h_u_cla24_and4545_y0, h_u_cla24_and4547_y0);
  and_gate and_gate_h_u_cla24_and4548_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4548_y0);
  and_gate and_gate_h_u_cla24_and4549_y0(h_u_cla24_and4548_y0, h_u_cla24_and4547_y0, h_u_cla24_and4549_y0);
  and_gate and_gate_h_u_cla24_and4550_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4550_y0);
  and_gate and_gate_h_u_cla24_and4551_y0(h_u_cla24_and4550_y0, h_u_cla24_and4549_y0, h_u_cla24_and4551_y0);
  and_gate and_gate_h_u_cla24_and4552_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4552_y0);
  and_gate and_gate_h_u_cla24_and4553_y0(h_u_cla24_and4552_y0, h_u_cla24_and4551_y0, h_u_cla24_and4553_y0);
  and_gate and_gate_h_u_cla24_and4554_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4554_y0);
  and_gate and_gate_h_u_cla24_and4555_y0(h_u_cla24_and4554_y0, h_u_cla24_and4553_y0, h_u_cla24_and4555_y0);
  and_gate and_gate_h_u_cla24_and4556_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4556_y0);
  and_gate and_gate_h_u_cla24_and4557_y0(h_u_cla24_and4556_y0, h_u_cla24_and4555_y0, h_u_cla24_and4557_y0);
  and_gate and_gate_h_u_cla24_and4558_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4558_y0);
  and_gate and_gate_h_u_cla24_and4559_y0(h_u_cla24_and4558_y0, h_u_cla24_and4557_y0, h_u_cla24_and4559_y0);
  and_gate and_gate_h_u_cla24_and4560_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4560_y0);
  and_gate and_gate_h_u_cla24_and4561_y0(h_u_cla24_and4560_y0, h_u_cla24_and4559_y0, h_u_cla24_and4561_y0);
  and_gate and_gate_h_u_cla24_and4562_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4562_y0);
  and_gate and_gate_h_u_cla24_and4563_y0(h_u_cla24_and4562_y0, h_u_cla24_and4561_y0, h_u_cla24_and4563_y0);
  and_gate and_gate_h_u_cla24_and4564_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4564_y0);
  and_gate and_gate_h_u_cla24_and4565_y0(h_u_cla24_and4564_y0, h_u_cla24_and4563_y0, h_u_cla24_and4565_y0);
  and_gate and_gate_h_u_cla24_and4566_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4566_y0);
  and_gate and_gate_h_u_cla24_and4567_y0(h_u_cla24_and4566_y0, h_u_cla24_and4565_y0, h_u_cla24_and4567_y0);
  and_gate and_gate_h_u_cla24_and4568_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4568_y0);
  and_gate and_gate_h_u_cla24_and4569_y0(h_u_cla24_and4568_y0, h_u_cla24_and4567_y0, h_u_cla24_and4569_y0);
  and_gate and_gate_h_u_cla24_and4570_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4570_y0);
  and_gate and_gate_h_u_cla24_and4571_y0(h_u_cla24_and4570_y0, h_u_cla24_and4569_y0, h_u_cla24_and4571_y0);
  and_gate and_gate_h_u_cla24_and4572_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4572_y0);
  and_gate and_gate_h_u_cla24_and4573_y0(h_u_cla24_and4572_y0, h_u_cla24_and4571_y0, h_u_cla24_and4573_y0);
  and_gate and_gate_h_u_cla24_and4574_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic4_y1, h_u_cla24_and4574_y0);
  and_gate and_gate_h_u_cla24_and4575_y0(h_u_cla24_and4574_y0, h_u_cla24_and4573_y0, h_u_cla24_and4575_y0);
  and_gate and_gate_h_u_cla24_and4576_y0(h_u_cla24_pg_logic6_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4576_y0);
  and_gate and_gate_h_u_cla24_and4577_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4577_y0);
  and_gate and_gate_h_u_cla24_and4578_y0(h_u_cla24_and4577_y0, h_u_cla24_and4576_y0, h_u_cla24_and4578_y0);
  and_gate and_gate_h_u_cla24_and4579_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4579_y0);
  and_gate and_gate_h_u_cla24_and4580_y0(h_u_cla24_and4579_y0, h_u_cla24_and4578_y0, h_u_cla24_and4580_y0);
  and_gate and_gate_h_u_cla24_and4581_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4581_y0);
  and_gate and_gate_h_u_cla24_and4582_y0(h_u_cla24_and4581_y0, h_u_cla24_and4580_y0, h_u_cla24_and4582_y0);
  and_gate and_gate_h_u_cla24_and4583_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4583_y0);
  and_gate and_gate_h_u_cla24_and4584_y0(h_u_cla24_and4583_y0, h_u_cla24_and4582_y0, h_u_cla24_and4584_y0);
  and_gate and_gate_h_u_cla24_and4585_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4585_y0);
  and_gate and_gate_h_u_cla24_and4586_y0(h_u_cla24_and4585_y0, h_u_cla24_and4584_y0, h_u_cla24_and4586_y0);
  and_gate and_gate_h_u_cla24_and4587_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4587_y0);
  and_gate and_gate_h_u_cla24_and4588_y0(h_u_cla24_and4587_y0, h_u_cla24_and4586_y0, h_u_cla24_and4588_y0);
  and_gate and_gate_h_u_cla24_and4589_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4589_y0);
  and_gate and_gate_h_u_cla24_and4590_y0(h_u_cla24_and4589_y0, h_u_cla24_and4588_y0, h_u_cla24_and4590_y0);
  and_gate and_gate_h_u_cla24_and4591_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4591_y0);
  and_gate and_gate_h_u_cla24_and4592_y0(h_u_cla24_and4591_y0, h_u_cla24_and4590_y0, h_u_cla24_and4592_y0);
  and_gate and_gate_h_u_cla24_and4593_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4593_y0);
  and_gate and_gate_h_u_cla24_and4594_y0(h_u_cla24_and4593_y0, h_u_cla24_and4592_y0, h_u_cla24_and4594_y0);
  and_gate and_gate_h_u_cla24_and4595_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4595_y0);
  and_gate and_gate_h_u_cla24_and4596_y0(h_u_cla24_and4595_y0, h_u_cla24_and4594_y0, h_u_cla24_and4596_y0);
  and_gate and_gate_h_u_cla24_and4597_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4597_y0);
  and_gate and_gate_h_u_cla24_and4598_y0(h_u_cla24_and4597_y0, h_u_cla24_and4596_y0, h_u_cla24_and4598_y0);
  and_gate and_gate_h_u_cla24_and4599_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4599_y0);
  and_gate and_gate_h_u_cla24_and4600_y0(h_u_cla24_and4599_y0, h_u_cla24_and4598_y0, h_u_cla24_and4600_y0);
  and_gate and_gate_h_u_cla24_and4601_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4601_y0);
  and_gate and_gate_h_u_cla24_and4602_y0(h_u_cla24_and4601_y0, h_u_cla24_and4600_y0, h_u_cla24_and4602_y0);
  and_gate and_gate_h_u_cla24_and4603_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4603_y0);
  and_gate and_gate_h_u_cla24_and4604_y0(h_u_cla24_and4603_y0, h_u_cla24_and4602_y0, h_u_cla24_and4604_y0);
  and_gate and_gate_h_u_cla24_and4605_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4605_y0);
  and_gate and_gate_h_u_cla24_and4606_y0(h_u_cla24_and4605_y0, h_u_cla24_and4604_y0, h_u_cla24_and4606_y0);
  and_gate and_gate_h_u_cla24_and4607_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4607_y0);
  and_gate and_gate_h_u_cla24_and4608_y0(h_u_cla24_and4607_y0, h_u_cla24_and4606_y0, h_u_cla24_and4608_y0);
  and_gate and_gate_h_u_cla24_and4609_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic5_y1, h_u_cla24_and4609_y0);
  and_gate and_gate_h_u_cla24_and4610_y0(h_u_cla24_and4609_y0, h_u_cla24_and4608_y0, h_u_cla24_and4610_y0);
  and_gate and_gate_h_u_cla24_and4611_y0(h_u_cla24_pg_logic7_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4611_y0);
  and_gate and_gate_h_u_cla24_and4612_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4612_y0);
  and_gate and_gate_h_u_cla24_and4613_y0(h_u_cla24_and4612_y0, h_u_cla24_and4611_y0, h_u_cla24_and4613_y0);
  and_gate and_gate_h_u_cla24_and4614_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4614_y0);
  and_gate and_gate_h_u_cla24_and4615_y0(h_u_cla24_and4614_y0, h_u_cla24_and4613_y0, h_u_cla24_and4615_y0);
  and_gate and_gate_h_u_cla24_and4616_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4616_y0);
  and_gate and_gate_h_u_cla24_and4617_y0(h_u_cla24_and4616_y0, h_u_cla24_and4615_y0, h_u_cla24_and4617_y0);
  and_gate and_gate_h_u_cla24_and4618_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4618_y0);
  and_gate and_gate_h_u_cla24_and4619_y0(h_u_cla24_and4618_y0, h_u_cla24_and4617_y0, h_u_cla24_and4619_y0);
  and_gate and_gate_h_u_cla24_and4620_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4620_y0);
  and_gate and_gate_h_u_cla24_and4621_y0(h_u_cla24_and4620_y0, h_u_cla24_and4619_y0, h_u_cla24_and4621_y0);
  and_gate and_gate_h_u_cla24_and4622_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4622_y0);
  and_gate and_gate_h_u_cla24_and4623_y0(h_u_cla24_and4622_y0, h_u_cla24_and4621_y0, h_u_cla24_and4623_y0);
  and_gate and_gate_h_u_cla24_and4624_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4624_y0);
  and_gate and_gate_h_u_cla24_and4625_y0(h_u_cla24_and4624_y0, h_u_cla24_and4623_y0, h_u_cla24_and4625_y0);
  and_gate and_gate_h_u_cla24_and4626_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4626_y0);
  and_gate and_gate_h_u_cla24_and4627_y0(h_u_cla24_and4626_y0, h_u_cla24_and4625_y0, h_u_cla24_and4627_y0);
  and_gate and_gate_h_u_cla24_and4628_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4628_y0);
  and_gate and_gate_h_u_cla24_and4629_y0(h_u_cla24_and4628_y0, h_u_cla24_and4627_y0, h_u_cla24_and4629_y0);
  and_gate and_gate_h_u_cla24_and4630_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4630_y0);
  and_gate and_gate_h_u_cla24_and4631_y0(h_u_cla24_and4630_y0, h_u_cla24_and4629_y0, h_u_cla24_and4631_y0);
  and_gate and_gate_h_u_cla24_and4632_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4632_y0);
  and_gate and_gate_h_u_cla24_and4633_y0(h_u_cla24_and4632_y0, h_u_cla24_and4631_y0, h_u_cla24_and4633_y0);
  and_gate and_gate_h_u_cla24_and4634_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4634_y0);
  and_gate and_gate_h_u_cla24_and4635_y0(h_u_cla24_and4634_y0, h_u_cla24_and4633_y0, h_u_cla24_and4635_y0);
  and_gate and_gate_h_u_cla24_and4636_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4636_y0);
  and_gate and_gate_h_u_cla24_and4637_y0(h_u_cla24_and4636_y0, h_u_cla24_and4635_y0, h_u_cla24_and4637_y0);
  and_gate and_gate_h_u_cla24_and4638_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4638_y0);
  and_gate and_gate_h_u_cla24_and4639_y0(h_u_cla24_and4638_y0, h_u_cla24_and4637_y0, h_u_cla24_and4639_y0);
  and_gate and_gate_h_u_cla24_and4640_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4640_y0);
  and_gate and_gate_h_u_cla24_and4641_y0(h_u_cla24_and4640_y0, h_u_cla24_and4639_y0, h_u_cla24_and4641_y0);
  and_gate and_gate_h_u_cla24_and4642_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic6_y1, h_u_cla24_and4642_y0);
  and_gate and_gate_h_u_cla24_and4643_y0(h_u_cla24_and4642_y0, h_u_cla24_and4641_y0, h_u_cla24_and4643_y0);
  and_gate and_gate_h_u_cla24_and4644_y0(h_u_cla24_pg_logic8_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4644_y0);
  and_gate and_gate_h_u_cla24_and4645_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4645_y0);
  and_gate and_gate_h_u_cla24_and4646_y0(h_u_cla24_and4645_y0, h_u_cla24_and4644_y0, h_u_cla24_and4646_y0);
  and_gate and_gate_h_u_cla24_and4647_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4647_y0);
  and_gate and_gate_h_u_cla24_and4648_y0(h_u_cla24_and4647_y0, h_u_cla24_and4646_y0, h_u_cla24_and4648_y0);
  and_gate and_gate_h_u_cla24_and4649_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4649_y0);
  and_gate and_gate_h_u_cla24_and4650_y0(h_u_cla24_and4649_y0, h_u_cla24_and4648_y0, h_u_cla24_and4650_y0);
  and_gate and_gate_h_u_cla24_and4651_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4651_y0);
  and_gate and_gate_h_u_cla24_and4652_y0(h_u_cla24_and4651_y0, h_u_cla24_and4650_y0, h_u_cla24_and4652_y0);
  and_gate and_gate_h_u_cla24_and4653_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4653_y0);
  and_gate and_gate_h_u_cla24_and4654_y0(h_u_cla24_and4653_y0, h_u_cla24_and4652_y0, h_u_cla24_and4654_y0);
  and_gate and_gate_h_u_cla24_and4655_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4655_y0);
  and_gate and_gate_h_u_cla24_and4656_y0(h_u_cla24_and4655_y0, h_u_cla24_and4654_y0, h_u_cla24_and4656_y0);
  and_gate and_gate_h_u_cla24_and4657_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4657_y0);
  and_gate and_gate_h_u_cla24_and4658_y0(h_u_cla24_and4657_y0, h_u_cla24_and4656_y0, h_u_cla24_and4658_y0);
  and_gate and_gate_h_u_cla24_and4659_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4659_y0);
  and_gate and_gate_h_u_cla24_and4660_y0(h_u_cla24_and4659_y0, h_u_cla24_and4658_y0, h_u_cla24_and4660_y0);
  and_gate and_gate_h_u_cla24_and4661_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4661_y0);
  and_gate and_gate_h_u_cla24_and4662_y0(h_u_cla24_and4661_y0, h_u_cla24_and4660_y0, h_u_cla24_and4662_y0);
  and_gate and_gate_h_u_cla24_and4663_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4663_y0);
  and_gate and_gate_h_u_cla24_and4664_y0(h_u_cla24_and4663_y0, h_u_cla24_and4662_y0, h_u_cla24_and4664_y0);
  and_gate and_gate_h_u_cla24_and4665_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4665_y0);
  and_gate and_gate_h_u_cla24_and4666_y0(h_u_cla24_and4665_y0, h_u_cla24_and4664_y0, h_u_cla24_and4666_y0);
  and_gate and_gate_h_u_cla24_and4667_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4667_y0);
  and_gate and_gate_h_u_cla24_and4668_y0(h_u_cla24_and4667_y0, h_u_cla24_and4666_y0, h_u_cla24_and4668_y0);
  and_gate and_gate_h_u_cla24_and4669_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4669_y0);
  and_gate and_gate_h_u_cla24_and4670_y0(h_u_cla24_and4669_y0, h_u_cla24_and4668_y0, h_u_cla24_and4670_y0);
  and_gate and_gate_h_u_cla24_and4671_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4671_y0);
  and_gate and_gate_h_u_cla24_and4672_y0(h_u_cla24_and4671_y0, h_u_cla24_and4670_y0, h_u_cla24_and4672_y0);
  and_gate and_gate_h_u_cla24_and4673_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic7_y1, h_u_cla24_and4673_y0);
  and_gate and_gate_h_u_cla24_and4674_y0(h_u_cla24_and4673_y0, h_u_cla24_and4672_y0, h_u_cla24_and4674_y0);
  and_gate and_gate_h_u_cla24_and4675_y0(h_u_cla24_pg_logic9_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4675_y0);
  and_gate and_gate_h_u_cla24_and4676_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4676_y0);
  and_gate and_gate_h_u_cla24_and4677_y0(h_u_cla24_and4676_y0, h_u_cla24_and4675_y0, h_u_cla24_and4677_y0);
  and_gate and_gate_h_u_cla24_and4678_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4678_y0);
  and_gate and_gate_h_u_cla24_and4679_y0(h_u_cla24_and4678_y0, h_u_cla24_and4677_y0, h_u_cla24_and4679_y0);
  and_gate and_gate_h_u_cla24_and4680_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4680_y0);
  and_gate and_gate_h_u_cla24_and4681_y0(h_u_cla24_and4680_y0, h_u_cla24_and4679_y0, h_u_cla24_and4681_y0);
  and_gate and_gate_h_u_cla24_and4682_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4682_y0);
  and_gate and_gate_h_u_cla24_and4683_y0(h_u_cla24_and4682_y0, h_u_cla24_and4681_y0, h_u_cla24_and4683_y0);
  and_gate and_gate_h_u_cla24_and4684_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4684_y0);
  and_gate and_gate_h_u_cla24_and4685_y0(h_u_cla24_and4684_y0, h_u_cla24_and4683_y0, h_u_cla24_and4685_y0);
  and_gate and_gate_h_u_cla24_and4686_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4686_y0);
  and_gate and_gate_h_u_cla24_and4687_y0(h_u_cla24_and4686_y0, h_u_cla24_and4685_y0, h_u_cla24_and4687_y0);
  and_gate and_gate_h_u_cla24_and4688_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4688_y0);
  and_gate and_gate_h_u_cla24_and4689_y0(h_u_cla24_and4688_y0, h_u_cla24_and4687_y0, h_u_cla24_and4689_y0);
  and_gate and_gate_h_u_cla24_and4690_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4690_y0);
  and_gate and_gate_h_u_cla24_and4691_y0(h_u_cla24_and4690_y0, h_u_cla24_and4689_y0, h_u_cla24_and4691_y0);
  and_gate and_gate_h_u_cla24_and4692_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4692_y0);
  and_gate and_gate_h_u_cla24_and4693_y0(h_u_cla24_and4692_y0, h_u_cla24_and4691_y0, h_u_cla24_and4693_y0);
  and_gate and_gate_h_u_cla24_and4694_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4694_y0);
  and_gate and_gate_h_u_cla24_and4695_y0(h_u_cla24_and4694_y0, h_u_cla24_and4693_y0, h_u_cla24_and4695_y0);
  and_gate and_gate_h_u_cla24_and4696_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4696_y0);
  and_gate and_gate_h_u_cla24_and4697_y0(h_u_cla24_and4696_y0, h_u_cla24_and4695_y0, h_u_cla24_and4697_y0);
  and_gate and_gate_h_u_cla24_and4698_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4698_y0);
  and_gate and_gate_h_u_cla24_and4699_y0(h_u_cla24_and4698_y0, h_u_cla24_and4697_y0, h_u_cla24_and4699_y0);
  and_gate and_gate_h_u_cla24_and4700_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4700_y0);
  and_gate and_gate_h_u_cla24_and4701_y0(h_u_cla24_and4700_y0, h_u_cla24_and4699_y0, h_u_cla24_and4701_y0);
  and_gate and_gate_h_u_cla24_and4702_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic8_y1, h_u_cla24_and4702_y0);
  and_gate and_gate_h_u_cla24_and4703_y0(h_u_cla24_and4702_y0, h_u_cla24_and4701_y0, h_u_cla24_and4703_y0);
  and_gate and_gate_h_u_cla24_and4704_y0(h_u_cla24_pg_logic10_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4704_y0);
  and_gate and_gate_h_u_cla24_and4705_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4705_y0);
  and_gate and_gate_h_u_cla24_and4706_y0(h_u_cla24_and4705_y0, h_u_cla24_and4704_y0, h_u_cla24_and4706_y0);
  and_gate and_gate_h_u_cla24_and4707_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4707_y0);
  and_gate and_gate_h_u_cla24_and4708_y0(h_u_cla24_and4707_y0, h_u_cla24_and4706_y0, h_u_cla24_and4708_y0);
  and_gate and_gate_h_u_cla24_and4709_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4709_y0);
  and_gate and_gate_h_u_cla24_and4710_y0(h_u_cla24_and4709_y0, h_u_cla24_and4708_y0, h_u_cla24_and4710_y0);
  and_gate and_gate_h_u_cla24_and4711_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4711_y0);
  and_gate and_gate_h_u_cla24_and4712_y0(h_u_cla24_and4711_y0, h_u_cla24_and4710_y0, h_u_cla24_and4712_y0);
  and_gate and_gate_h_u_cla24_and4713_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4713_y0);
  and_gate and_gate_h_u_cla24_and4714_y0(h_u_cla24_and4713_y0, h_u_cla24_and4712_y0, h_u_cla24_and4714_y0);
  and_gate and_gate_h_u_cla24_and4715_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4715_y0);
  and_gate and_gate_h_u_cla24_and4716_y0(h_u_cla24_and4715_y0, h_u_cla24_and4714_y0, h_u_cla24_and4716_y0);
  and_gate and_gate_h_u_cla24_and4717_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4717_y0);
  and_gate and_gate_h_u_cla24_and4718_y0(h_u_cla24_and4717_y0, h_u_cla24_and4716_y0, h_u_cla24_and4718_y0);
  and_gate and_gate_h_u_cla24_and4719_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4719_y0);
  and_gate and_gate_h_u_cla24_and4720_y0(h_u_cla24_and4719_y0, h_u_cla24_and4718_y0, h_u_cla24_and4720_y0);
  and_gate and_gate_h_u_cla24_and4721_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4721_y0);
  and_gate and_gate_h_u_cla24_and4722_y0(h_u_cla24_and4721_y0, h_u_cla24_and4720_y0, h_u_cla24_and4722_y0);
  and_gate and_gate_h_u_cla24_and4723_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4723_y0);
  and_gate and_gate_h_u_cla24_and4724_y0(h_u_cla24_and4723_y0, h_u_cla24_and4722_y0, h_u_cla24_and4724_y0);
  and_gate and_gate_h_u_cla24_and4725_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4725_y0);
  and_gate and_gate_h_u_cla24_and4726_y0(h_u_cla24_and4725_y0, h_u_cla24_and4724_y0, h_u_cla24_and4726_y0);
  and_gate and_gate_h_u_cla24_and4727_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4727_y0);
  and_gate and_gate_h_u_cla24_and4728_y0(h_u_cla24_and4727_y0, h_u_cla24_and4726_y0, h_u_cla24_and4728_y0);
  and_gate and_gate_h_u_cla24_and4729_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic9_y1, h_u_cla24_and4729_y0);
  and_gate and_gate_h_u_cla24_and4730_y0(h_u_cla24_and4729_y0, h_u_cla24_and4728_y0, h_u_cla24_and4730_y0);
  and_gate and_gate_h_u_cla24_and4731_y0(h_u_cla24_pg_logic11_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4731_y0);
  and_gate and_gate_h_u_cla24_and4732_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4732_y0);
  and_gate and_gate_h_u_cla24_and4733_y0(h_u_cla24_and4732_y0, h_u_cla24_and4731_y0, h_u_cla24_and4733_y0);
  and_gate and_gate_h_u_cla24_and4734_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4734_y0);
  and_gate and_gate_h_u_cla24_and4735_y0(h_u_cla24_and4734_y0, h_u_cla24_and4733_y0, h_u_cla24_and4735_y0);
  and_gate and_gate_h_u_cla24_and4736_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4736_y0);
  and_gate and_gate_h_u_cla24_and4737_y0(h_u_cla24_and4736_y0, h_u_cla24_and4735_y0, h_u_cla24_and4737_y0);
  and_gate and_gate_h_u_cla24_and4738_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4738_y0);
  and_gate and_gate_h_u_cla24_and4739_y0(h_u_cla24_and4738_y0, h_u_cla24_and4737_y0, h_u_cla24_and4739_y0);
  and_gate and_gate_h_u_cla24_and4740_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4740_y0);
  and_gate and_gate_h_u_cla24_and4741_y0(h_u_cla24_and4740_y0, h_u_cla24_and4739_y0, h_u_cla24_and4741_y0);
  and_gate and_gate_h_u_cla24_and4742_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4742_y0);
  and_gate and_gate_h_u_cla24_and4743_y0(h_u_cla24_and4742_y0, h_u_cla24_and4741_y0, h_u_cla24_and4743_y0);
  and_gate and_gate_h_u_cla24_and4744_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4744_y0);
  and_gate and_gate_h_u_cla24_and4745_y0(h_u_cla24_and4744_y0, h_u_cla24_and4743_y0, h_u_cla24_and4745_y0);
  and_gate and_gate_h_u_cla24_and4746_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4746_y0);
  and_gate and_gate_h_u_cla24_and4747_y0(h_u_cla24_and4746_y0, h_u_cla24_and4745_y0, h_u_cla24_and4747_y0);
  and_gate and_gate_h_u_cla24_and4748_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4748_y0);
  and_gate and_gate_h_u_cla24_and4749_y0(h_u_cla24_and4748_y0, h_u_cla24_and4747_y0, h_u_cla24_and4749_y0);
  and_gate and_gate_h_u_cla24_and4750_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4750_y0);
  and_gate and_gate_h_u_cla24_and4751_y0(h_u_cla24_and4750_y0, h_u_cla24_and4749_y0, h_u_cla24_and4751_y0);
  and_gate and_gate_h_u_cla24_and4752_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4752_y0);
  and_gate and_gate_h_u_cla24_and4753_y0(h_u_cla24_and4752_y0, h_u_cla24_and4751_y0, h_u_cla24_and4753_y0);
  and_gate and_gate_h_u_cla24_and4754_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic10_y1, h_u_cla24_and4754_y0);
  and_gate and_gate_h_u_cla24_and4755_y0(h_u_cla24_and4754_y0, h_u_cla24_and4753_y0, h_u_cla24_and4755_y0);
  and_gate and_gate_h_u_cla24_and4756_y0(h_u_cla24_pg_logic12_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4756_y0);
  and_gate and_gate_h_u_cla24_and4757_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4757_y0);
  and_gate and_gate_h_u_cla24_and4758_y0(h_u_cla24_and4757_y0, h_u_cla24_and4756_y0, h_u_cla24_and4758_y0);
  and_gate and_gate_h_u_cla24_and4759_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4759_y0);
  and_gate and_gate_h_u_cla24_and4760_y0(h_u_cla24_and4759_y0, h_u_cla24_and4758_y0, h_u_cla24_and4760_y0);
  and_gate and_gate_h_u_cla24_and4761_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4761_y0);
  and_gate and_gate_h_u_cla24_and4762_y0(h_u_cla24_and4761_y0, h_u_cla24_and4760_y0, h_u_cla24_and4762_y0);
  and_gate and_gate_h_u_cla24_and4763_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4763_y0);
  and_gate and_gate_h_u_cla24_and4764_y0(h_u_cla24_and4763_y0, h_u_cla24_and4762_y0, h_u_cla24_and4764_y0);
  and_gate and_gate_h_u_cla24_and4765_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4765_y0);
  and_gate and_gate_h_u_cla24_and4766_y0(h_u_cla24_and4765_y0, h_u_cla24_and4764_y0, h_u_cla24_and4766_y0);
  and_gate and_gate_h_u_cla24_and4767_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4767_y0);
  and_gate and_gate_h_u_cla24_and4768_y0(h_u_cla24_and4767_y0, h_u_cla24_and4766_y0, h_u_cla24_and4768_y0);
  and_gate and_gate_h_u_cla24_and4769_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4769_y0);
  and_gate and_gate_h_u_cla24_and4770_y0(h_u_cla24_and4769_y0, h_u_cla24_and4768_y0, h_u_cla24_and4770_y0);
  and_gate and_gate_h_u_cla24_and4771_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4771_y0);
  and_gate and_gate_h_u_cla24_and4772_y0(h_u_cla24_and4771_y0, h_u_cla24_and4770_y0, h_u_cla24_and4772_y0);
  and_gate and_gate_h_u_cla24_and4773_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4773_y0);
  and_gate and_gate_h_u_cla24_and4774_y0(h_u_cla24_and4773_y0, h_u_cla24_and4772_y0, h_u_cla24_and4774_y0);
  and_gate and_gate_h_u_cla24_and4775_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4775_y0);
  and_gate and_gate_h_u_cla24_and4776_y0(h_u_cla24_and4775_y0, h_u_cla24_and4774_y0, h_u_cla24_and4776_y0);
  and_gate and_gate_h_u_cla24_and4777_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic11_y1, h_u_cla24_and4777_y0);
  and_gate and_gate_h_u_cla24_and4778_y0(h_u_cla24_and4777_y0, h_u_cla24_and4776_y0, h_u_cla24_and4778_y0);
  and_gate and_gate_h_u_cla24_and4779_y0(h_u_cla24_pg_logic13_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4779_y0);
  and_gate and_gate_h_u_cla24_and4780_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4780_y0);
  and_gate and_gate_h_u_cla24_and4781_y0(h_u_cla24_and4780_y0, h_u_cla24_and4779_y0, h_u_cla24_and4781_y0);
  and_gate and_gate_h_u_cla24_and4782_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4782_y0);
  and_gate and_gate_h_u_cla24_and4783_y0(h_u_cla24_and4782_y0, h_u_cla24_and4781_y0, h_u_cla24_and4783_y0);
  and_gate and_gate_h_u_cla24_and4784_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4784_y0);
  and_gate and_gate_h_u_cla24_and4785_y0(h_u_cla24_and4784_y0, h_u_cla24_and4783_y0, h_u_cla24_and4785_y0);
  and_gate and_gate_h_u_cla24_and4786_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4786_y0);
  and_gate and_gate_h_u_cla24_and4787_y0(h_u_cla24_and4786_y0, h_u_cla24_and4785_y0, h_u_cla24_and4787_y0);
  and_gate and_gate_h_u_cla24_and4788_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4788_y0);
  and_gate and_gate_h_u_cla24_and4789_y0(h_u_cla24_and4788_y0, h_u_cla24_and4787_y0, h_u_cla24_and4789_y0);
  and_gate and_gate_h_u_cla24_and4790_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4790_y0);
  and_gate and_gate_h_u_cla24_and4791_y0(h_u_cla24_and4790_y0, h_u_cla24_and4789_y0, h_u_cla24_and4791_y0);
  and_gate and_gate_h_u_cla24_and4792_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4792_y0);
  and_gate and_gate_h_u_cla24_and4793_y0(h_u_cla24_and4792_y0, h_u_cla24_and4791_y0, h_u_cla24_and4793_y0);
  and_gate and_gate_h_u_cla24_and4794_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4794_y0);
  and_gate and_gate_h_u_cla24_and4795_y0(h_u_cla24_and4794_y0, h_u_cla24_and4793_y0, h_u_cla24_and4795_y0);
  and_gate and_gate_h_u_cla24_and4796_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4796_y0);
  and_gate and_gate_h_u_cla24_and4797_y0(h_u_cla24_and4796_y0, h_u_cla24_and4795_y0, h_u_cla24_and4797_y0);
  and_gate and_gate_h_u_cla24_and4798_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic12_y1, h_u_cla24_and4798_y0);
  and_gate and_gate_h_u_cla24_and4799_y0(h_u_cla24_and4798_y0, h_u_cla24_and4797_y0, h_u_cla24_and4799_y0);
  and_gate and_gate_h_u_cla24_and4800_y0(h_u_cla24_pg_logic14_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4800_y0);
  and_gate and_gate_h_u_cla24_and4801_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4801_y0);
  and_gate and_gate_h_u_cla24_and4802_y0(h_u_cla24_and4801_y0, h_u_cla24_and4800_y0, h_u_cla24_and4802_y0);
  and_gate and_gate_h_u_cla24_and4803_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4803_y0);
  and_gate and_gate_h_u_cla24_and4804_y0(h_u_cla24_and4803_y0, h_u_cla24_and4802_y0, h_u_cla24_and4804_y0);
  and_gate and_gate_h_u_cla24_and4805_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4805_y0);
  and_gate and_gate_h_u_cla24_and4806_y0(h_u_cla24_and4805_y0, h_u_cla24_and4804_y0, h_u_cla24_and4806_y0);
  and_gate and_gate_h_u_cla24_and4807_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4807_y0);
  and_gate and_gate_h_u_cla24_and4808_y0(h_u_cla24_and4807_y0, h_u_cla24_and4806_y0, h_u_cla24_and4808_y0);
  and_gate and_gate_h_u_cla24_and4809_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4809_y0);
  and_gate and_gate_h_u_cla24_and4810_y0(h_u_cla24_and4809_y0, h_u_cla24_and4808_y0, h_u_cla24_and4810_y0);
  and_gate and_gate_h_u_cla24_and4811_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4811_y0);
  and_gate and_gate_h_u_cla24_and4812_y0(h_u_cla24_and4811_y0, h_u_cla24_and4810_y0, h_u_cla24_and4812_y0);
  and_gate and_gate_h_u_cla24_and4813_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4813_y0);
  and_gate and_gate_h_u_cla24_and4814_y0(h_u_cla24_and4813_y0, h_u_cla24_and4812_y0, h_u_cla24_and4814_y0);
  and_gate and_gate_h_u_cla24_and4815_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4815_y0);
  and_gate and_gate_h_u_cla24_and4816_y0(h_u_cla24_and4815_y0, h_u_cla24_and4814_y0, h_u_cla24_and4816_y0);
  and_gate and_gate_h_u_cla24_and4817_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic13_y1, h_u_cla24_and4817_y0);
  and_gate and_gate_h_u_cla24_and4818_y0(h_u_cla24_and4817_y0, h_u_cla24_and4816_y0, h_u_cla24_and4818_y0);
  and_gate and_gate_h_u_cla24_and4819_y0(h_u_cla24_pg_logic15_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4819_y0);
  and_gate and_gate_h_u_cla24_and4820_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4820_y0);
  and_gate and_gate_h_u_cla24_and4821_y0(h_u_cla24_and4820_y0, h_u_cla24_and4819_y0, h_u_cla24_and4821_y0);
  and_gate and_gate_h_u_cla24_and4822_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4822_y0);
  and_gate and_gate_h_u_cla24_and4823_y0(h_u_cla24_and4822_y0, h_u_cla24_and4821_y0, h_u_cla24_and4823_y0);
  and_gate and_gate_h_u_cla24_and4824_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4824_y0);
  and_gate and_gate_h_u_cla24_and4825_y0(h_u_cla24_and4824_y0, h_u_cla24_and4823_y0, h_u_cla24_and4825_y0);
  and_gate and_gate_h_u_cla24_and4826_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4826_y0);
  and_gate and_gate_h_u_cla24_and4827_y0(h_u_cla24_and4826_y0, h_u_cla24_and4825_y0, h_u_cla24_and4827_y0);
  and_gate and_gate_h_u_cla24_and4828_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4828_y0);
  and_gate and_gate_h_u_cla24_and4829_y0(h_u_cla24_and4828_y0, h_u_cla24_and4827_y0, h_u_cla24_and4829_y0);
  and_gate and_gate_h_u_cla24_and4830_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4830_y0);
  and_gate and_gate_h_u_cla24_and4831_y0(h_u_cla24_and4830_y0, h_u_cla24_and4829_y0, h_u_cla24_and4831_y0);
  and_gate and_gate_h_u_cla24_and4832_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4832_y0);
  and_gate and_gate_h_u_cla24_and4833_y0(h_u_cla24_and4832_y0, h_u_cla24_and4831_y0, h_u_cla24_and4833_y0);
  and_gate and_gate_h_u_cla24_and4834_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic14_y1, h_u_cla24_and4834_y0);
  and_gate and_gate_h_u_cla24_and4835_y0(h_u_cla24_and4834_y0, h_u_cla24_and4833_y0, h_u_cla24_and4835_y0);
  and_gate and_gate_h_u_cla24_and4836_y0(h_u_cla24_pg_logic16_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4836_y0);
  and_gate and_gate_h_u_cla24_and4837_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4837_y0);
  and_gate and_gate_h_u_cla24_and4838_y0(h_u_cla24_and4837_y0, h_u_cla24_and4836_y0, h_u_cla24_and4838_y0);
  and_gate and_gate_h_u_cla24_and4839_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4839_y0);
  and_gate and_gate_h_u_cla24_and4840_y0(h_u_cla24_and4839_y0, h_u_cla24_and4838_y0, h_u_cla24_and4840_y0);
  and_gate and_gate_h_u_cla24_and4841_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4841_y0);
  and_gate and_gate_h_u_cla24_and4842_y0(h_u_cla24_and4841_y0, h_u_cla24_and4840_y0, h_u_cla24_and4842_y0);
  and_gate and_gate_h_u_cla24_and4843_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4843_y0);
  and_gate and_gate_h_u_cla24_and4844_y0(h_u_cla24_and4843_y0, h_u_cla24_and4842_y0, h_u_cla24_and4844_y0);
  and_gate and_gate_h_u_cla24_and4845_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4845_y0);
  and_gate and_gate_h_u_cla24_and4846_y0(h_u_cla24_and4845_y0, h_u_cla24_and4844_y0, h_u_cla24_and4846_y0);
  and_gate and_gate_h_u_cla24_and4847_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4847_y0);
  and_gate and_gate_h_u_cla24_and4848_y0(h_u_cla24_and4847_y0, h_u_cla24_and4846_y0, h_u_cla24_and4848_y0);
  and_gate and_gate_h_u_cla24_and4849_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic15_y1, h_u_cla24_and4849_y0);
  and_gate and_gate_h_u_cla24_and4850_y0(h_u_cla24_and4849_y0, h_u_cla24_and4848_y0, h_u_cla24_and4850_y0);
  and_gate and_gate_h_u_cla24_and4851_y0(h_u_cla24_pg_logic17_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4851_y0);
  and_gate and_gate_h_u_cla24_and4852_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4852_y0);
  and_gate and_gate_h_u_cla24_and4853_y0(h_u_cla24_and4852_y0, h_u_cla24_and4851_y0, h_u_cla24_and4853_y0);
  and_gate and_gate_h_u_cla24_and4854_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4854_y0);
  and_gate and_gate_h_u_cla24_and4855_y0(h_u_cla24_and4854_y0, h_u_cla24_and4853_y0, h_u_cla24_and4855_y0);
  and_gate and_gate_h_u_cla24_and4856_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4856_y0);
  and_gate and_gate_h_u_cla24_and4857_y0(h_u_cla24_and4856_y0, h_u_cla24_and4855_y0, h_u_cla24_and4857_y0);
  and_gate and_gate_h_u_cla24_and4858_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4858_y0);
  and_gate and_gate_h_u_cla24_and4859_y0(h_u_cla24_and4858_y0, h_u_cla24_and4857_y0, h_u_cla24_and4859_y0);
  and_gate and_gate_h_u_cla24_and4860_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4860_y0);
  and_gate and_gate_h_u_cla24_and4861_y0(h_u_cla24_and4860_y0, h_u_cla24_and4859_y0, h_u_cla24_and4861_y0);
  and_gate and_gate_h_u_cla24_and4862_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic16_y1, h_u_cla24_and4862_y0);
  and_gate and_gate_h_u_cla24_and4863_y0(h_u_cla24_and4862_y0, h_u_cla24_and4861_y0, h_u_cla24_and4863_y0);
  and_gate and_gate_h_u_cla24_and4864_y0(h_u_cla24_pg_logic18_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4864_y0);
  and_gate and_gate_h_u_cla24_and4865_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4865_y0);
  and_gate and_gate_h_u_cla24_and4866_y0(h_u_cla24_and4865_y0, h_u_cla24_and4864_y0, h_u_cla24_and4866_y0);
  and_gate and_gate_h_u_cla24_and4867_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4867_y0);
  and_gate and_gate_h_u_cla24_and4868_y0(h_u_cla24_and4867_y0, h_u_cla24_and4866_y0, h_u_cla24_and4868_y0);
  and_gate and_gate_h_u_cla24_and4869_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4869_y0);
  and_gate and_gate_h_u_cla24_and4870_y0(h_u_cla24_and4869_y0, h_u_cla24_and4868_y0, h_u_cla24_and4870_y0);
  and_gate and_gate_h_u_cla24_and4871_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4871_y0);
  and_gate and_gate_h_u_cla24_and4872_y0(h_u_cla24_and4871_y0, h_u_cla24_and4870_y0, h_u_cla24_and4872_y0);
  and_gate and_gate_h_u_cla24_and4873_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic17_y1, h_u_cla24_and4873_y0);
  and_gate and_gate_h_u_cla24_and4874_y0(h_u_cla24_and4873_y0, h_u_cla24_and4872_y0, h_u_cla24_and4874_y0);
  and_gate and_gate_h_u_cla24_and4875_y0(h_u_cla24_pg_logic19_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and4875_y0);
  and_gate and_gate_h_u_cla24_and4876_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and4876_y0);
  and_gate and_gate_h_u_cla24_and4877_y0(h_u_cla24_and4876_y0, h_u_cla24_and4875_y0, h_u_cla24_and4877_y0);
  and_gate and_gate_h_u_cla24_and4878_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and4878_y0);
  and_gate and_gate_h_u_cla24_and4879_y0(h_u_cla24_and4878_y0, h_u_cla24_and4877_y0, h_u_cla24_and4879_y0);
  and_gate and_gate_h_u_cla24_and4880_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and4880_y0);
  and_gate and_gate_h_u_cla24_and4881_y0(h_u_cla24_and4880_y0, h_u_cla24_and4879_y0, h_u_cla24_and4881_y0);
  and_gate and_gate_h_u_cla24_and4882_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic18_y1, h_u_cla24_and4882_y0);
  and_gate and_gate_h_u_cla24_and4883_y0(h_u_cla24_and4882_y0, h_u_cla24_and4881_y0, h_u_cla24_and4883_y0);
  and_gate and_gate_h_u_cla24_and4884_y0(h_u_cla24_pg_logic20_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and4884_y0);
  and_gate and_gate_h_u_cla24_and4885_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and4885_y0);
  and_gate and_gate_h_u_cla24_and4886_y0(h_u_cla24_and4885_y0, h_u_cla24_and4884_y0, h_u_cla24_and4886_y0);
  and_gate and_gate_h_u_cla24_and4887_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and4887_y0);
  and_gate and_gate_h_u_cla24_and4888_y0(h_u_cla24_and4887_y0, h_u_cla24_and4886_y0, h_u_cla24_and4888_y0);
  and_gate and_gate_h_u_cla24_and4889_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic19_y1, h_u_cla24_and4889_y0);
  and_gate and_gate_h_u_cla24_and4890_y0(h_u_cla24_and4889_y0, h_u_cla24_and4888_y0, h_u_cla24_and4890_y0);
  and_gate and_gate_h_u_cla24_and4891_y0(h_u_cla24_pg_logic21_y0, h_u_cla24_pg_logic20_y1, h_u_cla24_and4891_y0);
  and_gate and_gate_h_u_cla24_and4892_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic20_y1, h_u_cla24_and4892_y0);
  and_gate and_gate_h_u_cla24_and4893_y0(h_u_cla24_and4892_y0, h_u_cla24_and4891_y0, h_u_cla24_and4893_y0);
  and_gate and_gate_h_u_cla24_and4894_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic20_y1, h_u_cla24_and4894_y0);
  and_gate and_gate_h_u_cla24_and4895_y0(h_u_cla24_and4894_y0, h_u_cla24_and4893_y0, h_u_cla24_and4895_y0);
  and_gate and_gate_h_u_cla24_and4896_y0(h_u_cla24_pg_logic22_y0, h_u_cla24_pg_logic21_y1, h_u_cla24_and4896_y0);
  and_gate and_gate_h_u_cla24_and4897_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic21_y1, h_u_cla24_and4897_y0);
  and_gate and_gate_h_u_cla24_and4898_y0(h_u_cla24_and4897_y0, h_u_cla24_and4896_y0, h_u_cla24_and4898_y0);
  and_gate and_gate_h_u_cla24_and4899_y0(h_u_cla24_pg_logic23_y0, h_u_cla24_pg_logic22_y1, h_u_cla24_and4899_y0);
  or_gate or_gate_h_u_cla24_or276_y0(h_u_cla24_and4899_y0, h_u_cla24_and4370_y0, h_u_cla24_or276_y0);
  or_gate or_gate_h_u_cla24_or277_y0(h_u_cla24_or276_y0, h_u_cla24_and4415_y0, h_u_cla24_or277_y0);
  or_gate or_gate_h_u_cla24_or278_y0(h_u_cla24_or277_y0, h_u_cla24_and4458_y0, h_u_cla24_or278_y0);
  or_gate or_gate_h_u_cla24_or279_y0(h_u_cla24_or278_y0, h_u_cla24_and4499_y0, h_u_cla24_or279_y0);
  or_gate or_gate_h_u_cla24_or280_y0(h_u_cla24_or279_y0, h_u_cla24_and4538_y0, h_u_cla24_or280_y0);
  or_gate or_gate_h_u_cla24_or281_y0(h_u_cla24_or280_y0, h_u_cla24_and4575_y0, h_u_cla24_or281_y0);
  or_gate or_gate_h_u_cla24_or282_y0(h_u_cla24_or281_y0, h_u_cla24_and4610_y0, h_u_cla24_or282_y0);
  or_gate or_gate_h_u_cla24_or283_y0(h_u_cla24_or282_y0, h_u_cla24_and4643_y0, h_u_cla24_or283_y0);
  or_gate or_gate_h_u_cla24_or284_y0(h_u_cla24_or283_y0, h_u_cla24_and4674_y0, h_u_cla24_or284_y0);
  or_gate or_gate_h_u_cla24_or285_y0(h_u_cla24_or284_y0, h_u_cla24_and4703_y0, h_u_cla24_or285_y0);
  or_gate or_gate_h_u_cla24_or286_y0(h_u_cla24_or285_y0, h_u_cla24_and4730_y0, h_u_cla24_or286_y0);
  or_gate or_gate_h_u_cla24_or287_y0(h_u_cla24_or286_y0, h_u_cla24_and4755_y0, h_u_cla24_or287_y0);
  or_gate or_gate_h_u_cla24_or288_y0(h_u_cla24_or287_y0, h_u_cla24_and4778_y0, h_u_cla24_or288_y0);
  or_gate or_gate_h_u_cla24_or289_y0(h_u_cla24_or288_y0, h_u_cla24_and4799_y0, h_u_cla24_or289_y0);
  or_gate or_gate_h_u_cla24_or290_y0(h_u_cla24_or289_y0, h_u_cla24_and4818_y0, h_u_cla24_or290_y0);
  or_gate or_gate_h_u_cla24_or291_y0(h_u_cla24_or290_y0, h_u_cla24_and4835_y0, h_u_cla24_or291_y0);
  or_gate or_gate_h_u_cla24_or292_y0(h_u_cla24_or291_y0, h_u_cla24_and4850_y0, h_u_cla24_or292_y0);
  or_gate or_gate_h_u_cla24_or293_y0(h_u_cla24_or292_y0, h_u_cla24_and4863_y0, h_u_cla24_or293_y0);
  or_gate or_gate_h_u_cla24_or294_y0(h_u_cla24_or293_y0, h_u_cla24_and4874_y0, h_u_cla24_or294_y0);
  or_gate or_gate_h_u_cla24_or295_y0(h_u_cla24_or294_y0, h_u_cla24_and4883_y0, h_u_cla24_or295_y0);
  or_gate or_gate_h_u_cla24_or296_y0(h_u_cla24_or295_y0, h_u_cla24_and4890_y0, h_u_cla24_or296_y0);
  or_gate or_gate_h_u_cla24_or297_y0(h_u_cla24_or296_y0, h_u_cla24_and4895_y0, h_u_cla24_or297_y0);
  or_gate or_gate_h_u_cla24_or298_y0(h_u_cla24_or297_y0, h_u_cla24_and4898_y0, h_u_cla24_or298_y0);
  or_gate or_gate_h_u_cla24_or299_y0(h_u_cla24_pg_logic23_y1, h_u_cla24_or298_y0, h_u_cla24_or299_y0);

  assign out[0] = h_u_cla24_xor0_y0;
  assign out[1] = h_u_cla24_xor1_y0;
  assign out[2] = h_u_cla24_xor2_y0;
  assign out[3] = h_u_cla24_xor3_y0;
  assign out[4] = h_u_cla24_xor4_y0;
  assign out[5] = h_u_cla24_xor5_y0;
  assign out[6] = h_u_cla24_xor6_y0;
  assign out[7] = h_u_cla24_xor7_y0;
  assign out[8] = h_u_cla24_xor8_y0;
  assign out[9] = h_u_cla24_xor9_y0;
  assign out[10] = h_u_cla24_xor10_y0;
  assign out[11] = h_u_cla24_xor11_y0;
  assign out[12] = h_u_cla24_xor12_y0;
  assign out[13] = h_u_cla24_xor13_y0;
  assign out[14] = h_u_cla24_xor14_y0;
  assign out[15] = h_u_cla24_xor15_y0;
  assign out[16] = h_u_cla24_xor16_y0;
  assign out[17] = h_u_cla24_xor17_y0;
  assign out[18] = h_u_cla24_xor18_y0;
  assign out[19] = h_u_cla24_xor19_y0;
  assign out[20] = h_u_cla24_xor20_y0;
  assign out[21] = h_u_cla24_xor21_y0;
  assign out[22] = h_u_cla24_xor22_y0;
  assign out[23] = h_u_cla24_xor23_y0;
  assign out[24] = h_u_cla24_or299_y0;
endmodule