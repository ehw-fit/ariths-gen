module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(a[0], b[0], pg_logic_or0);
  and_gate and_gate_pg_logic_and0(a[0], b[0], pg_logic_and0);
  xor_gate xor_gate_pg_logic_xor0(a[0], b[0], pg_logic_xor0);
endmodule

module h_s_cla32(input [31:0] a, input [31:0] b, output [32:0] h_s_cla32_out);
  wire [0:0] h_s_cla32_pg_logic0_or0;
  wire [0:0] h_s_cla32_pg_logic0_and0;
  wire [0:0] h_s_cla32_pg_logic0_xor0;
  wire [0:0] h_s_cla32_pg_logic1_or0;
  wire [0:0] h_s_cla32_pg_logic1_and0;
  wire [0:0] h_s_cla32_pg_logic1_xor0;
  wire [0:0] h_s_cla32_xor1;
  wire [0:0] h_s_cla32_and0;
  wire [0:0] h_s_cla32_or0;
  wire [0:0] h_s_cla32_pg_logic2_or0;
  wire [0:0] h_s_cla32_pg_logic2_and0;
  wire [0:0] h_s_cla32_pg_logic2_xor0;
  wire [0:0] h_s_cla32_xor2;
  wire [0:0] h_s_cla32_and1;
  wire [0:0] h_s_cla32_and2;
  wire [0:0] h_s_cla32_and3;
  wire [0:0] h_s_cla32_and4;
  wire [0:0] h_s_cla32_or1;
  wire [0:0] h_s_cla32_or2;
  wire [0:0] h_s_cla32_pg_logic3_or0;
  wire [0:0] h_s_cla32_pg_logic3_and0;
  wire [0:0] h_s_cla32_pg_logic3_xor0;
  wire [0:0] h_s_cla32_xor3;
  wire [0:0] h_s_cla32_and5;
  wire [0:0] h_s_cla32_and6;
  wire [0:0] h_s_cla32_and7;
  wire [0:0] h_s_cla32_and8;
  wire [0:0] h_s_cla32_and9;
  wire [0:0] h_s_cla32_and10;
  wire [0:0] h_s_cla32_and11;
  wire [0:0] h_s_cla32_or3;
  wire [0:0] h_s_cla32_or4;
  wire [0:0] h_s_cla32_or5;
  wire [0:0] h_s_cla32_pg_logic4_or0;
  wire [0:0] h_s_cla32_pg_logic4_and0;
  wire [0:0] h_s_cla32_pg_logic4_xor0;
  wire [0:0] h_s_cla32_xor4;
  wire [0:0] h_s_cla32_and12;
  wire [0:0] h_s_cla32_or6;
  wire [0:0] h_s_cla32_pg_logic5_or0;
  wire [0:0] h_s_cla32_pg_logic5_and0;
  wire [0:0] h_s_cla32_pg_logic5_xor0;
  wire [0:0] h_s_cla32_xor5;
  wire [0:0] h_s_cla32_and13;
  wire [0:0] h_s_cla32_and14;
  wire [0:0] h_s_cla32_and15;
  wire [0:0] h_s_cla32_or7;
  wire [0:0] h_s_cla32_or8;
  wire [0:0] h_s_cla32_pg_logic6_or0;
  wire [0:0] h_s_cla32_pg_logic6_and0;
  wire [0:0] h_s_cla32_pg_logic6_xor0;
  wire [0:0] h_s_cla32_xor6;
  wire [0:0] h_s_cla32_and16;
  wire [0:0] h_s_cla32_and17;
  wire [0:0] h_s_cla32_and18;
  wire [0:0] h_s_cla32_and19;
  wire [0:0] h_s_cla32_and20;
  wire [0:0] h_s_cla32_and21;
  wire [0:0] h_s_cla32_or9;
  wire [0:0] h_s_cla32_or10;
  wire [0:0] h_s_cla32_or11;
  wire [0:0] h_s_cla32_pg_logic7_or0;
  wire [0:0] h_s_cla32_pg_logic7_and0;
  wire [0:0] h_s_cla32_pg_logic7_xor0;
  wire [0:0] h_s_cla32_xor7;
  wire [0:0] h_s_cla32_and22;
  wire [0:0] h_s_cla32_and23;
  wire [0:0] h_s_cla32_and24;
  wire [0:0] h_s_cla32_and25;
  wire [0:0] h_s_cla32_and26;
  wire [0:0] h_s_cla32_and27;
  wire [0:0] h_s_cla32_and28;
  wire [0:0] h_s_cla32_and29;
  wire [0:0] h_s_cla32_and30;
  wire [0:0] h_s_cla32_and31;
  wire [0:0] h_s_cla32_or12;
  wire [0:0] h_s_cla32_or13;
  wire [0:0] h_s_cla32_or14;
  wire [0:0] h_s_cla32_or15;
  wire [0:0] h_s_cla32_pg_logic8_or0;
  wire [0:0] h_s_cla32_pg_logic8_and0;
  wire [0:0] h_s_cla32_pg_logic8_xor0;
  wire [0:0] h_s_cla32_xor8;
  wire [0:0] h_s_cla32_and32;
  wire [0:0] h_s_cla32_or16;
  wire [0:0] h_s_cla32_pg_logic9_or0;
  wire [0:0] h_s_cla32_pg_logic9_and0;
  wire [0:0] h_s_cla32_pg_logic9_xor0;
  wire [0:0] h_s_cla32_xor9;
  wire [0:0] h_s_cla32_and33;
  wire [0:0] h_s_cla32_and34;
  wire [0:0] h_s_cla32_and35;
  wire [0:0] h_s_cla32_or17;
  wire [0:0] h_s_cla32_or18;
  wire [0:0] h_s_cla32_pg_logic10_or0;
  wire [0:0] h_s_cla32_pg_logic10_and0;
  wire [0:0] h_s_cla32_pg_logic10_xor0;
  wire [0:0] h_s_cla32_xor10;
  wire [0:0] h_s_cla32_and36;
  wire [0:0] h_s_cla32_and37;
  wire [0:0] h_s_cla32_and38;
  wire [0:0] h_s_cla32_and39;
  wire [0:0] h_s_cla32_and40;
  wire [0:0] h_s_cla32_and41;
  wire [0:0] h_s_cla32_or19;
  wire [0:0] h_s_cla32_or20;
  wire [0:0] h_s_cla32_or21;
  wire [0:0] h_s_cla32_pg_logic11_or0;
  wire [0:0] h_s_cla32_pg_logic11_and0;
  wire [0:0] h_s_cla32_pg_logic11_xor0;
  wire [0:0] h_s_cla32_xor11;
  wire [0:0] h_s_cla32_and42;
  wire [0:0] h_s_cla32_and43;
  wire [0:0] h_s_cla32_and44;
  wire [0:0] h_s_cla32_and45;
  wire [0:0] h_s_cla32_and46;
  wire [0:0] h_s_cla32_and47;
  wire [0:0] h_s_cla32_and48;
  wire [0:0] h_s_cla32_and49;
  wire [0:0] h_s_cla32_and50;
  wire [0:0] h_s_cla32_and51;
  wire [0:0] h_s_cla32_or22;
  wire [0:0] h_s_cla32_or23;
  wire [0:0] h_s_cla32_or24;
  wire [0:0] h_s_cla32_or25;
  wire [0:0] h_s_cla32_pg_logic12_or0;
  wire [0:0] h_s_cla32_pg_logic12_and0;
  wire [0:0] h_s_cla32_pg_logic12_xor0;
  wire [0:0] h_s_cla32_xor12;
  wire [0:0] h_s_cla32_and52;
  wire [0:0] h_s_cla32_or26;
  wire [0:0] h_s_cla32_pg_logic13_or0;
  wire [0:0] h_s_cla32_pg_logic13_and0;
  wire [0:0] h_s_cla32_pg_logic13_xor0;
  wire [0:0] h_s_cla32_xor13;
  wire [0:0] h_s_cla32_and53;
  wire [0:0] h_s_cla32_and54;
  wire [0:0] h_s_cla32_and55;
  wire [0:0] h_s_cla32_or27;
  wire [0:0] h_s_cla32_or28;
  wire [0:0] h_s_cla32_pg_logic14_or0;
  wire [0:0] h_s_cla32_pg_logic14_and0;
  wire [0:0] h_s_cla32_pg_logic14_xor0;
  wire [0:0] h_s_cla32_xor14;
  wire [0:0] h_s_cla32_and56;
  wire [0:0] h_s_cla32_and57;
  wire [0:0] h_s_cla32_and58;
  wire [0:0] h_s_cla32_and59;
  wire [0:0] h_s_cla32_and60;
  wire [0:0] h_s_cla32_and61;
  wire [0:0] h_s_cla32_or29;
  wire [0:0] h_s_cla32_or30;
  wire [0:0] h_s_cla32_or31;
  wire [0:0] h_s_cla32_pg_logic15_or0;
  wire [0:0] h_s_cla32_pg_logic15_and0;
  wire [0:0] h_s_cla32_pg_logic15_xor0;
  wire [0:0] h_s_cla32_xor15;
  wire [0:0] h_s_cla32_and62;
  wire [0:0] h_s_cla32_and63;
  wire [0:0] h_s_cla32_and64;
  wire [0:0] h_s_cla32_and65;
  wire [0:0] h_s_cla32_and66;
  wire [0:0] h_s_cla32_and67;
  wire [0:0] h_s_cla32_and68;
  wire [0:0] h_s_cla32_and69;
  wire [0:0] h_s_cla32_and70;
  wire [0:0] h_s_cla32_and71;
  wire [0:0] h_s_cla32_or32;
  wire [0:0] h_s_cla32_or33;
  wire [0:0] h_s_cla32_or34;
  wire [0:0] h_s_cla32_or35;
  wire [0:0] h_s_cla32_pg_logic16_or0;
  wire [0:0] h_s_cla32_pg_logic16_and0;
  wire [0:0] h_s_cla32_pg_logic16_xor0;
  wire [0:0] h_s_cla32_xor16;
  wire [0:0] h_s_cla32_and72;
  wire [0:0] h_s_cla32_or36;
  wire [0:0] h_s_cla32_pg_logic17_or0;
  wire [0:0] h_s_cla32_pg_logic17_and0;
  wire [0:0] h_s_cla32_pg_logic17_xor0;
  wire [0:0] h_s_cla32_xor17;
  wire [0:0] h_s_cla32_and73;
  wire [0:0] h_s_cla32_and74;
  wire [0:0] h_s_cla32_and75;
  wire [0:0] h_s_cla32_or37;
  wire [0:0] h_s_cla32_or38;
  wire [0:0] h_s_cla32_pg_logic18_or0;
  wire [0:0] h_s_cla32_pg_logic18_and0;
  wire [0:0] h_s_cla32_pg_logic18_xor0;
  wire [0:0] h_s_cla32_xor18;
  wire [0:0] h_s_cla32_and76;
  wire [0:0] h_s_cla32_and77;
  wire [0:0] h_s_cla32_and78;
  wire [0:0] h_s_cla32_and79;
  wire [0:0] h_s_cla32_and80;
  wire [0:0] h_s_cla32_and81;
  wire [0:0] h_s_cla32_or39;
  wire [0:0] h_s_cla32_or40;
  wire [0:0] h_s_cla32_or41;
  wire [0:0] h_s_cla32_pg_logic19_or0;
  wire [0:0] h_s_cla32_pg_logic19_and0;
  wire [0:0] h_s_cla32_pg_logic19_xor0;
  wire [0:0] h_s_cla32_xor19;
  wire [0:0] h_s_cla32_and82;
  wire [0:0] h_s_cla32_and83;
  wire [0:0] h_s_cla32_and84;
  wire [0:0] h_s_cla32_and85;
  wire [0:0] h_s_cla32_and86;
  wire [0:0] h_s_cla32_and87;
  wire [0:0] h_s_cla32_and88;
  wire [0:0] h_s_cla32_and89;
  wire [0:0] h_s_cla32_and90;
  wire [0:0] h_s_cla32_and91;
  wire [0:0] h_s_cla32_or42;
  wire [0:0] h_s_cla32_or43;
  wire [0:0] h_s_cla32_or44;
  wire [0:0] h_s_cla32_or45;
  wire [0:0] h_s_cla32_pg_logic20_or0;
  wire [0:0] h_s_cla32_pg_logic20_and0;
  wire [0:0] h_s_cla32_pg_logic20_xor0;
  wire [0:0] h_s_cla32_xor20;
  wire [0:0] h_s_cla32_and92;
  wire [0:0] h_s_cla32_or46;
  wire [0:0] h_s_cla32_pg_logic21_or0;
  wire [0:0] h_s_cla32_pg_logic21_and0;
  wire [0:0] h_s_cla32_pg_logic21_xor0;
  wire [0:0] h_s_cla32_xor21;
  wire [0:0] h_s_cla32_and93;
  wire [0:0] h_s_cla32_and94;
  wire [0:0] h_s_cla32_and95;
  wire [0:0] h_s_cla32_or47;
  wire [0:0] h_s_cla32_or48;
  wire [0:0] h_s_cla32_pg_logic22_or0;
  wire [0:0] h_s_cla32_pg_logic22_and0;
  wire [0:0] h_s_cla32_pg_logic22_xor0;
  wire [0:0] h_s_cla32_xor22;
  wire [0:0] h_s_cla32_and96;
  wire [0:0] h_s_cla32_and97;
  wire [0:0] h_s_cla32_and98;
  wire [0:0] h_s_cla32_and99;
  wire [0:0] h_s_cla32_and100;
  wire [0:0] h_s_cla32_and101;
  wire [0:0] h_s_cla32_or49;
  wire [0:0] h_s_cla32_or50;
  wire [0:0] h_s_cla32_or51;
  wire [0:0] h_s_cla32_pg_logic23_or0;
  wire [0:0] h_s_cla32_pg_logic23_and0;
  wire [0:0] h_s_cla32_pg_logic23_xor0;
  wire [0:0] h_s_cla32_xor23;
  wire [0:0] h_s_cla32_and102;
  wire [0:0] h_s_cla32_and103;
  wire [0:0] h_s_cla32_and104;
  wire [0:0] h_s_cla32_and105;
  wire [0:0] h_s_cla32_and106;
  wire [0:0] h_s_cla32_and107;
  wire [0:0] h_s_cla32_and108;
  wire [0:0] h_s_cla32_and109;
  wire [0:0] h_s_cla32_and110;
  wire [0:0] h_s_cla32_and111;
  wire [0:0] h_s_cla32_or52;
  wire [0:0] h_s_cla32_or53;
  wire [0:0] h_s_cla32_or54;
  wire [0:0] h_s_cla32_or55;
  wire [0:0] h_s_cla32_pg_logic24_or0;
  wire [0:0] h_s_cla32_pg_logic24_and0;
  wire [0:0] h_s_cla32_pg_logic24_xor0;
  wire [0:0] h_s_cla32_xor24;
  wire [0:0] h_s_cla32_and112;
  wire [0:0] h_s_cla32_or56;
  wire [0:0] h_s_cla32_pg_logic25_or0;
  wire [0:0] h_s_cla32_pg_logic25_and0;
  wire [0:0] h_s_cla32_pg_logic25_xor0;
  wire [0:0] h_s_cla32_xor25;
  wire [0:0] h_s_cla32_and113;
  wire [0:0] h_s_cla32_and114;
  wire [0:0] h_s_cla32_and115;
  wire [0:0] h_s_cla32_or57;
  wire [0:0] h_s_cla32_or58;
  wire [0:0] h_s_cla32_pg_logic26_or0;
  wire [0:0] h_s_cla32_pg_logic26_and0;
  wire [0:0] h_s_cla32_pg_logic26_xor0;
  wire [0:0] h_s_cla32_xor26;
  wire [0:0] h_s_cla32_and116;
  wire [0:0] h_s_cla32_and117;
  wire [0:0] h_s_cla32_and118;
  wire [0:0] h_s_cla32_and119;
  wire [0:0] h_s_cla32_and120;
  wire [0:0] h_s_cla32_and121;
  wire [0:0] h_s_cla32_or59;
  wire [0:0] h_s_cla32_or60;
  wire [0:0] h_s_cla32_or61;
  wire [0:0] h_s_cla32_pg_logic27_or0;
  wire [0:0] h_s_cla32_pg_logic27_and0;
  wire [0:0] h_s_cla32_pg_logic27_xor0;
  wire [0:0] h_s_cla32_xor27;
  wire [0:0] h_s_cla32_and122;
  wire [0:0] h_s_cla32_and123;
  wire [0:0] h_s_cla32_and124;
  wire [0:0] h_s_cla32_and125;
  wire [0:0] h_s_cla32_and126;
  wire [0:0] h_s_cla32_and127;
  wire [0:0] h_s_cla32_and128;
  wire [0:0] h_s_cla32_and129;
  wire [0:0] h_s_cla32_and130;
  wire [0:0] h_s_cla32_and131;
  wire [0:0] h_s_cla32_or62;
  wire [0:0] h_s_cla32_or63;
  wire [0:0] h_s_cla32_or64;
  wire [0:0] h_s_cla32_or65;
  wire [0:0] h_s_cla32_pg_logic28_or0;
  wire [0:0] h_s_cla32_pg_logic28_and0;
  wire [0:0] h_s_cla32_pg_logic28_xor0;
  wire [0:0] h_s_cla32_xor28;
  wire [0:0] h_s_cla32_and132;
  wire [0:0] h_s_cla32_or66;
  wire [0:0] h_s_cla32_pg_logic29_or0;
  wire [0:0] h_s_cla32_pg_logic29_and0;
  wire [0:0] h_s_cla32_pg_logic29_xor0;
  wire [0:0] h_s_cla32_xor29;
  wire [0:0] h_s_cla32_and133;
  wire [0:0] h_s_cla32_and134;
  wire [0:0] h_s_cla32_and135;
  wire [0:0] h_s_cla32_or67;
  wire [0:0] h_s_cla32_or68;
  wire [0:0] h_s_cla32_pg_logic30_or0;
  wire [0:0] h_s_cla32_pg_logic30_and0;
  wire [0:0] h_s_cla32_pg_logic30_xor0;
  wire [0:0] h_s_cla32_xor30;
  wire [0:0] h_s_cla32_and136;
  wire [0:0] h_s_cla32_and137;
  wire [0:0] h_s_cla32_and138;
  wire [0:0] h_s_cla32_and139;
  wire [0:0] h_s_cla32_and140;
  wire [0:0] h_s_cla32_and141;
  wire [0:0] h_s_cla32_or69;
  wire [0:0] h_s_cla32_or70;
  wire [0:0] h_s_cla32_or71;
  wire [0:0] h_s_cla32_pg_logic31_or0;
  wire [0:0] h_s_cla32_pg_logic31_and0;
  wire [0:0] h_s_cla32_pg_logic31_xor0;
  wire [0:0] h_s_cla32_xor31;
  wire [0:0] h_s_cla32_and142;
  wire [0:0] h_s_cla32_and143;
  wire [0:0] h_s_cla32_and144;
  wire [0:0] h_s_cla32_and145;
  wire [0:0] h_s_cla32_and146;
  wire [0:0] h_s_cla32_and147;
  wire [0:0] h_s_cla32_and148;
  wire [0:0] h_s_cla32_and149;
  wire [0:0] h_s_cla32_and150;
  wire [0:0] h_s_cla32_and151;
  wire [0:0] h_s_cla32_or72;
  wire [0:0] h_s_cla32_or73;
  wire [0:0] h_s_cla32_or74;
  wire [0:0] h_s_cla32_or75;
  wire [0:0] h_s_cla32_xor32;
  wire [0:0] h_s_cla32_xor33;

  pg_logic pg_logic_h_s_cla32_pg_logic0_out(a[0], b[0], h_s_cla32_pg_logic0_or0, h_s_cla32_pg_logic0_and0, h_s_cla32_pg_logic0_xor0);
  pg_logic pg_logic_h_s_cla32_pg_logic1_out(a[1], b[1], h_s_cla32_pg_logic1_or0, h_s_cla32_pg_logic1_and0, h_s_cla32_pg_logic1_xor0);
  xor_gate xor_gate_h_s_cla32_xor1(h_s_cla32_pg_logic1_xor0[0], h_s_cla32_pg_logic0_and0[0], h_s_cla32_xor1);
  and_gate and_gate_h_s_cla32_and0(h_s_cla32_pg_logic0_and0[0], h_s_cla32_pg_logic1_or0[0], h_s_cla32_and0);
  or_gate or_gate_h_s_cla32_or0(h_s_cla32_pg_logic1_and0[0], h_s_cla32_and0[0], h_s_cla32_or0);
  pg_logic pg_logic_h_s_cla32_pg_logic2_out(a[2], b[2], h_s_cla32_pg_logic2_or0, h_s_cla32_pg_logic2_and0, h_s_cla32_pg_logic2_xor0);
  xor_gate xor_gate_h_s_cla32_xor2(h_s_cla32_pg_logic2_xor0[0], h_s_cla32_or0[0], h_s_cla32_xor2);
  and_gate and_gate_h_s_cla32_and1(h_s_cla32_pg_logic2_or0[0], h_s_cla32_pg_logic0_or0[0], h_s_cla32_and1);
  and_gate and_gate_h_s_cla32_and2(h_s_cla32_pg_logic0_and0[0], h_s_cla32_pg_logic2_or0[0], h_s_cla32_and2);
  and_gate and_gate_h_s_cla32_and3(h_s_cla32_and2[0], h_s_cla32_pg_logic1_or0[0], h_s_cla32_and3);
  and_gate and_gate_h_s_cla32_and4(h_s_cla32_pg_logic1_and0[0], h_s_cla32_pg_logic2_or0[0], h_s_cla32_and4);
  or_gate or_gate_h_s_cla32_or1(h_s_cla32_and3[0], h_s_cla32_and4[0], h_s_cla32_or1);
  or_gate or_gate_h_s_cla32_or2(h_s_cla32_pg_logic2_and0[0], h_s_cla32_or1[0], h_s_cla32_or2);
  pg_logic pg_logic_h_s_cla32_pg_logic3_out(a[3], b[3], h_s_cla32_pg_logic3_or0, h_s_cla32_pg_logic3_and0, h_s_cla32_pg_logic3_xor0);
  xor_gate xor_gate_h_s_cla32_xor3(h_s_cla32_pg_logic3_xor0[0], h_s_cla32_or2[0], h_s_cla32_xor3);
  and_gate and_gate_h_s_cla32_and5(h_s_cla32_pg_logic3_or0[0], h_s_cla32_pg_logic1_or0[0], h_s_cla32_and5);
  and_gate and_gate_h_s_cla32_and6(h_s_cla32_pg_logic0_and0[0], h_s_cla32_pg_logic2_or0[0], h_s_cla32_and6);
  and_gate and_gate_h_s_cla32_and7(h_s_cla32_pg_logic3_or0[0], h_s_cla32_pg_logic1_or0[0], h_s_cla32_and7);
  and_gate and_gate_h_s_cla32_and8(h_s_cla32_and6[0], h_s_cla32_and7[0], h_s_cla32_and8);
  and_gate and_gate_h_s_cla32_and9(h_s_cla32_pg_logic1_and0[0], h_s_cla32_pg_logic3_or0[0], h_s_cla32_and9);
  and_gate and_gate_h_s_cla32_and10(h_s_cla32_and9[0], h_s_cla32_pg_logic2_or0[0], h_s_cla32_and10);
  and_gate and_gate_h_s_cla32_and11(h_s_cla32_pg_logic2_and0[0], h_s_cla32_pg_logic3_or0[0], h_s_cla32_and11);
  or_gate or_gate_h_s_cla32_or3(h_s_cla32_and8[0], h_s_cla32_and11[0], h_s_cla32_or3);
  or_gate or_gate_h_s_cla32_or4(h_s_cla32_and10[0], h_s_cla32_or3[0], h_s_cla32_or4);
  or_gate or_gate_h_s_cla32_or5(h_s_cla32_pg_logic3_and0[0], h_s_cla32_or4[0], h_s_cla32_or5);
  pg_logic pg_logic_h_s_cla32_pg_logic4_out(a[4], b[4], h_s_cla32_pg_logic4_or0, h_s_cla32_pg_logic4_and0, h_s_cla32_pg_logic4_xor0);
  xor_gate xor_gate_h_s_cla32_xor4(h_s_cla32_pg_logic4_xor0[0], h_s_cla32_or5[0], h_s_cla32_xor4);
  and_gate and_gate_h_s_cla32_and12(h_s_cla32_or5[0], h_s_cla32_pg_logic4_or0[0], h_s_cla32_and12);
  or_gate or_gate_h_s_cla32_or6(h_s_cla32_pg_logic4_and0[0], h_s_cla32_and12[0], h_s_cla32_or6);
  pg_logic pg_logic_h_s_cla32_pg_logic5_out(a[5], b[5], h_s_cla32_pg_logic5_or0, h_s_cla32_pg_logic5_and0, h_s_cla32_pg_logic5_xor0);
  xor_gate xor_gate_h_s_cla32_xor5(h_s_cla32_pg_logic5_xor0[0], h_s_cla32_or6[0], h_s_cla32_xor5);
  and_gate and_gate_h_s_cla32_and13(h_s_cla32_or5[0], h_s_cla32_pg_logic5_or0[0], h_s_cla32_and13);
  and_gate and_gate_h_s_cla32_and14(h_s_cla32_and13[0], h_s_cla32_pg_logic4_or0[0], h_s_cla32_and14);
  and_gate and_gate_h_s_cla32_and15(h_s_cla32_pg_logic4_and0[0], h_s_cla32_pg_logic5_or0[0], h_s_cla32_and15);
  or_gate or_gate_h_s_cla32_or7(h_s_cla32_and14[0], h_s_cla32_and15[0], h_s_cla32_or7);
  or_gate or_gate_h_s_cla32_or8(h_s_cla32_pg_logic5_and0[0], h_s_cla32_or7[0], h_s_cla32_or8);
  pg_logic pg_logic_h_s_cla32_pg_logic6_out(a[6], b[6], h_s_cla32_pg_logic6_or0, h_s_cla32_pg_logic6_and0, h_s_cla32_pg_logic6_xor0);
  xor_gate xor_gate_h_s_cla32_xor6(h_s_cla32_pg_logic6_xor0[0], h_s_cla32_or8[0], h_s_cla32_xor6);
  and_gate and_gate_h_s_cla32_and16(h_s_cla32_or5[0], h_s_cla32_pg_logic5_or0[0], h_s_cla32_and16);
  and_gate and_gate_h_s_cla32_and17(h_s_cla32_pg_logic6_or0[0], h_s_cla32_pg_logic4_or0[0], h_s_cla32_and17);
  and_gate and_gate_h_s_cla32_and18(h_s_cla32_and16[0], h_s_cla32_and17[0], h_s_cla32_and18);
  and_gate and_gate_h_s_cla32_and19(h_s_cla32_pg_logic4_and0[0], h_s_cla32_pg_logic6_or0[0], h_s_cla32_and19);
  and_gate and_gate_h_s_cla32_and20(h_s_cla32_and19[0], h_s_cla32_pg_logic5_or0[0], h_s_cla32_and20);
  and_gate and_gate_h_s_cla32_and21(h_s_cla32_pg_logic5_and0[0], h_s_cla32_pg_logic6_or0[0], h_s_cla32_and21);
  or_gate or_gate_h_s_cla32_or9(h_s_cla32_and18[0], h_s_cla32_and20[0], h_s_cla32_or9);
  or_gate or_gate_h_s_cla32_or10(h_s_cla32_or9[0], h_s_cla32_and21[0], h_s_cla32_or10);
  or_gate or_gate_h_s_cla32_or11(h_s_cla32_pg_logic6_and0[0], h_s_cla32_or10[0], h_s_cla32_or11);
  pg_logic pg_logic_h_s_cla32_pg_logic7_out(a[7], b[7], h_s_cla32_pg_logic7_or0, h_s_cla32_pg_logic7_and0, h_s_cla32_pg_logic7_xor0);
  xor_gate xor_gate_h_s_cla32_xor7(h_s_cla32_pg_logic7_xor0[0], h_s_cla32_or11[0], h_s_cla32_xor7);
  and_gate and_gate_h_s_cla32_and22(h_s_cla32_or5[0], h_s_cla32_pg_logic6_or0[0], h_s_cla32_and22);
  and_gate and_gate_h_s_cla32_and23(h_s_cla32_pg_logic7_or0[0], h_s_cla32_pg_logic5_or0[0], h_s_cla32_and23);
  and_gate and_gate_h_s_cla32_and24(h_s_cla32_and22[0], h_s_cla32_and23[0], h_s_cla32_and24);
  and_gate and_gate_h_s_cla32_and25(h_s_cla32_and24[0], h_s_cla32_pg_logic4_or0[0], h_s_cla32_and25);
  and_gate and_gate_h_s_cla32_and26(h_s_cla32_pg_logic4_and0[0], h_s_cla32_pg_logic6_or0[0], h_s_cla32_and26);
  and_gate and_gate_h_s_cla32_and27(h_s_cla32_pg_logic7_or0[0], h_s_cla32_pg_logic5_or0[0], h_s_cla32_and27);
  and_gate and_gate_h_s_cla32_and28(h_s_cla32_and26[0], h_s_cla32_and27[0], h_s_cla32_and28);
  and_gate and_gate_h_s_cla32_and29(h_s_cla32_pg_logic5_and0[0], h_s_cla32_pg_logic7_or0[0], h_s_cla32_and29);
  and_gate and_gate_h_s_cla32_and30(h_s_cla32_and29[0], h_s_cla32_pg_logic6_or0[0], h_s_cla32_and30);
  and_gate and_gate_h_s_cla32_and31(h_s_cla32_pg_logic6_and0[0], h_s_cla32_pg_logic7_or0[0], h_s_cla32_and31);
  or_gate or_gate_h_s_cla32_or12(h_s_cla32_and25[0], h_s_cla32_and30[0], h_s_cla32_or12);
  or_gate or_gate_h_s_cla32_or13(h_s_cla32_and28[0], h_s_cla32_and31[0], h_s_cla32_or13);
  or_gate or_gate_h_s_cla32_or14(h_s_cla32_or12[0], h_s_cla32_or13[0], h_s_cla32_or14);
  or_gate or_gate_h_s_cla32_or15(h_s_cla32_pg_logic7_and0[0], h_s_cla32_or14[0], h_s_cla32_or15);
  pg_logic pg_logic_h_s_cla32_pg_logic8_out(a[8], b[8], h_s_cla32_pg_logic8_or0, h_s_cla32_pg_logic8_and0, h_s_cla32_pg_logic8_xor0);
  xor_gate xor_gate_h_s_cla32_xor8(h_s_cla32_pg_logic8_xor0[0], h_s_cla32_or15[0], h_s_cla32_xor8);
  and_gate and_gate_h_s_cla32_and32(h_s_cla32_or15[0], h_s_cla32_pg_logic8_or0[0], h_s_cla32_and32);
  or_gate or_gate_h_s_cla32_or16(h_s_cla32_pg_logic8_and0[0], h_s_cla32_and32[0], h_s_cla32_or16);
  pg_logic pg_logic_h_s_cla32_pg_logic9_out(a[9], b[9], h_s_cla32_pg_logic9_or0, h_s_cla32_pg_logic9_and0, h_s_cla32_pg_logic9_xor0);
  xor_gate xor_gate_h_s_cla32_xor9(h_s_cla32_pg_logic9_xor0[0], h_s_cla32_or16[0], h_s_cla32_xor9);
  and_gate and_gate_h_s_cla32_and33(h_s_cla32_or15[0], h_s_cla32_pg_logic9_or0[0], h_s_cla32_and33);
  and_gate and_gate_h_s_cla32_and34(h_s_cla32_and33[0], h_s_cla32_pg_logic8_or0[0], h_s_cla32_and34);
  and_gate and_gate_h_s_cla32_and35(h_s_cla32_pg_logic8_and0[0], h_s_cla32_pg_logic9_or0[0], h_s_cla32_and35);
  or_gate or_gate_h_s_cla32_or17(h_s_cla32_and34[0], h_s_cla32_and35[0], h_s_cla32_or17);
  or_gate or_gate_h_s_cla32_or18(h_s_cla32_pg_logic9_and0[0], h_s_cla32_or17[0], h_s_cla32_or18);
  pg_logic pg_logic_h_s_cla32_pg_logic10_out(a[10], b[10], h_s_cla32_pg_logic10_or0, h_s_cla32_pg_logic10_and0, h_s_cla32_pg_logic10_xor0);
  xor_gate xor_gate_h_s_cla32_xor10(h_s_cla32_pg_logic10_xor0[0], h_s_cla32_or18[0], h_s_cla32_xor10);
  and_gate and_gate_h_s_cla32_and36(h_s_cla32_or15[0], h_s_cla32_pg_logic9_or0[0], h_s_cla32_and36);
  and_gate and_gate_h_s_cla32_and37(h_s_cla32_pg_logic10_or0[0], h_s_cla32_pg_logic8_or0[0], h_s_cla32_and37);
  and_gate and_gate_h_s_cla32_and38(h_s_cla32_and36[0], h_s_cla32_and37[0], h_s_cla32_and38);
  and_gate and_gate_h_s_cla32_and39(h_s_cla32_pg_logic8_and0[0], h_s_cla32_pg_logic10_or0[0], h_s_cla32_and39);
  and_gate and_gate_h_s_cla32_and40(h_s_cla32_and39[0], h_s_cla32_pg_logic9_or0[0], h_s_cla32_and40);
  and_gate and_gate_h_s_cla32_and41(h_s_cla32_pg_logic9_and0[0], h_s_cla32_pg_logic10_or0[0], h_s_cla32_and41);
  or_gate or_gate_h_s_cla32_or19(h_s_cla32_and38[0], h_s_cla32_and40[0], h_s_cla32_or19);
  or_gate or_gate_h_s_cla32_or20(h_s_cla32_or19[0], h_s_cla32_and41[0], h_s_cla32_or20);
  or_gate or_gate_h_s_cla32_or21(h_s_cla32_pg_logic10_and0[0], h_s_cla32_or20[0], h_s_cla32_or21);
  pg_logic pg_logic_h_s_cla32_pg_logic11_out(a[11], b[11], h_s_cla32_pg_logic11_or0, h_s_cla32_pg_logic11_and0, h_s_cla32_pg_logic11_xor0);
  xor_gate xor_gate_h_s_cla32_xor11(h_s_cla32_pg_logic11_xor0[0], h_s_cla32_or21[0], h_s_cla32_xor11);
  and_gate and_gate_h_s_cla32_and42(h_s_cla32_or15[0], h_s_cla32_pg_logic10_or0[0], h_s_cla32_and42);
  and_gate and_gate_h_s_cla32_and43(h_s_cla32_pg_logic11_or0[0], h_s_cla32_pg_logic9_or0[0], h_s_cla32_and43);
  and_gate and_gate_h_s_cla32_and44(h_s_cla32_and42[0], h_s_cla32_and43[0], h_s_cla32_and44);
  and_gate and_gate_h_s_cla32_and45(h_s_cla32_and44[0], h_s_cla32_pg_logic8_or0[0], h_s_cla32_and45);
  and_gate and_gate_h_s_cla32_and46(h_s_cla32_pg_logic8_and0[0], h_s_cla32_pg_logic10_or0[0], h_s_cla32_and46);
  and_gate and_gate_h_s_cla32_and47(h_s_cla32_pg_logic11_or0[0], h_s_cla32_pg_logic9_or0[0], h_s_cla32_and47);
  and_gate and_gate_h_s_cla32_and48(h_s_cla32_and46[0], h_s_cla32_and47[0], h_s_cla32_and48);
  and_gate and_gate_h_s_cla32_and49(h_s_cla32_pg_logic9_and0[0], h_s_cla32_pg_logic11_or0[0], h_s_cla32_and49);
  and_gate and_gate_h_s_cla32_and50(h_s_cla32_and49[0], h_s_cla32_pg_logic10_or0[0], h_s_cla32_and50);
  and_gate and_gate_h_s_cla32_and51(h_s_cla32_pg_logic10_and0[0], h_s_cla32_pg_logic11_or0[0], h_s_cla32_and51);
  or_gate or_gate_h_s_cla32_or22(h_s_cla32_and45[0], h_s_cla32_and50[0], h_s_cla32_or22);
  or_gate or_gate_h_s_cla32_or23(h_s_cla32_and48[0], h_s_cla32_and51[0], h_s_cla32_or23);
  or_gate or_gate_h_s_cla32_or24(h_s_cla32_or22[0], h_s_cla32_or23[0], h_s_cla32_or24);
  or_gate or_gate_h_s_cla32_or25(h_s_cla32_pg_logic11_and0[0], h_s_cla32_or24[0], h_s_cla32_or25);
  pg_logic pg_logic_h_s_cla32_pg_logic12_out(a[12], b[12], h_s_cla32_pg_logic12_or0, h_s_cla32_pg_logic12_and0, h_s_cla32_pg_logic12_xor0);
  xor_gate xor_gate_h_s_cla32_xor12(h_s_cla32_pg_logic12_xor0[0], h_s_cla32_or25[0], h_s_cla32_xor12);
  and_gate and_gate_h_s_cla32_and52(h_s_cla32_or25[0], h_s_cla32_pg_logic12_or0[0], h_s_cla32_and52);
  or_gate or_gate_h_s_cla32_or26(h_s_cla32_pg_logic12_and0[0], h_s_cla32_and52[0], h_s_cla32_or26);
  pg_logic pg_logic_h_s_cla32_pg_logic13_out(a[13], b[13], h_s_cla32_pg_logic13_or0, h_s_cla32_pg_logic13_and0, h_s_cla32_pg_logic13_xor0);
  xor_gate xor_gate_h_s_cla32_xor13(h_s_cla32_pg_logic13_xor0[0], h_s_cla32_or26[0], h_s_cla32_xor13);
  and_gate and_gate_h_s_cla32_and53(h_s_cla32_or25[0], h_s_cla32_pg_logic13_or0[0], h_s_cla32_and53);
  and_gate and_gate_h_s_cla32_and54(h_s_cla32_and53[0], h_s_cla32_pg_logic12_or0[0], h_s_cla32_and54);
  and_gate and_gate_h_s_cla32_and55(h_s_cla32_pg_logic12_and0[0], h_s_cla32_pg_logic13_or0[0], h_s_cla32_and55);
  or_gate or_gate_h_s_cla32_or27(h_s_cla32_and54[0], h_s_cla32_and55[0], h_s_cla32_or27);
  or_gate or_gate_h_s_cla32_or28(h_s_cla32_pg_logic13_and0[0], h_s_cla32_or27[0], h_s_cla32_or28);
  pg_logic pg_logic_h_s_cla32_pg_logic14_out(a[14], b[14], h_s_cla32_pg_logic14_or0, h_s_cla32_pg_logic14_and0, h_s_cla32_pg_logic14_xor0);
  xor_gate xor_gate_h_s_cla32_xor14(h_s_cla32_pg_logic14_xor0[0], h_s_cla32_or28[0], h_s_cla32_xor14);
  and_gate and_gate_h_s_cla32_and56(h_s_cla32_or25[0], h_s_cla32_pg_logic13_or0[0], h_s_cla32_and56);
  and_gate and_gate_h_s_cla32_and57(h_s_cla32_pg_logic14_or0[0], h_s_cla32_pg_logic12_or0[0], h_s_cla32_and57);
  and_gate and_gate_h_s_cla32_and58(h_s_cla32_and56[0], h_s_cla32_and57[0], h_s_cla32_and58);
  and_gate and_gate_h_s_cla32_and59(h_s_cla32_pg_logic12_and0[0], h_s_cla32_pg_logic14_or0[0], h_s_cla32_and59);
  and_gate and_gate_h_s_cla32_and60(h_s_cla32_and59[0], h_s_cla32_pg_logic13_or0[0], h_s_cla32_and60);
  and_gate and_gate_h_s_cla32_and61(h_s_cla32_pg_logic13_and0[0], h_s_cla32_pg_logic14_or0[0], h_s_cla32_and61);
  or_gate or_gate_h_s_cla32_or29(h_s_cla32_and58[0], h_s_cla32_and60[0], h_s_cla32_or29);
  or_gate or_gate_h_s_cla32_or30(h_s_cla32_or29[0], h_s_cla32_and61[0], h_s_cla32_or30);
  or_gate or_gate_h_s_cla32_or31(h_s_cla32_pg_logic14_and0[0], h_s_cla32_or30[0], h_s_cla32_or31);
  pg_logic pg_logic_h_s_cla32_pg_logic15_out(a[15], b[15], h_s_cla32_pg_logic15_or0, h_s_cla32_pg_logic15_and0, h_s_cla32_pg_logic15_xor0);
  xor_gate xor_gate_h_s_cla32_xor15(h_s_cla32_pg_logic15_xor0[0], h_s_cla32_or31[0], h_s_cla32_xor15);
  and_gate and_gate_h_s_cla32_and62(h_s_cla32_or25[0], h_s_cla32_pg_logic14_or0[0], h_s_cla32_and62);
  and_gate and_gate_h_s_cla32_and63(h_s_cla32_pg_logic15_or0[0], h_s_cla32_pg_logic13_or0[0], h_s_cla32_and63);
  and_gate and_gate_h_s_cla32_and64(h_s_cla32_and62[0], h_s_cla32_and63[0], h_s_cla32_and64);
  and_gate and_gate_h_s_cla32_and65(h_s_cla32_and64[0], h_s_cla32_pg_logic12_or0[0], h_s_cla32_and65);
  and_gate and_gate_h_s_cla32_and66(h_s_cla32_pg_logic12_and0[0], h_s_cla32_pg_logic14_or0[0], h_s_cla32_and66);
  and_gate and_gate_h_s_cla32_and67(h_s_cla32_pg_logic15_or0[0], h_s_cla32_pg_logic13_or0[0], h_s_cla32_and67);
  and_gate and_gate_h_s_cla32_and68(h_s_cla32_and66[0], h_s_cla32_and67[0], h_s_cla32_and68);
  and_gate and_gate_h_s_cla32_and69(h_s_cla32_pg_logic13_and0[0], h_s_cla32_pg_logic15_or0[0], h_s_cla32_and69);
  and_gate and_gate_h_s_cla32_and70(h_s_cla32_and69[0], h_s_cla32_pg_logic14_or0[0], h_s_cla32_and70);
  and_gate and_gate_h_s_cla32_and71(h_s_cla32_pg_logic14_and0[0], h_s_cla32_pg_logic15_or0[0], h_s_cla32_and71);
  or_gate or_gate_h_s_cla32_or32(h_s_cla32_and65[0], h_s_cla32_and70[0], h_s_cla32_or32);
  or_gate or_gate_h_s_cla32_or33(h_s_cla32_and68[0], h_s_cla32_and71[0], h_s_cla32_or33);
  or_gate or_gate_h_s_cla32_or34(h_s_cla32_or32[0], h_s_cla32_or33[0], h_s_cla32_or34);
  or_gate or_gate_h_s_cla32_or35(h_s_cla32_pg_logic15_and0[0], h_s_cla32_or34[0], h_s_cla32_or35);
  pg_logic pg_logic_h_s_cla32_pg_logic16_out(a[16], b[16], h_s_cla32_pg_logic16_or0, h_s_cla32_pg_logic16_and0, h_s_cla32_pg_logic16_xor0);
  xor_gate xor_gate_h_s_cla32_xor16(h_s_cla32_pg_logic16_xor0[0], h_s_cla32_or35[0], h_s_cla32_xor16);
  and_gate and_gate_h_s_cla32_and72(h_s_cla32_or35[0], h_s_cla32_pg_logic16_or0[0], h_s_cla32_and72);
  or_gate or_gate_h_s_cla32_or36(h_s_cla32_pg_logic16_and0[0], h_s_cla32_and72[0], h_s_cla32_or36);
  pg_logic pg_logic_h_s_cla32_pg_logic17_out(a[17], b[17], h_s_cla32_pg_logic17_or0, h_s_cla32_pg_logic17_and0, h_s_cla32_pg_logic17_xor0);
  xor_gate xor_gate_h_s_cla32_xor17(h_s_cla32_pg_logic17_xor0[0], h_s_cla32_or36[0], h_s_cla32_xor17);
  and_gate and_gate_h_s_cla32_and73(h_s_cla32_or35[0], h_s_cla32_pg_logic17_or0[0], h_s_cla32_and73);
  and_gate and_gate_h_s_cla32_and74(h_s_cla32_and73[0], h_s_cla32_pg_logic16_or0[0], h_s_cla32_and74);
  and_gate and_gate_h_s_cla32_and75(h_s_cla32_pg_logic16_and0[0], h_s_cla32_pg_logic17_or0[0], h_s_cla32_and75);
  or_gate or_gate_h_s_cla32_or37(h_s_cla32_and74[0], h_s_cla32_and75[0], h_s_cla32_or37);
  or_gate or_gate_h_s_cla32_or38(h_s_cla32_pg_logic17_and0[0], h_s_cla32_or37[0], h_s_cla32_or38);
  pg_logic pg_logic_h_s_cla32_pg_logic18_out(a[18], b[18], h_s_cla32_pg_logic18_or0, h_s_cla32_pg_logic18_and0, h_s_cla32_pg_logic18_xor0);
  xor_gate xor_gate_h_s_cla32_xor18(h_s_cla32_pg_logic18_xor0[0], h_s_cla32_or38[0], h_s_cla32_xor18);
  and_gate and_gate_h_s_cla32_and76(h_s_cla32_or35[0], h_s_cla32_pg_logic17_or0[0], h_s_cla32_and76);
  and_gate and_gate_h_s_cla32_and77(h_s_cla32_pg_logic18_or0[0], h_s_cla32_pg_logic16_or0[0], h_s_cla32_and77);
  and_gate and_gate_h_s_cla32_and78(h_s_cla32_and76[0], h_s_cla32_and77[0], h_s_cla32_and78);
  and_gate and_gate_h_s_cla32_and79(h_s_cla32_pg_logic16_and0[0], h_s_cla32_pg_logic18_or0[0], h_s_cla32_and79);
  and_gate and_gate_h_s_cla32_and80(h_s_cla32_and79[0], h_s_cla32_pg_logic17_or0[0], h_s_cla32_and80);
  and_gate and_gate_h_s_cla32_and81(h_s_cla32_pg_logic17_and0[0], h_s_cla32_pg_logic18_or0[0], h_s_cla32_and81);
  or_gate or_gate_h_s_cla32_or39(h_s_cla32_and78[0], h_s_cla32_and80[0], h_s_cla32_or39);
  or_gate or_gate_h_s_cla32_or40(h_s_cla32_or39[0], h_s_cla32_and81[0], h_s_cla32_or40);
  or_gate or_gate_h_s_cla32_or41(h_s_cla32_pg_logic18_and0[0], h_s_cla32_or40[0], h_s_cla32_or41);
  pg_logic pg_logic_h_s_cla32_pg_logic19_out(a[19], b[19], h_s_cla32_pg_logic19_or0, h_s_cla32_pg_logic19_and0, h_s_cla32_pg_logic19_xor0);
  xor_gate xor_gate_h_s_cla32_xor19(h_s_cla32_pg_logic19_xor0[0], h_s_cla32_or41[0], h_s_cla32_xor19);
  and_gate and_gate_h_s_cla32_and82(h_s_cla32_or35[0], h_s_cla32_pg_logic18_or0[0], h_s_cla32_and82);
  and_gate and_gate_h_s_cla32_and83(h_s_cla32_pg_logic19_or0[0], h_s_cla32_pg_logic17_or0[0], h_s_cla32_and83);
  and_gate and_gate_h_s_cla32_and84(h_s_cla32_and82[0], h_s_cla32_and83[0], h_s_cla32_and84);
  and_gate and_gate_h_s_cla32_and85(h_s_cla32_and84[0], h_s_cla32_pg_logic16_or0[0], h_s_cla32_and85);
  and_gate and_gate_h_s_cla32_and86(h_s_cla32_pg_logic16_and0[0], h_s_cla32_pg_logic18_or0[0], h_s_cla32_and86);
  and_gate and_gate_h_s_cla32_and87(h_s_cla32_pg_logic19_or0[0], h_s_cla32_pg_logic17_or0[0], h_s_cla32_and87);
  and_gate and_gate_h_s_cla32_and88(h_s_cla32_and86[0], h_s_cla32_and87[0], h_s_cla32_and88);
  and_gate and_gate_h_s_cla32_and89(h_s_cla32_pg_logic17_and0[0], h_s_cla32_pg_logic19_or0[0], h_s_cla32_and89);
  and_gate and_gate_h_s_cla32_and90(h_s_cla32_and89[0], h_s_cla32_pg_logic18_or0[0], h_s_cla32_and90);
  and_gate and_gate_h_s_cla32_and91(h_s_cla32_pg_logic18_and0[0], h_s_cla32_pg_logic19_or0[0], h_s_cla32_and91);
  or_gate or_gate_h_s_cla32_or42(h_s_cla32_and85[0], h_s_cla32_and90[0], h_s_cla32_or42);
  or_gate or_gate_h_s_cla32_or43(h_s_cla32_and88[0], h_s_cla32_and91[0], h_s_cla32_or43);
  or_gate or_gate_h_s_cla32_or44(h_s_cla32_or42[0], h_s_cla32_or43[0], h_s_cla32_or44);
  or_gate or_gate_h_s_cla32_or45(h_s_cla32_pg_logic19_and0[0], h_s_cla32_or44[0], h_s_cla32_or45);
  pg_logic pg_logic_h_s_cla32_pg_logic20_out(a[20], b[20], h_s_cla32_pg_logic20_or0, h_s_cla32_pg_logic20_and0, h_s_cla32_pg_logic20_xor0);
  xor_gate xor_gate_h_s_cla32_xor20(h_s_cla32_pg_logic20_xor0[0], h_s_cla32_or45[0], h_s_cla32_xor20);
  and_gate and_gate_h_s_cla32_and92(h_s_cla32_or45[0], h_s_cla32_pg_logic20_or0[0], h_s_cla32_and92);
  or_gate or_gate_h_s_cla32_or46(h_s_cla32_pg_logic20_and0[0], h_s_cla32_and92[0], h_s_cla32_or46);
  pg_logic pg_logic_h_s_cla32_pg_logic21_out(a[21], b[21], h_s_cla32_pg_logic21_or0, h_s_cla32_pg_logic21_and0, h_s_cla32_pg_logic21_xor0);
  xor_gate xor_gate_h_s_cla32_xor21(h_s_cla32_pg_logic21_xor0[0], h_s_cla32_or46[0], h_s_cla32_xor21);
  and_gate and_gate_h_s_cla32_and93(h_s_cla32_or45[0], h_s_cla32_pg_logic21_or0[0], h_s_cla32_and93);
  and_gate and_gate_h_s_cla32_and94(h_s_cla32_and93[0], h_s_cla32_pg_logic20_or0[0], h_s_cla32_and94);
  and_gate and_gate_h_s_cla32_and95(h_s_cla32_pg_logic20_and0[0], h_s_cla32_pg_logic21_or0[0], h_s_cla32_and95);
  or_gate or_gate_h_s_cla32_or47(h_s_cla32_and94[0], h_s_cla32_and95[0], h_s_cla32_or47);
  or_gate or_gate_h_s_cla32_or48(h_s_cla32_pg_logic21_and0[0], h_s_cla32_or47[0], h_s_cla32_or48);
  pg_logic pg_logic_h_s_cla32_pg_logic22_out(a[22], b[22], h_s_cla32_pg_logic22_or0, h_s_cla32_pg_logic22_and0, h_s_cla32_pg_logic22_xor0);
  xor_gate xor_gate_h_s_cla32_xor22(h_s_cla32_pg_logic22_xor0[0], h_s_cla32_or48[0], h_s_cla32_xor22);
  and_gate and_gate_h_s_cla32_and96(h_s_cla32_or45[0], h_s_cla32_pg_logic21_or0[0], h_s_cla32_and96);
  and_gate and_gate_h_s_cla32_and97(h_s_cla32_pg_logic22_or0[0], h_s_cla32_pg_logic20_or0[0], h_s_cla32_and97);
  and_gate and_gate_h_s_cla32_and98(h_s_cla32_and96[0], h_s_cla32_and97[0], h_s_cla32_and98);
  and_gate and_gate_h_s_cla32_and99(h_s_cla32_pg_logic20_and0[0], h_s_cla32_pg_logic22_or0[0], h_s_cla32_and99);
  and_gate and_gate_h_s_cla32_and100(h_s_cla32_and99[0], h_s_cla32_pg_logic21_or0[0], h_s_cla32_and100);
  and_gate and_gate_h_s_cla32_and101(h_s_cla32_pg_logic21_and0[0], h_s_cla32_pg_logic22_or0[0], h_s_cla32_and101);
  or_gate or_gate_h_s_cla32_or49(h_s_cla32_and98[0], h_s_cla32_and100[0], h_s_cla32_or49);
  or_gate or_gate_h_s_cla32_or50(h_s_cla32_or49[0], h_s_cla32_and101[0], h_s_cla32_or50);
  or_gate or_gate_h_s_cla32_or51(h_s_cla32_pg_logic22_and0[0], h_s_cla32_or50[0], h_s_cla32_or51);
  pg_logic pg_logic_h_s_cla32_pg_logic23_out(a[23], b[23], h_s_cla32_pg_logic23_or0, h_s_cla32_pg_logic23_and0, h_s_cla32_pg_logic23_xor0);
  xor_gate xor_gate_h_s_cla32_xor23(h_s_cla32_pg_logic23_xor0[0], h_s_cla32_or51[0], h_s_cla32_xor23);
  and_gate and_gate_h_s_cla32_and102(h_s_cla32_or45[0], h_s_cla32_pg_logic22_or0[0], h_s_cla32_and102);
  and_gate and_gate_h_s_cla32_and103(h_s_cla32_pg_logic23_or0[0], h_s_cla32_pg_logic21_or0[0], h_s_cla32_and103);
  and_gate and_gate_h_s_cla32_and104(h_s_cla32_and102[0], h_s_cla32_and103[0], h_s_cla32_and104);
  and_gate and_gate_h_s_cla32_and105(h_s_cla32_and104[0], h_s_cla32_pg_logic20_or0[0], h_s_cla32_and105);
  and_gate and_gate_h_s_cla32_and106(h_s_cla32_pg_logic20_and0[0], h_s_cla32_pg_logic22_or0[0], h_s_cla32_and106);
  and_gate and_gate_h_s_cla32_and107(h_s_cla32_pg_logic23_or0[0], h_s_cla32_pg_logic21_or0[0], h_s_cla32_and107);
  and_gate and_gate_h_s_cla32_and108(h_s_cla32_and106[0], h_s_cla32_and107[0], h_s_cla32_and108);
  and_gate and_gate_h_s_cla32_and109(h_s_cla32_pg_logic21_and0[0], h_s_cla32_pg_logic23_or0[0], h_s_cla32_and109);
  and_gate and_gate_h_s_cla32_and110(h_s_cla32_and109[0], h_s_cla32_pg_logic22_or0[0], h_s_cla32_and110);
  and_gate and_gate_h_s_cla32_and111(h_s_cla32_pg_logic22_and0[0], h_s_cla32_pg_logic23_or0[0], h_s_cla32_and111);
  or_gate or_gate_h_s_cla32_or52(h_s_cla32_and105[0], h_s_cla32_and110[0], h_s_cla32_or52);
  or_gate or_gate_h_s_cla32_or53(h_s_cla32_and108[0], h_s_cla32_and111[0], h_s_cla32_or53);
  or_gate or_gate_h_s_cla32_or54(h_s_cla32_or52[0], h_s_cla32_or53[0], h_s_cla32_or54);
  or_gate or_gate_h_s_cla32_or55(h_s_cla32_pg_logic23_and0[0], h_s_cla32_or54[0], h_s_cla32_or55);
  pg_logic pg_logic_h_s_cla32_pg_logic24_out(a[24], b[24], h_s_cla32_pg_logic24_or0, h_s_cla32_pg_logic24_and0, h_s_cla32_pg_logic24_xor0);
  xor_gate xor_gate_h_s_cla32_xor24(h_s_cla32_pg_logic24_xor0[0], h_s_cla32_or55[0], h_s_cla32_xor24);
  and_gate and_gate_h_s_cla32_and112(h_s_cla32_or55[0], h_s_cla32_pg_logic24_or0[0], h_s_cla32_and112);
  or_gate or_gate_h_s_cla32_or56(h_s_cla32_pg_logic24_and0[0], h_s_cla32_and112[0], h_s_cla32_or56);
  pg_logic pg_logic_h_s_cla32_pg_logic25_out(a[25], b[25], h_s_cla32_pg_logic25_or0, h_s_cla32_pg_logic25_and0, h_s_cla32_pg_logic25_xor0);
  xor_gate xor_gate_h_s_cla32_xor25(h_s_cla32_pg_logic25_xor0[0], h_s_cla32_or56[0], h_s_cla32_xor25);
  and_gate and_gate_h_s_cla32_and113(h_s_cla32_or55[0], h_s_cla32_pg_logic25_or0[0], h_s_cla32_and113);
  and_gate and_gate_h_s_cla32_and114(h_s_cla32_and113[0], h_s_cla32_pg_logic24_or0[0], h_s_cla32_and114);
  and_gate and_gate_h_s_cla32_and115(h_s_cla32_pg_logic24_and0[0], h_s_cla32_pg_logic25_or0[0], h_s_cla32_and115);
  or_gate or_gate_h_s_cla32_or57(h_s_cla32_and114[0], h_s_cla32_and115[0], h_s_cla32_or57);
  or_gate or_gate_h_s_cla32_or58(h_s_cla32_pg_logic25_and0[0], h_s_cla32_or57[0], h_s_cla32_or58);
  pg_logic pg_logic_h_s_cla32_pg_logic26_out(a[26], b[26], h_s_cla32_pg_logic26_or0, h_s_cla32_pg_logic26_and0, h_s_cla32_pg_logic26_xor0);
  xor_gate xor_gate_h_s_cla32_xor26(h_s_cla32_pg_logic26_xor0[0], h_s_cla32_or58[0], h_s_cla32_xor26);
  and_gate and_gate_h_s_cla32_and116(h_s_cla32_or55[0], h_s_cla32_pg_logic25_or0[0], h_s_cla32_and116);
  and_gate and_gate_h_s_cla32_and117(h_s_cla32_pg_logic26_or0[0], h_s_cla32_pg_logic24_or0[0], h_s_cla32_and117);
  and_gate and_gate_h_s_cla32_and118(h_s_cla32_and116[0], h_s_cla32_and117[0], h_s_cla32_and118);
  and_gate and_gate_h_s_cla32_and119(h_s_cla32_pg_logic24_and0[0], h_s_cla32_pg_logic26_or0[0], h_s_cla32_and119);
  and_gate and_gate_h_s_cla32_and120(h_s_cla32_and119[0], h_s_cla32_pg_logic25_or0[0], h_s_cla32_and120);
  and_gate and_gate_h_s_cla32_and121(h_s_cla32_pg_logic25_and0[0], h_s_cla32_pg_logic26_or0[0], h_s_cla32_and121);
  or_gate or_gate_h_s_cla32_or59(h_s_cla32_and118[0], h_s_cla32_and120[0], h_s_cla32_or59);
  or_gate or_gate_h_s_cla32_or60(h_s_cla32_or59[0], h_s_cla32_and121[0], h_s_cla32_or60);
  or_gate or_gate_h_s_cla32_or61(h_s_cla32_pg_logic26_and0[0], h_s_cla32_or60[0], h_s_cla32_or61);
  pg_logic pg_logic_h_s_cla32_pg_logic27_out(a[27], b[27], h_s_cla32_pg_logic27_or0, h_s_cla32_pg_logic27_and0, h_s_cla32_pg_logic27_xor0);
  xor_gate xor_gate_h_s_cla32_xor27(h_s_cla32_pg_logic27_xor0[0], h_s_cla32_or61[0], h_s_cla32_xor27);
  and_gate and_gate_h_s_cla32_and122(h_s_cla32_or55[0], h_s_cla32_pg_logic26_or0[0], h_s_cla32_and122);
  and_gate and_gate_h_s_cla32_and123(h_s_cla32_pg_logic27_or0[0], h_s_cla32_pg_logic25_or0[0], h_s_cla32_and123);
  and_gate and_gate_h_s_cla32_and124(h_s_cla32_and122[0], h_s_cla32_and123[0], h_s_cla32_and124);
  and_gate and_gate_h_s_cla32_and125(h_s_cla32_and124[0], h_s_cla32_pg_logic24_or0[0], h_s_cla32_and125);
  and_gate and_gate_h_s_cla32_and126(h_s_cla32_pg_logic24_and0[0], h_s_cla32_pg_logic26_or0[0], h_s_cla32_and126);
  and_gate and_gate_h_s_cla32_and127(h_s_cla32_pg_logic27_or0[0], h_s_cla32_pg_logic25_or0[0], h_s_cla32_and127);
  and_gate and_gate_h_s_cla32_and128(h_s_cla32_and126[0], h_s_cla32_and127[0], h_s_cla32_and128);
  and_gate and_gate_h_s_cla32_and129(h_s_cla32_pg_logic25_and0[0], h_s_cla32_pg_logic27_or0[0], h_s_cla32_and129);
  and_gate and_gate_h_s_cla32_and130(h_s_cla32_and129[0], h_s_cla32_pg_logic26_or0[0], h_s_cla32_and130);
  and_gate and_gate_h_s_cla32_and131(h_s_cla32_pg_logic26_and0[0], h_s_cla32_pg_logic27_or0[0], h_s_cla32_and131);
  or_gate or_gate_h_s_cla32_or62(h_s_cla32_and125[0], h_s_cla32_and130[0], h_s_cla32_or62);
  or_gate or_gate_h_s_cla32_or63(h_s_cla32_and128[0], h_s_cla32_and131[0], h_s_cla32_or63);
  or_gate or_gate_h_s_cla32_or64(h_s_cla32_or62[0], h_s_cla32_or63[0], h_s_cla32_or64);
  or_gate or_gate_h_s_cla32_or65(h_s_cla32_pg_logic27_and0[0], h_s_cla32_or64[0], h_s_cla32_or65);
  pg_logic pg_logic_h_s_cla32_pg_logic28_out(a[28], b[28], h_s_cla32_pg_logic28_or0, h_s_cla32_pg_logic28_and0, h_s_cla32_pg_logic28_xor0);
  xor_gate xor_gate_h_s_cla32_xor28(h_s_cla32_pg_logic28_xor0[0], h_s_cla32_or65[0], h_s_cla32_xor28);
  and_gate and_gate_h_s_cla32_and132(h_s_cla32_or65[0], h_s_cla32_pg_logic28_or0[0], h_s_cla32_and132);
  or_gate or_gate_h_s_cla32_or66(h_s_cla32_pg_logic28_and0[0], h_s_cla32_and132[0], h_s_cla32_or66);
  pg_logic pg_logic_h_s_cla32_pg_logic29_out(a[29], b[29], h_s_cla32_pg_logic29_or0, h_s_cla32_pg_logic29_and0, h_s_cla32_pg_logic29_xor0);
  xor_gate xor_gate_h_s_cla32_xor29(h_s_cla32_pg_logic29_xor0[0], h_s_cla32_or66[0], h_s_cla32_xor29);
  and_gate and_gate_h_s_cla32_and133(h_s_cla32_or65[0], h_s_cla32_pg_logic29_or0[0], h_s_cla32_and133);
  and_gate and_gate_h_s_cla32_and134(h_s_cla32_and133[0], h_s_cla32_pg_logic28_or0[0], h_s_cla32_and134);
  and_gate and_gate_h_s_cla32_and135(h_s_cla32_pg_logic28_and0[0], h_s_cla32_pg_logic29_or0[0], h_s_cla32_and135);
  or_gate or_gate_h_s_cla32_or67(h_s_cla32_and134[0], h_s_cla32_and135[0], h_s_cla32_or67);
  or_gate or_gate_h_s_cla32_or68(h_s_cla32_pg_logic29_and0[0], h_s_cla32_or67[0], h_s_cla32_or68);
  pg_logic pg_logic_h_s_cla32_pg_logic30_out(a[30], b[30], h_s_cla32_pg_logic30_or0, h_s_cla32_pg_logic30_and0, h_s_cla32_pg_logic30_xor0);
  xor_gate xor_gate_h_s_cla32_xor30(h_s_cla32_pg_logic30_xor0[0], h_s_cla32_or68[0], h_s_cla32_xor30);
  and_gate and_gate_h_s_cla32_and136(h_s_cla32_or65[0], h_s_cla32_pg_logic29_or0[0], h_s_cla32_and136);
  and_gate and_gate_h_s_cla32_and137(h_s_cla32_pg_logic30_or0[0], h_s_cla32_pg_logic28_or0[0], h_s_cla32_and137);
  and_gate and_gate_h_s_cla32_and138(h_s_cla32_and136[0], h_s_cla32_and137[0], h_s_cla32_and138);
  and_gate and_gate_h_s_cla32_and139(h_s_cla32_pg_logic28_and0[0], h_s_cla32_pg_logic30_or0[0], h_s_cla32_and139);
  and_gate and_gate_h_s_cla32_and140(h_s_cla32_and139[0], h_s_cla32_pg_logic29_or0[0], h_s_cla32_and140);
  and_gate and_gate_h_s_cla32_and141(h_s_cla32_pg_logic29_and0[0], h_s_cla32_pg_logic30_or0[0], h_s_cla32_and141);
  or_gate or_gate_h_s_cla32_or69(h_s_cla32_and138[0], h_s_cla32_and140[0], h_s_cla32_or69);
  or_gate or_gate_h_s_cla32_or70(h_s_cla32_or69[0], h_s_cla32_and141[0], h_s_cla32_or70);
  or_gate or_gate_h_s_cla32_or71(h_s_cla32_pg_logic30_and0[0], h_s_cla32_or70[0], h_s_cla32_or71);
  pg_logic pg_logic_h_s_cla32_pg_logic31_out(a[31], b[31], h_s_cla32_pg_logic31_or0, h_s_cla32_pg_logic31_and0, h_s_cla32_pg_logic31_xor0);
  xor_gate xor_gate_h_s_cla32_xor31(h_s_cla32_pg_logic31_xor0[0], h_s_cla32_or71[0], h_s_cla32_xor31);
  and_gate and_gate_h_s_cla32_and142(h_s_cla32_or65[0], h_s_cla32_pg_logic30_or0[0], h_s_cla32_and142);
  and_gate and_gate_h_s_cla32_and143(h_s_cla32_pg_logic31_or0[0], h_s_cla32_pg_logic29_or0[0], h_s_cla32_and143);
  and_gate and_gate_h_s_cla32_and144(h_s_cla32_and142[0], h_s_cla32_and143[0], h_s_cla32_and144);
  and_gate and_gate_h_s_cla32_and145(h_s_cla32_and144[0], h_s_cla32_pg_logic28_or0[0], h_s_cla32_and145);
  and_gate and_gate_h_s_cla32_and146(h_s_cla32_pg_logic28_and0[0], h_s_cla32_pg_logic30_or0[0], h_s_cla32_and146);
  and_gate and_gate_h_s_cla32_and147(h_s_cla32_pg_logic31_or0[0], h_s_cla32_pg_logic29_or0[0], h_s_cla32_and147);
  and_gate and_gate_h_s_cla32_and148(h_s_cla32_and146[0], h_s_cla32_and147[0], h_s_cla32_and148);
  and_gate and_gate_h_s_cla32_and149(h_s_cla32_pg_logic29_and0[0], h_s_cla32_pg_logic31_or0[0], h_s_cla32_and149);
  and_gate and_gate_h_s_cla32_and150(h_s_cla32_and149[0], h_s_cla32_pg_logic30_or0[0], h_s_cla32_and150);
  and_gate and_gate_h_s_cla32_and151(h_s_cla32_pg_logic30_and0[0], h_s_cla32_pg_logic31_or0[0], h_s_cla32_and151);
  or_gate or_gate_h_s_cla32_or72(h_s_cla32_and145[0], h_s_cla32_and150[0], h_s_cla32_or72);
  or_gate or_gate_h_s_cla32_or73(h_s_cla32_and148[0], h_s_cla32_and151[0], h_s_cla32_or73);
  or_gate or_gate_h_s_cla32_or74(h_s_cla32_or72[0], h_s_cla32_or73[0], h_s_cla32_or74);
  or_gate or_gate_h_s_cla32_or75(h_s_cla32_pg_logic31_and0[0], h_s_cla32_or74[0], h_s_cla32_or75);
  xor_gate xor_gate_h_s_cla32_xor32(a[31], b[31], h_s_cla32_xor32);
  xor_gate xor_gate_h_s_cla32_xor33(h_s_cla32_xor32[0], h_s_cla32_or75[0], h_s_cla32_xor33);

  assign h_s_cla32_out[0] = h_s_cla32_pg_logic0_xor0[0];
  assign h_s_cla32_out[1] = h_s_cla32_xor1[0];
  assign h_s_cla32_out[2] = h_s_cla32_xor2[0];
  assign h_s_cla32_out[3] = h_s_cla32_xor3[0];
  assign h_s_cla32_out[4] = h_s_cla32_xor4[0];
  assign h_s_cla32_out[5] = h_s_cla32_xor5[0];
  assign h_s_cla32_out[6] = h_s_cla32_xor6[0];
  assign h_s_cla32_out[7] = h_s_cla32_xor7[0];
  assign h_s_cla32_out[8] = h_s_cla32_xor8[0];
  assign h_s_cla32_out[9] = h_s_cla32_xor9[0];
  assign h_s_cla32_out[10] = h_s_cla32_xor10[0];
  assign h_s_cla32_out[11] = h_s_cla32_xor11[0];
  assign h_s_cla32_out[12] = h_s_cla32_xor12[0];
  assign h_s_cla32_out[13] = h_s_cla32_xor13[0];
  assign h_s_cla32_out[14] = h_s_cla32_xor14[0];
  assign h_s_cla32_out[15] = h_s_cla32_xor15[0];
  assign h_s_cla32_out[16] = h_s_cla32_xor16[0];
  assign h_s_cla32_out[17] = h_s_cla32_xor17[0];
  assign h_s_cla32_out[18] = h_s_cla32_xor18[0];
  assign h_s_cla32_out[19] = h_s_cla32_xor19[0];
  assign h_s_cla32_out[20] = h_s_cla32_xor20[0];
  assign h_s_cla32_out[21] = h_s_cla32_xor21[0];
  assign h_s_cla32_out[22] = h_s_cla32_xor22[0];
  assign h_s_cla32_out[23] = h_s_cla32_xor23[0];
  assign h_s_cla32_out[24] = h_s_cla32_xor24[0];
  assign h_s_cla32_out[25] = h_s_cla32_xor25[0];
  assign h_s_cla32_out[26] = h_s_cla32_xor26[0];
  assign h_s_cla32_out[27] = h_s_cla32_xor27[0];
  assign h_s_cla32_out[28] = h_s_cla32_xor28[0];
  assign h_s_cla32_out[29] = h_s_cla32_xor29[0];
  assign h_s_cla32_out[30] = h_s_cla32_xor30[0];
  assign h_s_cla32_out[31] = h_s_cla32_xor31[0];
  assign h_s_cla32_out[32] = h_s_cla32_xor33[0];
endmodule