module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module mux2to1(input [0:0] d0, input [0:0] d1, input [0:0] sel, output [0:0] mux2to1_xor0);
  wire [0:0] mux2to1_and0;
  wire [0:0] mux2to1_not0;
  wire [0:0] mux2to1_and1;
  and_gate and_gate_mux2to1_and0(.a(d1[0]), .b(sel[0]), .out(mux2to1_and0));
  not_gate not_gate_mux2to1_not0(.a(sel[0]), .out(mux2to1_not0));
  and_gate and_gate_mux2to1_and1(.a(d0[0]), .b(mux2to1_not0[0]), .out(mux2to1_and1));
  xor_gate xor_gate_mux2to1_xor0(.a(mux2to1_and0[0]), .b(mux2to1_and1[0]), .out(mux2to1_xor0));
endmodule

module u_cska32(input [31:0] a, input [31:0] b, output [32:0] u_cska32_out);
  wire [0:0] u_cska32_xor0;
  wire [0:0] u_cska32_ha0_xor0;
  wire [0:0] u_cska32_ha0_and0;
  wire [0:0] u_cska32_xor1;
  wire [0:0] u_cska32_fa0_xor1;
  wire [0:0] u_cska32_fa0_or0;
  wire [0:0] u_cska32_xor2;
  wire [0:0] u_cska32_fa1_xor1;
  wire [0:0] u_cska32_fa1_or0;
  wire [0:0] u_cska32_xor3;
  wire [0:0] u_cska32_fa2_xor1;
  wire [0:0] u_cska32_fa2_or0;
  wire [0:0] u_cska32_and_propagate00;
  wire [0:0] u_cska32_and_propagate01;
  wire [0:0] u_cska32_and_propagate02;
  wire [0:0] u_cska32_mux2to10_and1;
  wire [0:0] u_cska32_xor4;
  wire [0:0] u_cska32_fa3_xor1;
  wire [0:0] u_cska32_fa3_or0;
  wire [0:0] u_cska32_xor5;
  wire [0:0] u_cska32_fa4_xor1;
  wire [0:0] u_cska32_fa4_or0;
  wire [0:0] u_cska32_xor6;
  wire [0:0] u_cska32_fa5_xor1;
  wire [0:0] u_cska32_fa5_or0;
  wire [0:0] u_cska32_xor7;
  wire [0:0] u_cska32_fa6_xor1;
  wire [0:0] u_cska32_fa6_or0;
  wire [0:0] u_cska32_and_propagate13;
  wire [0:0] u_cska32_and_propagate14;
  wire [0:0] u_cska32_and_propagate15;
  wire [0:0] u_cska32_mux2to11_xor0;
  wire [0:0] u_cska32_xor8;
  wire [0:0] u_cska32_fa7_xor1;
  wire [0:0] u_cska32_fa7_or0;
  wire [0:0] u_cska32_xor9;
  wire [0:0] u_cska32_fa8_xor1;
  wire [0:0] u_cska32_fa8_or0;
  wire [0:0] u_cska32_xor10;
  wire [0:0] u_cska32_fa9_xor1;
  wire [0:0] u_cska32_fa9_or0;
  wire [0:0] u_cska32_xor11;
  wire [0:0] u_cska32_fa10_xor1;
  wire [0:0] u_cska32_fa10_or0;
  wire [0:0] u_cska32_and_propagate26;
  wire [0:0] u_cska32_and_propagate27;
  wire [0:0] u_cska32_and_propagate28;
  wire [0:0] u_cska32_mux2to12_xor0;
  wire [0:0] u_cska32_xor12;
  wire [0:0] u_cska32_fa11_xor1;
  wire [0:0] u_cska32_fa11_or0;
  wire [0:0] u_cska32_xor13;
  wire [0:0] u_cska32_fa12_xor1;
  wire [0:0] u_cska32_fa12_or0;
  wire [0:0] u_cska32_xor14;
  wire [0:0] u_cska32_fa13_xor1;
  wire [0:0] u_cska32_fa13_or0;
  wire [0:0] u_cska32_xor15;
  wire [0:0] u_cska32_fa14_xor1;
  wire [0:0] u_cska32_fa14_or0;
  wire [0:0] u_cska32_and_propagate39;
  wire [0:0] u_cska32_and_propagate310;
  wire [0:0] u_cska32_and_propagate311;
  wire [0:0] u_cska32_mux2to13_xor0;
  wire [0:0] u_cska32_xor16;
  wire [0:0] u_cska32_fa15_xor1;
  wire [0:0] u_cska32_fa15_or0;
  wire [0:0] u_cska32_xor17;
  wire [0:0] u_cska32_fa16_xor1;
  wire [0:0] u_cska32_fa16_or0;
  wire [0:0] u_cska32_xor18;
  wire [0:0] u_cska32_fa17_xor1;
  wire [0:0] u_cska32_fa17_or0;
  wire [0:0] u_cska32_xor19;
  wire [0:0] u_cska32_fa18_xor1;
  wire [0:0] u_cska32_fa18_or0;
  wire [0:0] u_cska32_and_propagate412;
  wire [0:0] u_cska32_and_propagate413;
  wire [0:0] u_cska32_and_propagate414;
  wire [0:0] u_cska32_mux2to14_xor0;
  wire [0:0] u_cska32_xor20;
  wire [0:0] u_cska32_fa19_xor1;
  wire [0:0] u_cska32_fa19_or0;
  wire [0:0] u_cska32_xor21;
  wire [0:0] u_cska32_fa20_xor1;
  wire [0:0] u_cska32_fa20_or0;
  wire [0:0] u_cska32_xor22;
  wire [0:0] u_cska32_fa21_xor1;
  wire [0:0] u_cska32_fa21_or0;
  wire [0:0] u_cska32_xor23;
  wire [0:0] u_cska32_fa22_xor1;
  wire [0:0] u_cska32_fa22_or0;
  wire [0:0] u_cska32_and_propagate515;
  wire [0:0] u_cska32_and_propagate516;
  wire [0:0] u_cska32_and_propagate517;
  wire [0:0] u_cska32_mux2to15_xor0;
  wire [0:0] u_cska32_xor24;
  wire [0:0] u_cska32_fa23_xor1;
  wire [0:0] u_cska32_fa23_or0;
  wire [0:0] u_cska32_xor25;
  wire [0:0] u_cska32_fa24_xor1;
  wire [0:0] u_cska32_fa24_or0;
  wire [0:0] u_cska32_xor26;
  wire [0:0] u_cska32_fa25_xor1;
  wire [0:0] u_cska32_fa25_or0;
  wire [0:0] u_cska32_xor27;
  wire [0:0] u_cska32_fa26_xor1;
  wire [0:0] u_cska32_fa26_or0;
  wire [0:0] u_cska32_and_propagate618;
  wire [0:0] u_cska32_and_propagate619;
  wire [0:0] u_cska32_and_propagate620;
  wire [0:0] u_cska32_mux2to16_xor0;
  wire [0:0] u_cska32_xor28;
  wire [0:0] u_cska32_fa27_xor1;
  wire [0:0] u_cska32_fa27_or0;
  wire [0:0] u_cska32_xor29;
  wire [0:0] u_cska32_fa28_xor1;
  wire [0:0] u_cska32_fa28_or0;
  wire [0:0] u_cska32_xor30;
  wire [0:0] u_cska32_fa29_xor1;
  wire [0:0] u_cska32_fa29_or0;
  wire [0:0] u_cska32_xor31;
  wire [0:0] u_cska32_fa30_xor1;
  wire [0:0] u_cska32_fa30_or0;
  wire [0:0] u_cska32_and_propagate721;
  wire [0:0] u_cska32_and_propagate722;
  wire [0:0] u_cska32_and_propagate723;
  wire [0:0] u_cska32_mux2to17_xor0;

  xor_gate xor_gate_u_cska32_xor0(.a(a[0]), .b(b[0]), .out(u_cska32_xor0));
  ha ha_u_cska32_ha0_out(.a(a[0]), .b(b[0]), .ha_xor0(u_cska32_ha0_xor0), .ha_and0(u_cska32_ha0_and0));
  xor_gate xor_gate_u_cska32_xor1(.a(a[1]), .b(b[1]), .out(u_cska32_xor1));
  fa fa_u_cska32_fa0_out(.a(a[1]), .b(b[1]), .cin(u_cska32_ha0_and0[0]), .fa_xor1(u_cska32_fa0_xor1), .fa_or0(u_cska32_fa0_or0));
  xor_gate xor_gate_u_cska32_xor2(.a(a[2]), .b(b[2]), .out(u_cska32_xor2));
  fa fa_u_cska32_fa1_out(.a(a[2]), .b(b[2]), .cin(u_cska32_fa0_or0[0]), .fa_xor1(u_cska32_fa1_xor1), .fa_or0(u_cska32_fa1_or0));
  xor_gate xor_gate_u_cska32_xor3(.a(a[3]), .b(b[3]), .out(u_cska32_xor3));
  fa fa_u_cska32_fa2_out(.a(a[3]), .b(b[3]), .cin(u_cska32_fa1_or0[0]), .fa_xor1(u_cska32_fa2_xor1), .fa_or0(u_cska32_fa2_or0));
  and_gate and_gate_u_cska32_and_propagate00(.a(u_cska32_xor0[0]), .b(u_cska32_xor2[0]), .out(u_cska32_and_propagate00));
  and_gate and_gate_u_cska32_and_propagate01(.a(u_cska32_xor1[0]), .b(u_cska32_xor3[0]), .out(u_cska32_and_propagate01));
  and_gate and_gate_u_cska32_and_propagate02(.a(u_cska32_and_propagate00[0]), .b(u_cska32_and_propagate01[0]), .out(u_cska32_and_propagate02));
  mux2to1 mux2to1_u_cska32_mux2to10_out(.d0(u_cska32_fa2_or0[0]), .d1(1'b0), .sel(u_cska32_and_propagate02[0]), .mux2to1_xor0(u_cska32_mux2to10_and1));
  xor_gate xor_gate_u_cska32_xor4(.a(a[4]), .b(b[4]), .out(u_cska32_xor4));
  fa fa_u_cska32_fa3_out(.a(a[4]), .b(b[4]), .cin(u_cska32_mux2to10_and1[0]), .fa_xor1(u_cska32_fa3_xor1), .fa_or0(u_cska32_fa3_or0));
  xor_gate xor_gate_u_cska32_xor5(.a(a[5]), .b(b[5]), .out(u_cska32_xor5));
  fa fa_u_cska32_fa4_out(.a(a[5]), .b(b[5]), .cin(u_cska32_fa3_or0[0]), .fa_xor1(u_cska32_fa4_xor1), .fa_or0(u_cska32_fa4_or0));
  xor_gate xor_gate_u_cska32_xor6(.a(a[6]), .b(b[6]), .out(u_cska32_xor6));
  fa fa_u_cska32_fa5_out(.a(a[6]), .b(b[6]), .cin(u_cska32_fa4_or0[0]), .fa_xor1(u_cska32_fa5_xor1), .fa_or0(u_cska32_fa5_or0));
  xor_gate xor_gate_u_cska32_xor7(.a(a[7]), .b(b[7]), .out(u_cska32_xor7));
  fa fa_u_cska32_fa6_out(.a(a[7]), .b(b[7]), .cin(u_cska32_fa5_or0[0]), .fa_xor1(u_cska32_fa6_xor1), .fa_or0(u_cska32_fa6_or0));
  and_gate and_gate_u_cska32_and_propagate13(.a(u_cska32_xor4[0]), .b(u_cska32_xor6[0]), .out(u_cska32_and_propagate13));
  and_gate and_gate_u_cska32_and_propagate14(.a(u_cska32_xor5[0]), .b(u_cska32_xor7[0]), .out(u_cska32_and_propagate14));
  and_gate and_gate_u_cska32_and_propagate15(.a(u_cska32_and_propagate13[0]), .b(u_cska32_and_propagate14[0]), .out(u_cska32_and_propagate15));
  mux2to1 mux2to1_u_cska32_mux2to11_out(.d0(u_cska32_fa6_or0[0]), .d1(u_cska32_mux2to10_and1[0]), .sel(u_cska32_and_propagate15[0]), .mux2to1_xor0(u_cska32_mux2to11_xor0));
  xor_gate xor_gate_u_cska32_xor8(.a(a[8]), .b(b[8]), .out(u_cska32_xor8));
  fa fa_u_cska32_fa7_out(.a(a[8]), .b(b[8]), .cin(u_cska32_mux2to11_xor0[0]), .fa_xor1(u_cska32_fa7_xor1), .fa_or0(u_cska32_fa7_or0));
  xor_gate xor_gate_u_cska32_xor9(.a(a[9]), .b(b[9]), .out(u_cska32_xor9));
  fa fa_u_cska32_fa8_out(.a(a[9]), .b(b[9]), .cin(u_cska32_fa7_or0[0]), .fa_xor1(u_cska32_fa8_xor1), .fa_or0(u_cska32_fa8_or0));
  xor_gate xor_gate_u_cska32_xor10(.a(a[10]), .b(b[10]), .out(u_cska32_xor10));
  fa fa_u_cska32_fa9_out(.a(a[10]), .b(b[10]), .cin(u_cska32_fa8_or0[0]), .fa_xor1(u_cska32_fa9_xor1), .fa_or0(u_cska32_fa9_or0));
  xor_gate xor_gate_u_cska32_xor11(.a(a[11]), .b(b[11]), .out(u_cska32_xor11));
  fa fa_u_cska32_fa10_out(.a(a[11]), .b(b[11]), .cin(u_cska32_fa9_or0[0]), .fa_xor1(u_cska32_fa10_xor1), .fa_or0(u_cska32_fa10_or0));
  and_gate and_gate_u_cska32_and_propagate26(.a(u_cska32_xor8[0]), .b(u_cska32_xor10[0]), .out(u_cska32_and_propagate26));
  and_gate and_gate_u_cska32_and_propagate27(.a(u_cska32_xor9[0]), .b(u_cska32_xor11[0]), .out(u_cska32_and_propagate27));
  and_gate and_gate_u_cska32_and_propagate28(.a(u_cska32_and_propagate26[0]), .b(u_cska32_and_propagate27[0]), .out(u_cska32_and_propagate28));
  mux2to1 mux2to1_u_cska32_mux2to12_out(.d0(u_cska32_fa10_or0[0]), .d1(u_cska32_mux2to11_xor0[0]), .sel(u_cska32_and_propagate28[0]), .mux2to1_xor0(u_cska32_mux2to12_xor0));
  xor_gate xor_gate_u_cska32_xor12(.a(a[12]), .b(b[12]), .out(u_cska32_xor12));
  fa fa_u_cska32_fa11_out(.a(a[12]), .b(b[12]), .cin(u_cska32_mux2to12_xor0[0]), .fa_xor1(u_cska32_fa11_xor1), .fa_or0(u_cska32_fa11_or0));
  xor_gate xor_gate_u_cska32_xor13(.a(a[13]), .b(b[13]), .out(u_cska32_xor13));
  fa fa_u_cska32_fa12_out(.a(a[13]), .b(b[13]), .cin(u_cska32_fa11_or0[0]), .fa_xor1(u_cska32_fa12_xor1), .fa_or0(u_cska32_fa12_or0));
  xor_gate xor_gate_u_cska32_xor14(.a(a[14]), .b(b[14]), .out(u_cska32_xor14));
  fa fa_u_cska32_fa13_out(.a(a[14]), .b(b[14]), .cin(u_cska32_fa12_or0[0]), .fa_xor1(u_cska32_fa13_xor1), .fa_or0(u_cska32_fa13_or0));
  xor_gate xor_gate_u_cska32_xor15(.a(a[15]), .b(b[15]), .out(u_cska32_xor15));
  fa fa_u_cska32_fa14_out(.a(a[15]), .b(b[15]), .cin(u_cska32_fa13_or0[0]), .fa_xor1(u_cska32_fa14_xor1), .fa_or0(u_cska32_fa14_or0));
  and_gate and_gate_u_cska32_and_propagate39(.a(u_cska32_xor12[0]), .b(u_cska32_xor14[0]), .out(u_cska32_and_propagate39));
  and_gate and_gate_u_cska32_and_propagate310(.a(u_cska32_xor13[0]), .b(u_cska32_xor15[0]), .out(u_cska32_and_propagate310));
  and_gate and_gate_u_cska32_and_propagate311(.a(u_cska32_and_propagate39[0]), .b(u_cska32_and_propagate310[0]), .out(u_cska32_and_propagate311));
  mux2to1 mux2to1_u_cska32_mux2to13_out(.d0(u_cska32_fa14_or0[0]), .d1(u_cska32_mux2to12_xor0[0]), .sel(u_cska32_and_propagate311[0]), .mux2to1_xor0(u_cska32_mux2to13_xor0));
  xor_gate xor_gate_u_cska32_xor16(.a(a[16]), .b(b[16]), .out(u_cska32_xor16));
  fa fa_u_cska32_fa15_out(.a(a[16]), .b(b[16]), .cin(u_cska32_mux2to13_xor0[0]), .fa_xor1(u_cska32_fa15_xor1), .fa_or0(u_cska32_fa15_or0));
  xor_gate xor_gate_u_cska32_xor17(.a(a[17]), .b(b[17]), .out(u_cska32_xor17));
  fa fa_u_cska32_fa16_out(.a(a[17]), .b(b[17]), .cin(u_cska32_fa15_or0[0]), .fa_xor1(u_cska32_fa16_xor1), .fa_or0(u_cska32_fa16_or0));
  xor_gate xor_gate_u_cska32_xor18(.a(a[18]), .b(b[18]), .out(u_cska32_xor18));
  fa fa_u_cska32_fa17_out(.a(a[18]), .b(b[18]), .cin(u_cska32_fa16_or0[0]), .fa_xor1(u_cska32_fa17_xor1), .fa_or0(u_cska32_fa17_or0));
  xor_gate xor_gate_u_cska32_xor19(.a(a[19]), .b(b[19]), .out(u_cska32_xor19));
  fa fa_u_cska32_fa18_out(.a(a[19]), .b(b[19]), .cin(u_cska32_fa17_or0[0]), .fa_xor1(u_cska32_fa18_xor1), .fa_or0(u_cska32_fa18_or0));
  and_gate and_gate_u_cska32_and_propagate412(.a(u_cska32_xor16[0]), .b(u_cska32_xor18[0]), .out(u_cska32_and_propagate412));
  and_gate and_gate_u_cska32_and_propagate413(.a(u_cska32_xor17[0]), .b(u_cska32_xor19[0]), .out(u_cska32_and_propagate413));
  and_gate and_gate_u_cska32_and_propagate414(.a(u_cska32_and_propagate412[0]), .b(u_cska32_and_propagate413[0]), .out(u_cska32_and_propagate414));
  mux2to1 mux2to1_u_cska32_mux2to14_out(.d0(u_cska32_fa18_or0[0]), .d1(u_cska32_mux2to13_xor0[0]), .sel(u_cska32_and_propagate414[0]), .mux2to1_xor0(u_cska32_mux2to14_xor0));
  xor_gate xor_gate_u_cska32_xor20(.a(a[20]), .b(b[20]), .out(u_cska32_xor20));
  fa fa_u_cska32_fa19_out(.a(a[20]), .b(b[20]), .cin(u_cska32_mux2to14_xor0[0]), .fa_xor1(u_cska32_fa19_xor1), .fa_or0(u_cska32_fa19_or0));
  xor_gate xor_gate_u_cska32_xor21(.a(a[21]), .b(b[21]), .out(u_cska32_xor21));
  fa fa_u_cska32_fa20_out(.a(a[21]), .b(b[21]), .cin(u_cska32_fa19_or0[0]), .fa_xor1(u_cska32_fa20_xor1), .fa_or0(u_cska32_fa20_or0));
  xor_gate xor_gate_u_cska32_xor22(.a(a[22]), .b(b[22]), .out(u_cska32_xor22));
  fa fa_u_cska32_fa21_out(.a(a[22]), .b(b[22]), .cin(u_cska32_fa20_or0[0]), .fa_xor1(u_cska32_fa21_xor1), .fa_or0(u_cska32_fa21_or0));
  xor_gate xor_gate_u_cska32_xor23(.a(a[23]), .b(b[23]), .out(u_cska32_xor23));
  fa fa_u_cska32_fa22_out(.a(a[23]), .b(b[23]), .cin(u_cska32_fa21_or0[0]), .fa_xor1(u_cska32_fa22_xor1), .fa_or0(u_cska32_fa22_or0));
  and_gate and_gate_u_cska32_and_propagate515(.a(u_cska32_xor20[0]), .b(u_cska32_xor22[0]), .out(u_cska32_and_propagate515));
  and_gate and_gate_u_cska32_and_propagate516(.a(u_cska32_xor21[0]), .b(u_cska32_xor23[0]), .out(u_cska32_and_propagate516));
  and_gate and_gate_u_cska32_and_propagate517(.a(u_cska32_and_propagate515[0]), .b(u_cska32_and_propagate516[0]), .out(u_cska32_and_propagate517));
  mux2to1 mux2to1_u_cska32_mux2to15_out(.d0(u_cska32_fa22_or0[0]), .d1(u_cska32_mux2to14_xor0[0]), .sel(u_cska32_and_propagate517[0]), .mux2to1_xor0(u_cska32_mux2to15_xor0));
  xor_gate xor_gate_u_cska32_xor24(.a(a[24]), .b(b[24]), .out(u_cska32_xor24));
  fa fa_u_cska32_fa23_out(.a(a[24]), .b(b[24]), .cin(u_cska32_mux2to15_xor0[0]), .fa_xor1(u_cska32_fa23_xor1), .fa_or0(u_cska32_fa23_or0));
  xor_gate xor_gate_u_cska32_xor25(.a(a[25]), .b(b[25]), .out(u_cska32_xor25));
  fa fa_u_cska32_fa24_out(.a(a[25]), .b(b[25]), .cin(u_cska32_fa23_or0[0]), .fa_xor1(u_cska32_fa24_xor1), .fa_or0(u_cska32_fa24_or0));
  xor_gate xor_gate_u_cska32_xor26(.a(a[26]), .b(b[26]), .out(u_cska32_xor26));
  fa fa_u_cska32_fa25_out(.a(a[26]), .b(b[26]), .cin(u_cska32_fa24_or0[0]), .fa_xor1(u_cska32_fa25_xor1), .fa_or0(u_cska32_fa25_or0));
  xor_gate xor_gate_u_cska32_xor27(.a(a[27]), .b(b[27]), .out(u_cska32_xor27));
  fa fa_u_cska32_fa26_out(.a(a[27]), .b(b[27]), .cin(u_cska32_fa25_or0[0]), .fa_xor1(u_cska32_fa26_xor1), .fa_or0(u_cska32_fa26_or0));
  and_gate and_gate_u_cska32_and_propagate618(.a(u_cska32_xor24[0]), .b(u_cska32_xor26[0]), .out(u_cska32_and_propagate618));
  and_gate and_gate_u_cska32_and_propagate619(.a(u_cska32_xor25[0]), .b(u_cska32_xor27[0]), .out(u_cska32_and_propagate619));
  and_gate and_gate_u_cska32_and_propagate620(.a(u_cska32_and_propagate618[0]), .b(u_cska32_and_propagate619[0]), .out(u_cska32_and_propagate620));
  mux2to1 mux2to1_u_cska32_mux2to16_out(.d0(u_cska32_fa26_or0[0]), .d1(u_cska32_mux2to15_xor0[0]), .sel(u_cska32_and_propagate620[0]), .mux2to1_xor0(u_cska32_mux2to16_xor0));
  xor_gate xor_gate_u_cska32_xor28(.a(a[28]), .b(b[28]), .out(u_cska32_xor28));
  fa fa_u_cska32_fa27_out(.a(a[28]), .b(b[28]), .cin(u_cska32_mux2to16_xor0[0]), .fa_xor1(u_cska32_fa27_xor1), .fa_or0(u_cska32_fa27_or0));
  xor_gate xor_gate_u_cska32_xor29(.a(a[29]), .b(b[29]), .out(u_cska32_xor29));
  fa fa_u_cska32_fa28_out(.a(a[29]), .b(b[29]), .cin(u_cska32_fa27_or0[0]), .fa_xor1(u_cska32_fa28_xor1), .fa_or0(u_cska32_fa28_or0));
  xor_gate xor_gate_u_cska32_xor30(.a(a[30]), .b(b[30]), .out(u_cska32_xor30));
  fa fa_u_cska32_fa29_out(.a(a[30]), .b(b[30]), .cin(u_cska32_fa28_or0[0]), .fa_xor1(u_cska32_fa29_xor1), .fa_or0(u_cska32_fa29_or0));
  xor_gate xor_gate_u_cska32_xor31(.a(a[31]), .b(b[31]), .out(u_cska32_xor31));
  fa fa_u_cska32_fa30_out(.a(a[31]), .b(b[31]), .cin(u_cska32_fa29_or0[0]), .fa_xor1(u_cska32_fa30_xor1), .fa_or0(u_cska32_fa30_or0));
  and_gate and_gate_u_cska32_and_propagate721(.a(u_cska32_xor28[0]), .b(u_cska32_xor30[0]), .out(u_cska32_and_propagate721));
  and_gate and_gate_u_cska32_and_propagate722(.a(u_cska32_xor29[0]), .b(u_cska32_xor31[0]), .out(u_cska32_and_propagate722));
  and_gate and_gate_u_cska32_and_propagate723(.a(u_cska32_and_propagate721[0]), .b(u_cska32_and_propagate722[0]), .out(u_cska32_and_propagate723));
  mux2to1 mux2to1_u_cska32_mux2to17_out(.d0(u_cska32_fa30_or0[0]), .d1(u_cska32_mux2to16_xor0[0]), .sel(u_cska32_and_propagate723[0]), .mux2to1_xor0(u_cska32_mux2to17_xor0));

  assign u_cska32_out[0] = u_cska32_ha0_xor0[0];
  assign u_cska32_out[1] = u_cska32_fa0_xor1[0];
  assign u_cska32_out[2] = u_cska32_fa1_xor1[0];
  assign u_cska32_out[3] = u_cska32_fa2_xor1[0];
  assign u_cska32_out[4] = u_cska32_fa3_xor1[0];
  assign u_cska32_out[5] = u_cska32_fa4_xor1[0];
  assign u_cska32_out[6] = u_cska32_fa5_xor1[0];
  assign u_cska32_out[7] = u_cska32_fa6_xor1[0];
  assign u_cska32_out[8] = u_cska32_fa7_xor1[0];
  assign u_cska32_out[9] = u_cska32_fa8_xor1[0];
  assign u_cska32_out[10] = u_cska32_fa9_xor1[0];
  assign u_cska32_out[11] = u_cska32_fa10_xor1[0];
  assign u_cska32_out[12] = u_cska32_fa11_xor1[0];
  assign u_cska32_out[13] = u_cska32_fa12_xor1[0];
  assign u_cska32_out[14] = u_cska32_fa13_xor1[0];
  assign u_cska32_out[15] = u_cska32_fa14_xor1[0];
  assign u_cska32_out[16] = u_cska32_fa15_xor1[0];
  assign u_cska32_out[17] = u_cska32_fa16_xor1[0];
  assign u_cska32_out[18] = u_cska32_fa17_xor1[0];
  assign u_cska32_out[19] = u_cska32_fa18_xor1[0];
  assign u_cska32_out[20] = u_cska32_fa19_xor1[0];
  assign u_cska32_out[21] = u_cska32_fa20_xor1[0];
  assign u_cska32_out[22] = u_cska32_fa21_xor1[0];
  assign u_cska32_out[23] = u_cska32_fa22_xor1[0];
  assign u_cska32_out[24] = u_cska32_fa23_xor1[0];
  assign u_cska32_out[25] = u_cska32_fa24_xor1[0];
  assign u_cska32_out[26] = u_cska32_fa25_xor1[0];
  assign u_cska32_out[27] = u_cska32_fa26_xor1[0];
  assign u_cska32_out[28] = u_cska32_fa27_xor1[0];
  assign u_cska32_out[29] = u_cska32_fa28_xor1[0];
  assign u_cska32_out[30] = u_cska32_fa29_xor1[0];
  assign u_cska32_out[31] = u_cska32_fa30_xor1[0];
  assign u_cska32_out[32] = u_cska32_mux2to17_xor0[0];
endmodule

module u_csamul_cska32(input [31:0] a, input [31:0] b, output [63:0] u_csamul_cska32_out);
  wire [0:0] u_csamul_cska32_and0_0;
  wire [0:0] u_csamul_cska32_and1_0;
  wire [0:0] u_csamul_cska32_and2_0;
  wire [0:0] u_csamul_cska32_and3_0;
  wire [0:0] u_csamul_cska32_and4_0;
  wire [0:0] u_csamul_cska32_and5_0;
  wire [0:0] u_csamul_cska32_and6_0;
  wire [0:0] u_csamul_cska32_and7_0;
  wire [0:0] u_csamul_cska32_and8_0;
  wire [0:0] u_csamul_cska32_and9_0;
  wire [0:0] u_csamul_cska32_and10_0;
  wire [0:0] u_csamul_cska32_and11_0;
  wire [0:0] u_csamul_cska32_and12_0;
  wire [0:0] u_csamul_cska32_and13_0;
  wire [0:0] u_csamul_cska32_and14_0;
  wire [0:0] u_csamul_cska32_and15_0;
  wire [0:0] u_csamul_cska32_and16_0;
  wire [0:0] u_csamul_cska32_and17_0;
  wire [0:0] u_csamul_cska32_and18_0;
  wire [0:0] u_csamul_cska32_and19_0;
  wire [0:0] u_csamul_cska32_and20_0;
  wire [0:0] u_csamul_cska32_and21_0;
  wire [0:0] u_csamul_cska32_and22_0;
  wire [0:0] u_csamul_cska32_and23_0;
  wire [0:0] u_csamul_cska32_and24_0;
  wire [0:0] u_csamul_cska32_and25_0;
  wire [0:0] u_csamul_cska32_and26_0;
  wire [0:0] u_csamul_cska32_and27_0;
  wire [0:0] u_csamul_cska32_and28_0;
  wire [0:0] u_csamul_cska32_and29_0;
  wire [0:0] u_csamul_cska32_and30_0;
  wire [0:0] u_csamul_cska32_and31_0;
  wire [0:0] u_csamul_cska32_and0_1;
  wire [0:0] u_csamul_cska32_ha0_1_xor0;
  wire [0:0] u_csamul_cska32_ha0_1_and0;
  wire [0:0] u_csamul_cska32_and1_1;
  wire [0:0] u_csamul_cska32_ha1_1_xor0;
  wire [0:0] u_csamul_cska32_ha1_1_and0;
  wire [0:0] u_csamul_cska32_and2_1;
  wire [0:0] u_csamul_cska32_ha2_1_xor0;
  wire [0:0] u_csamul_cska32_ha2_1_and0;
  wire [0:0] u_csamul_cska32_and3_1;
  wire [0:0] u_csamul_cska32_ha3_1_xor0;
  wire [0:0] u_csamul_cska32_ha3_1_and0;
  wire [0:0] u_csamul_cska32_and4_1;
  wire [0:0] u_csamul_cska32_ha4_1_xor0;
  wire [0:0] u_csamul_cska32_ha4_1_and0;
  wire [0:0] u_csamul_cska32_and5_1;
  wire [0:0] u_csamul_cska32_ha5_1_xor0;
  wire [0:0] u_csamul_cska32_ha5_1_and0;
  wire [0:0] u_csamul_cska32_and6_1;
  wire [0:0] u_csamul_cska32_ha6_1_xor0;
  wire [0:0] u_csamul_cska32_ha6_1_and0;
  wire [0:0] u_csamul_cska32_and7_1;
  wire [0:0] u_csamul_cska32_ha7_1_xor0;
  wire [0:0] u_csamul_cska32_ha7_1_and0;
  wire [0:0] u_csamul_cska32_and8_1;
  wire [0:0] u_csamul_cska32_ha8_1_xor0;
  wire [0:0] u_csamul_cska32_ha8_1_and0;
  wire [0:0] u_csamul_cska32_and9_1;
  wire [0:0] u_csamul_cska32_ha9_1_xor0;
  wire [0:0] u_csamul_cska32_ha9_1_and0;
  wire [0:0] u_csamul_cska32_and10_1;
  wire [0:0] u_csamul_cska32_ha10_1_xor0;
  wire [0:0] u_csamul_cska32_ha10_1_and0;
  wire [0:0] u_csamul_cska32_and11_1;
  wire [0:0] u_csamul_cska32_ha11_1_xor0;
  wire [0:0] u_csamul_cska32_ha11_1_and0;
  wire [0:0] u_csamul_cska32_and12_1;
  wire [0:0] u_csamul_cska32_ha12_1_xor0;
  wire [0:0] u_csamul_cska32_ha12_1_and0;
  wire [0:0] u_csamul_cska32_and13_1;
  wire [0:0] u_csamul_cska32_ha13_1_xor0;
  wire [0:0] u_csamul_cska32_ha13_1_and0;
  wire [0:0] u_csamul_cska32_and14_1;
  wire [0:0] u_csamul_cska32_ha14_1_xor0;
  wire [0:0] u_csamul_cska32_ha14_1_and0;
  wire [0:0] u_csamul_cska32_and15_1;
  wire [0:0] u_csamul_cska32_ha15_1_xor0;
  wire [0:0] u_csamul_cska32_ha15_1_and0;
  wire [0:0] u_csamul_cska32_and16_1;
  wire [0:0] u_csamul_cska32_ha16_1_xor0;
  wire [0:0] u_csamul_cska32_ha16_1_and0;
  wire [0:0] u_csamul_cska32_and17_1;
  wire [0:0] u_csamul_cska32_ha17_1_xor0;
  wire [0:0] u_csamul_cska32_ha17_1_and0;
  wire [0:0] u_csamul_cska32_and18_1;
  wire [0:0] u_csamul_cska32_ha18_1_xor0;
  wire [0:0] u_csamul_cska32_ha18_1_and0;
  wire [0:0] u_csamul_cska32_and19_1;
  wire [0:0] u_csamul_cska32_ha19_1_xor0;
  wire [0:0] u_csamul_cska32_ha19_1_and0;
  wire [0:0] u_csamul_cska32_and20_1;
  wire [0:0] u_csamul_cska32_ha20_1_xor0;
  wire [0:0] u_csamul_cska32_ha20_1_and0;
  wire [0:0] u_csamul_cska32_and21_1;
  wire [0:0] u_csamul_cska32_ha21_1_xor0;
  wire [0:0] u_csamul_cska32_ha21_1_and0;
  wire [0:0] u_csamul_cska32_and22_1;
  wire [0:0] u_csamul_cska32_ha22_1_xor0;
  wire [0:0] u_csamul_cska32_ha22_1_and0;
  wire [0:0] u_csamul_cska32_and23_1;
  wire [0:0] u_csamul_cska32_ha23_1_xor0;
  wire [0:0] u_csamul_cska32_ha23_1_and0;
  wire [0:0] u_csamul_cska32_and24_1;
  wire [0:0] u_csamul_cska32_ha24_1_xor0;
  wire [0:0] u_csamul_cska32_ha24_1_and0;
  wire [0:0] u_csamul_cska32_and25_1;
  wire [0:0] u_csamul_cska32_ha25_1_xor0;
  wire [0:0] u_csamul_cska32_ha25_1_and0;
  wire [0:0] u_csamul_cska32_and26_1;
  wire [0:0] u_csamul_cska32_ha26_1_xor0;
  wire [0:0] u_csamul_cska32_ha26_1_and0;
  wire [0:0] u_csamul_cska32_and27_1;
  wire [0:0] u_csamul_cska32_ha27_1_xor0;
  wire [0:0] u_csamul_cska32_ha27_1_and0;
  wire [0:0] u_csamul_cska32_and28_1;
  wire [0:0] u_csamul_cska32_ha28_1_xor0;
  wire [0:0] u_csamul_cska32_ha28_1_and0;
  wire [0:0] u_csamul_cska32_and29_1;
  wire [0:0] u_csamul_cska32_ha29_1_xor0;
  wire [0:0] u_csamul_cska32_ha29_1_and0;
  wire [0:0] u_csamul_cska32_and30_1;
  wire [0:0] u_csamul_cska32_ha30_1_xor0;
  wire [0:0] u_csamul_cska32_ha30_1_and0;
  wire [0:0] u_csamul_cska32_and31_1;
  wire [0:0] u_csamul_cska32_and0_2;
  wire [0:0] u_csamul_cska32_fa0_2_xor1;
  wire [0:0] u_csamul_cska32_fa0_2_or0;
  wire [0:0] u_csamul_cska32_and1_2;
  wire [0:0] u_csamul_cska32_fa1_2_xor1;
  wire [0:0] u_csamul_cska32_fa1_2_or0;
  wire [0:0] u_csamul_cska32_and2_2;
  wire [0:0] u_csamul_cska32_fa2_2_xor1;
  wire [0:0] u_csamul_cska32_fa2_2_or0;
  wire [0:0] u_csamul_cska32_and3_2;
  wire [0:0] u_csamul_cska32_fa3_2_xor1;
  wire [0:0] u_csamul_cska32_fa3_2_or0;
  wire [0:0] u_csamul_cska32_and4_2;
  wire [0:0] u_csamul_cska32_fa4_2_xor1;
  wire [0:0] u_csamul_cska32_fa4_2_or0;
  wire [0:0] u_csamul_cska32_and5_2;
  wire [0:0] u_csamul_cska32_fa5_2_xor1;
  wire [0:0] u_csamul_cska32_fa5_2_or0;
  wire [0:0] u_csamul_cska32_and6_2;
  wire [0:0] u_csamul_cska32_fa6_2_xor1;
  wire [0:0] u_csamul_cska32_fa6_2_or0;
  wire [0:0] u_csamul_cska32_and7_2;
  wire [0:0] u_csamul_cska32_fa7_2_xor1;
  wire [0:0] u_csamul_cska32_fa7_2_or0;
  wire [0:0] u_csamul_cska32_and8_2;
  wire [0:0] u_csamul_cska32_fa8_2_xor1;
  wire [0:0] u_csamul_cska32_fa8_2_or0;
  wire [0:0] u_csamul_cska32_and9_2;
  wire [0:0] u_csamul_cska32_fa9_2_xor1;
  wire [0:0] u_csamul_cska32_fa9_2_or0;
  wire [0:0] u_csamul_cska32_and10_2;
  wire [0:0] u_csamul_cska32_fa10_2_xor1;
  wire [0:0] u_csamul_cska32_fa10_2_or0;
  wire [0:0] u_csamul_cska32_and11_2;
  wire [0:0] u_csamul_cska32_fa11_2_xor1;
  wire [0:0] u_csamul_cska32_fa11_2_or0;
  wire [0:0] u_csamul_cska32_and12_2;
  wire [0:0] u_csamul_cska32_fa12_2_xor1;
  wire [0:0] u_csamul_cska32_fa12_2_or0;
  wire [0:0] u_csamul_cska32_and13_2;
  wire [0:0] u_csamul_cska32_fa13_2_xor1;
  wire [0:0] u_csamul_cska32_fa13_2_or0;
  wire [0:0] u_csamul_cska32_and14_2;
  wire [0:0] u_csamul_cska32_fa14_2_xor1;
  wire [0:0] u_csamul_cska32_fa14_2_or0;
  wire [0:0] u_csamul_cska32_and15_2;
  wire [0:0] u_csamul_cska32_fa15_2_xor1;
  wire [0:0] u_csamul_cska32_fa15_2_or0;
  wire [0:0] u_csamul_cska32_and16_2;
  wire [0:0] u_csamul_cska32_fa16_2_xor1;
  wire [0:0] u_csamul_cska32_fa16_2_or0;
  wire [0:0] u_csamul_cska32_and17_2;
  wire [0:0] u_csamul_cska32_fa17_2_xor1;
  wire [0:0] u_csamul_cska32_fa17_2_or0;
  wire [0:0] u_csamul_cska32_and18_2;
  wire [0:0] u_csamul_cska32_fa18_2_xor1;
  wire [0:0] u_csamul_cska32_fa18_2_or0;
  wire [0:0] u_csamul_cska32_and19_2;
  wire [0:0] u_csamul_cska32_fa19_2_xor1;
  wire [0:0] u_csamul_cska32_fa19_2_or0;
  wire [0:0] u_csamul_cska32_and20_2;
  wire [0:0] u_csamul_cska32_fa20_2_xor1;
  wire [0:0] u_csamul_cska32_fa20_2_or0;
  wire [0:0] u_csamul_cska32_and21_2;
  wire [0:0] u_csamul_cska32_fa21_2_xor1;
  wire [0:0] u_csamul_cska32_fa21_2_or0;
  wire [0:0] u_csamul_cska32_and22_2;
  wire [0:0] u_csamul_cska32_fa22_2_xor1;
  wire [0:0] u_csamul_cska32_fa22_2_or0;
  wire [0:0] u_csamul_cska32_and23_2;
  wire [0:0] u_csamul_cska32_fa23_2_xor1;
  wire [0:0] u_csamul_cska32_fa23_2_or0;
  wire [0:0] u_csamul_cska32_and24_2;
  wire [0:0] u_csamul_cska32_fa24_2_xor1;
  wire [0:0] u_csamul_cska32_fa24_2_or0;
  wire [0:0] u_csamul_cska32_and25_2;
  wire [0:0] u_csamul_cska32_fa25_2_xor1;
  wire [0:0] u_csamul_cska32_fa25_2_or0;
  wire [0:0] u_csamul_cska32_and26_2;
  wire [0:0] u_csamul_cska32_fa26_2_xor1;
  wire [0:0] u_csamul_cska32_fa26_2_or0;
  wire [0:0] u_csamul_cska32_and27_2;
  wire [0:0] u_csamul_cska32_fa27_2_xor1;
  wire [0:0] u_csamul_cska32_fa27_2_or0;
  wire [0:0] u_csamul_cska32_and28_2;
  wire [0:0] u_csamul_cska32_fa28_2_xor1;
  wire [0:0] u_csamul_cska32_fa28_2_or0;
  wire [0:0] u_csamul_cska32_and29_2;
  wire [0:0] u_csamul_cska32_fa29_2_xor1;
  wire [0:0] u_csamul_cska32_fa29_2_or0;
  wire [0:0] u_csamul_cska32_and30_2;
  wire [0:0] u_csamul_cska32_fa30_2_xor1;
  wire [0:0] u_csamul_cska32_fa30_2_or0;
  wire [0:0] u_csamul_cska32_and31_2;
  wire [0:0] u_csamul_cska32_and0_3;
  wire [0:0] u_csamul_cska32_fa0_3_xor1;
  wire [0:0] u_csamul_cska32_fa0_3_or0;
  wire [0:0] u_csamul_cska32_and1_3;
  wire [0:0] u_csamul_cska32_fa1_3_xor1;
  wire [0:0] u_csamul_cska32_fa1_3_or0;
  wire [0:0] u_csamul_cska32_and2_3;
  wire [0:0] u_csamul_cska32_fa2_3_xor1;
  wire [0:0] u_csamul_cska32_fa2_3_or0;
  wire [0:0] u_csamul_cska32_and3_3;
  wire [0:0] u_csamul_cska32_fa3_3_xor1;
  wire [0:0] u_csamul_cska32_fa3_3_or0;
  wire [0:0] u_csamul_cska32_and4_3;
  wire [0:0] u_csamul_cska32_fa4_3_xor1;
  wire [0:0] u_csamul_cska32_fa4_3_or0;
  wire [0:0] u_csamul_cska32_and5_3;
  wire [0:0] u_csamul_cska32_fa5_3_xor1;
  wire [0:0] u_csamul_cska32_fa5_3_or0;
  wire [0:0] u_csamul_cska32_and6_3;
  wire [0:0] u_csamul_cska32_fa6_3_xor1;
  wire [0:0] u_csamul_cska32_fa6_3_or0;
  wire [0:0] u_csamul_cska32_and7_3;
  wire [0:0] u_csamul_cska32_fa7_3_xor1;
  wire [0:0] u_csamul_cska32_fa7_3_or0;
  wire [0:0] u_csamul_cska32_and8_3;
  wire [0:0] u_csamul_cska32_fa8_3_xor1;
  wire [0:0] u_csamul_cska32_fa8_3_or0;
  wire [0:0] u_csamul_cska32_and9_3;
  wire [0:0] u_csamul_cska32_fa9_3_xor1;
  wire [0:0] u_csamul_cska32_fa9_3_or0;
  wire [0:0] u_csamul_cska32_and10_3;
  wire [0:0] u_csamul_cska32_fa10_3_xor1;
  wire [0:0] u_csamul_cska32_fa10_3_or0;
  wire [0:0] u_csamul_cska32_and11_3;
  wire [0:0] u_csamul_cska32_fa11_3_xor1;
  wire [0:0] u_csamul_cska32_fa11_3_or0;
  wire [0:0] u_csamul_cska32_and12_3;
  wire [0:0] u_csamul_cska32_fa12_3_xor1;
  wire [0:0] u_csamul_cska32_fa12_3_or0;
  wire [0:0] u_csamul_cska32_and13_3;
  wire [0:0] u_csamul_cska32_fa13_3_xor1;
  wire [0:0] u_csamul_cska32_fa13_3_or0;
  wire [0:0] u_csamul_cska32_and14_3;
  wire [0:0] u_csamul_cska32_fa14_3_xor1;
  wire [0:0] u_csamul_cska32_fa14_3_or0;
  wire [0:0] u_csamul_cska32_and15_3;
  wire [0:0] u_csamul_cska32_fa15_3_xor1;
  wire [0:0] u_csamul_cska32_fa15_3_or0;
  wire [0:0] u_csamul_cska32_and16_3;
  wire [0:0] u_csamul_cska32_fa16_3_xor1;
  wire [0:0] u_csamul_cska32_fa16_3_or0;
  wire [0:0] u_csamul_cska32_and17_3;
  wire [0:0] u_csamul_cska32_fa17_3_xor1;
  wire [0:0] u_csamul_cska32_fa17_3_or0;
  wire [0:0] u_csamul_cska32_and18_3;
  wire [0:0] u_csamul_cska32_fa18_3_xor1;
  wire [0:0] u_csamul_cska32_fa18_3_or0;
  wire [0:0] u_csamul_cska32_and19_3;
  wire [0:0] u_csamul_cska32_fa19_3_xor1;
  wire [0:0] u_csamul_cska32_fa19_3_or0;
  wire [0:0] u_csamul_cska32_and20_3;
  wire [0:0] u_csamul_cska32_fa20_3_xor1;
  wire [0:0] u_csamul_cska32_fa20_3_or0;
  wire [0:0] u_csamul_cska32_and21_3;
  wire [0:0] u_csamul_cska32_fa21_3_xor1;
  wire [0:0] u_csamul_cska32_fa21_3_or0;
  wire [0:0] u_csamul_cska32_and22_3;
  wire [0:0] u_csamul_cska32_fa22_3_xor1;
  wire [0:0] u_csamul_cska32_fa22_3_or0;
  wire [0:0] u_csamul_cska32_and23_3;
  wire [0:0] u_csamul_cska32_fa23_3_xor1;
  wire [0:0] u_csamul_cska32_fa23_3_or0;
  wire [0:0] u_csamul_cska32_and24_3;
  wire [0:0] u_csamul_cska32_fa24_3_xor1;
  wire [0:0] u_csamul_cska32_fa24_3_or0;
  wire [0:0] u_csamul_cska32_and25_3;
  wire [0:0] u_csamul_cska32_fa25_3_xor1;
  wire [0:0] u_csamul_cska32_fa25_3_or0;
  wire [0:0] u_csamul_cska32_and26_3;
  wire [0:0] u_csamul_cska32_fa26_3_xor1;
  wire [0:0] u_csamul_cska32_fa26_3_or0;
  wire [0:0] u_csamul_cska32_and27_3;
  wire [0:0] u_csamul_cska32_fa27_3_xor1;
  wire [0:0] u_csamul_cska32_fa27_3_or0;
  wire [0:0] u_csamul_cska32_and28_3;
  wire [0:0] u_csamul_cska32_fa28_3_xor1;
  wire [0:0] u_csamul_cska32_fa28_3_or0;
  wire [0:0] u_csamul_cska32_and29_3;
  wire [0:0] u_csamul_cska32_fa29_3_xor1;
  wire [0:0] u_csamul_cska32_fa29_3_or0;
  wire [0:0] u_csamul_cska32_and30_3;
  wire [0:0] u_csamul_cska32_fa30_3_xor1;
  wire [0:0] u_csamul_cska32_fa30_3_or0;
  wire [0:0] u_csamul_cska32_and31_3;
  wire [0:0] u_csamul_cska32_and0_4;
  wire [0:0] u_csamul_cska32_fa0_4_xor1;
  wire [0:0] u_csamul_cska32_fa0_4_or0;
  wire [0:0] u_csamul_cska32_and1_4;
  wire [0:0] u_csamul_cska32_fa1_4_xor1;
  wire [0:0] u_csamul_cska32_fa1_4_or0;
  wire [0:0] u_csamul_cska32_and2_4;
  wire [0:0] u_csamul_cska32_fa2_4_xor1;
  wire [0:0] u_csamul_cska32_fa2_4_or0;
  wire [0:0] u_csamul_cska32_and3_4;
  wire [0:0] u_csamul_cska32_fa3_4_xor1;
  wire [0:0] u_csamul_cska32_fa3_4_or0;
  wire [0:0] u_csamul_cska32_and4_4;
  wire [0:0] u_csamul_cska32_fa4_4_xor1;
  wire [0:0] u_csamul_cska32_fa4_4_or0;
  wire [0:0] u_csamul_cska32_and5_4;
  wire [0:0] u_csamul_cska32_fa5_4_xor1;
  wire [0:0] u_csamul_cska32_fa5_4_or0;
  wire [0:0] u_csamul_cska32_and6_4;
  wire [0:0] u_csamul_cska32_fa6_4_xor1;
  wire [0:0] u_csamul_cska32_fa6_4_or0;
  wire [0:0] u_csamul_cska32_and7_4;
  wire [0:0] u_csamul_cska32_fa7_4_xor1;
  wire [0:0] u_csamul_cska32_fa7_4_or0;
  wire [0:0] u_csamul_cska32_and8_4;
  wire [0:0] u_csamul_cska32_fa8_4_xor1;
  wire [0:0] u_csamul_cska32_fa8_4_or0;
  wire [0:0] u_csamul_cska32_and9_4;
  wire [0:0] u_csamul_cska32_fa9_4_xor1;
  wire [0:0] u_csamul_cska32_fa9_4_or0;
  wire [0:0] u_csamul_cska32_and10_4;
  wire [0:0] u_csamul_cska32_fa10_4_xor1;
  wire [0:0] u_csamul_cska32_fa10_4_or0;
  wire [0:0] u_csamul_cska32_and11_4;
  wire [0:0] u_csamul_cska32_fa11_4_xor1;
  wire [0:0] u_csamul_cska32_fa11_4_or0;
  wire [0:0] u_csamul_cska32_and12_4;
  wire [0:0] u_csamul_cska32_fa12_4_xor1;
  wire [0:0] u_csamul_cska32_fa12_4_or0;
  wire [0:0] u_csamul_cska32_and13_4;
  wire [0:0] u_csamul_cska32_fa13_4_xor1;
  wire [0:0] u_csamul_cska32_fa13_4_or0;
  wire [0:0] u_csamul_cska32_and14_4;
  wire [0:0] u_csamul_cska32_fa14_4_xor1;
  wire [0:0] u_csamul_cska32_fa14_4_or0;
  wire [0:0] u_csamul_cska32_and15_4;
  wire [0:0] u_csamul_cska32_fa15_4_xor1;
  wire [0:0] u_csamul_cska32_fa15_4_or0;
  wire [0:0] u_csamul_cska32_and16_4;
  wire [0:0] u_csamul_cska32_fa16_4_xor1;
  wire [0:0] u_csamul_cska32_fa16_4_or0;
  wire [0:0] u_csamul_cska32_and17_4;
  wire [0:0] u_csamul_cska32_fa17_4_xor1;
  wire [0:0] u_csamul_cska32_fa17_4_or0;
  wire [0:0] u_csamul_cska32_and18_4;
  wire [0:0] u_csamul_cska32_fa18_4_xor1;
  wire [0:0] u_csamul_cska32_fa18_4_or0;
  wire [0:0] u_csamul_cska32_and19_4;
  wire [0:0] u_csamul_cska32_fa19_4_xor1;
  wire [0:0] u_csamul_cska32_fa19_4_or0;
  wire [0:0] u_csamul_cska32_and20_4;
  wire [0:0] u_csamul_cska32_fa20_4_xor1;
  wire [0:0] u_csamul_cska32_fa20_4_or0;
  wire [0:0] u_csamul_cska32_and21_4;
  wire [0:0] u_csamul_cska32_fa21_4_xor1;
  wire [0:0] u_csamul_cska32_fa21_4_or0;
  wire [0:0] u_csamul_cska32_and22_4;
  wire [0:0] u_csamul_cska32_fa22_4_xor1;
  wire [0:0] u_csamul_cska32_fa22_4_or0;
  wire [0:0] u_csamul_cska32_and23_4;
  wire [0:0] u_csamul_cska32_fa23_4_xor1;
  wire [0:0] u_csamul_cska32_fa23_4_or0;
  wire [0:0] u_csamul_cska32_and24_4;
  wire [0:0] u_csamul_cska32_fa24_4_xor1;
  wire [0:0] u_csamul_cska32_fa24_4_or0;
  wire [0:0] u_csamul_cska32_and25_4;
  wire [0:0] u_csamul_cska32_fa25_4_xor1;
  wire [0:0] u_csamul_cska32_fa25_4_or0;
  wire [0:0] u_csamul_cska32_and26_4;
  wire [0:0] u_csamul_cska32_fa26_4_xor1;
  wire [0:0] u_csamul_cska32_fa26_4_or0;
  wire [0:0] u_csamul_cska32_and27_4;
  wire [0:0] u_csamul_cska32_fa27_4_xor1;
  wire [0:0] u_csamul_cska32_fa27_4_or0;
  wire [0:0] u_csamul_cska32_and28_4;
  wire [0:0] u_csamul_cska32_fa28_4_xor1;
  wire [0:0] u_csamul_cska32_fa28_4_or0;
  wire [0:0] u_csamul_cska32_and29_4;
  wire [0:0] u_csamul_cska32_fa29_4_xor1;
  wire [0:0] u_csamul_cska32_fa29_4_or0;
  wire [0:0] u_csamul_cska32_and30_4;
  wire [0:0] u_csamul_cska32_fa30_4_xor1;
  wire [0:0] u_csamul_cska32_fa30_4_or0;
  wire [0:0] u_csamul_cska32_and31_4;
  wire [0:0] u_csamul_cska32_and0_5;
  wire [0:0] u_csamul_cska32_fa0_5_xor1;
  wire [0:0] u_csamul_cska32_fa0_5_or0;
  wire [0:0] u_csamul_cska32_and1_5;
  wire [0:0] u_csamul_cska32_fa1_5_xor1;
  wire [0:0] u_csamul_cska32_fa1_5_or0;
  wire [0:0] u_csamul_cska32_and2_5;
  wire [0:0] u_csamul_cska32_fa2_5_xor1;
  wire [0:0] u_csamul_cska32_fa2_5_or0;
  wire [0:0] u_csamul_cska32_and3_5;
  wire [0:0] u_csamul_cska32_fa3_5_xor1;
  wire [0:0] u_csamul_cska32_fa3_5_or0;
  wire [0:0] u_csamul_cska32_and4_5;
  wire [0:0] u_csamul_cska32_fa4_5_xor1;
  wire [0:0] u_csamul_cska32_fa4_5_or0;
  wire [0:0] u_csamul_cska32_and5_5;
  wire [0:0] u_csamul_cska32_fa5_5_xor1;
  wire [0:0] u_csamul_cska32_fa5_5_or0;
  wire [0:0] u_csamul_cska32_and6_5;
  wire [0:0] u_csamul_cska32_fa6_5_xor1;
  wire [0:0] u_csamul_cska32_fa6_5_or0;
  wire [0:0] u_csamul_cska32_and7_5;
  wire [0:0] u_csamul_cska32_fa7_5_xor1;
  wire [0:0] u_csamul_cska32_fa7_5_or0;
  wire [0:0] u_csamul_cska32_and8_5;
  wire [0:0] u_csamul_cska32_fa8_5_xor1;
  wire [0:0] u_csamul_cska32_fa8_5_or0;
  wire [0:0] u_csamul_cska32_and9_5;
  wire [0:0] u_csamul_cska32_fa9_5_xor1;
  wire [0:0] u_csamul_cska32_fa9_5_or0;
  wire [0:0] u_csamul_cska32_and10_5;
  wire [0:0] u_csamul_cska32_fa10_5_xor1;
  wire [0:0] u_csamul_cska32_fa10_5_or0;
  wire [0:0] u_csamul_cska32_and11_5;
  wire [0:0] u_csamul_cska32_fa11_5_xor1;
  wire [0:0] u_csamul_cska32_fa11_5_or0;
  wire [0:0] u_csamul_cska32_and12_5;
  wire [0:0] u_csamul_cska32_fa12_5_xor1;
  wire [0:0] u_csamul_cska32_fa12_5_or0;
  wire [0:0] u_csamul_cska32_and13_5;
  wire [0:0] u_csamul_cska32_fa13_5_xor1;
  wire [0:0] u_csamul_cska32_fa13_5_or0;
  wire [0:0] u_csamul_cska32_and14_5;
  wire [0:0] u_csamul_cska32_fa14_5_xor1;
  wire [0:0] u_csamul_cska32_fa14_5_or0;
  wire [0:0] u_csamul_cska32_and15_5;
  wire [0:0] u_csamul_cska32_fa15_5_xor1;
  wire [0:0] u_csamul_cska32_fa15_5_or0;
  wire [0:0] u_csamul_cska32_and16_5;
  wire [0:0] u_csamul_cska32_fa16_5_xor1;
  wire [0:0] u_csamul_cska32_fa16_5_or0;
  wire [0:0] u_csamul_cska32_and17_5;
  wire [0:0] u_csamul_cska32_fa17_5_xor1;
  wire [0:0] u_csamul_cska32_fa17_5_or0;
  wire [0:0] u_csamul_cska32_and18_5;
  wire [0:0] u_csamul_cska32_fa18_5_xor1;
  wire [0:0] u_csamul_cska32_fa18_5_or0;
  wire [0:0] u_csamul_cska32_and19_5;
  wire [0:0] u_csamul_cska32_fa19_5_xor1;
  wire [0:0] u_csamul_cska32_fa19_5_or0;
  wire [0:0] u_csamul_cska32_and20_5;
  wire [0:0] u_csamul_cska32_fa20_5_xor1;
  wire [0:0] u_csamul_cska32_fa20_5_or0;
  wire [0:0] u_csamul_cska32_and21_5;
  wire [0:0] u_csamul_cska32_fa21_5_xor1;
  wire [0:0] u_csamul_cska32_fa21_5_or0;
  wire [0:0] u_csamul_cska32_and22_5;
  wire [0:0] u_csamul_cska32_fa22_5_xor1;
  wire [0:0] u_csamul_cska32_fa22_5_or0;
  wire [0:0] u_csamul_cska32_and23_5;
  wire [0:0] u_csamul_cska32_fa23_5_xor1;
  wire [0:0] u_csamul_cska32_fa23_5_or0;
  wire [0:0] u_csamul_cska32_and24_5;
  wire [0:0] u_csamul_cska32_fa24_5_xor1;
  wire [0:0] u_csamul_cska32_fa24_5_or0;
  wire [0:0] u_csamul_cska32_and25_5;
  wire [0:0] u_csamul_cska32_fa25_5_xor1;
  wire [0:0] u_csamul_cska32_fa25_5_or0;
  wire [0:0] u_csamul_cska32_and26_5;
  wire [0:0] u_csamul_cska32_fa26_5_xor1;
  wire [0:0] u_csamul_cska32_fa26_5_or0;
  wire [0:0] u_csamul_cska32_and27_5;
  wire [0:0] u_csamul_cska32_fa27_5_xor1;
  wire [0:0] u_csamul_cska32_fa27_5_or0;
  wire [0:0] u_csamul_cska32_and28_5;
  wire [0:0] u_csamul_cska32_fa28_5_xor1;
  wire [0:0] u_csamul_cska32_fa28_5_or0;
  wire [0:0] u_csamul_cska32_and29_5;
  wire [0:0] u_csamul_cska32_fa29_5_xor1;
  wire [0:0] u_csamul_cska32_fa29_5_or0;
  wire [0:0] u_csamul_cska32_and30_5;
  wire [0:0] u_csamul_cska32_fa30_5_xor1;
  wire [0:0] u_csamul_cska32_fa30_5_or0;
  wire [0:0] u_csamul_cska32_and31_5;
  wire [0:0] u_csamul_cska32_and0_6;
  wire [0:0] u_csamul_cska32_fa0_6_xor1;
  wire [0:0] u_csamul_cska32_fa0_6_or0;
  wire [0:0] u_csamul_cska32_and1_6;
  wire [0:0] u_csamul_cska32_fa1_6_xor1;
  wire [0:0] u_csamul_cska32_fa1_6_or0;
  wire [0:0] u_csamul_cska32_and2_6;
  wire [0:0] u_csamul_cska32_fa2_6_xor1;
  wire [0:0] u_csamul_cska32_fa2_6_or0;
  wire [0:0] u_csamul_cska32_and3_6;
  wire [0:0] u_csamul_cska32_fa3_6_xor1;
  wire [0:0] u_csamul_cska32_fa3_6_or0;
  wire [0:0] u_csamul_cska32_and4_6;
  wire [0:0] u_csamul_cska32_fa4_6_xor1;
  wire [0:0] u_csamul_cska32_fa4_6_or0;
  wire [0:0] u_csamul_cska32_and5_6;
  wire [0:0] u_csamul_cska32_fa5_6_xor1;
  wire [0:0] u_csamul_cska32_fa5_6_or0;
  wire [0:0] u_csamul_cska32_and6_6;
  wire [0:0] u_csamul_cska32_fa6_6_xor1;
  wire [0:0] u_csamul_cska32_fa6_6_or0;
  wire [0:0] u_csamul_cska32_and7_6;
  wire [0:0] u_csamul_cska32_fa7_6_xor1;
  wire [0:0] u_csamul_cska32_fa7_6_or0;
  wire [0:0] u_csamul_cska32_and8_6;
  wire [0:0] u_csamul_cska32_fa8_6_xor1;
  wire [0:0] u_csamul_cska32_fa8_6_or0;
  wire [0:0] u_csamul_cska32_and9_6;
  wire [0:0] u_csamul_cska32_fa9_6_xor1;
  wire [0:0] u_csamul_cska32_fa9_6_or0;
  wire [0:0] u_csamul_cska32_and10_6;
  wire [0:0] u_csamul_cska32_fa10_6_xor1;
  wire [0:0] u_csamul_cska32_fa10_6_or0;
  wire [0:0] u_csamul_cska32_and11_6;
  wire [0:0] u_csamul_cska32_fa11_6_xor1;
  wire [0:0] u_csamul_cska32_fa11_6_or0;
  wire [0:0] u_csamul_cska32_and12_6;
  wire [0:0] u_csamul_cska32_fa12_6_xor1;
  wire [0:0] u_csamul_cska32_fa12_6_or0;
  wire [0:0] u_csamul_cska32_and13_6;
  wire [0:0] u_csamul_cska32_fa13_6_xor1;
  wire [0:0] u_csamul_cska32_fa13_6_or0;
  wire [0:0] u_csamul_cska32_and14_6;
  wire [0:0] u_csamul_cska32_fa14_6_xor1;
  wire [0:0] u_csamul_cska32_fa14_6_or0;
  wire [0:0] u_csamul_cska32_and15_6;
  wire [0:0] u_csamul_cska32_fa15_6_xor1;
  wire [0:0] u_csamul_cska32_fa15_6_or0;
  wire [0:0] u_csamul_cska32_and16_6;
  wire [0:0] u_csamul_cska32_fa16_6_xor1;
  wire [0:0] u_csamul_cska32_fa16_6_or0;
  wire [0:0] u_csamul_cska32_and17_6;
  wire [0:0] u_csamul_cska32_fa17_6_xor1;
  wire [0:0] u_csamul_cska32_fa17_6_or0;
  wire [0:0] u_csamul_cska32_and18_6;
  wire [0:0] u_csamul_cska32_fa18_6_xor1;
  wire [0:0] u_csamul_cska32_fa18_6_or0;
  wire [0:0] u_csamul_cska32_and19_6;
  wire [0:0] u_csamul_cska32_fa19_6_xor1;
  wire [0:0] u_csamul_cska32_fa19_6_or0;
  wire [0:0] u_csamul_cska32_and20_6;
  wire [0:0] u_csamul_cska32_fa20_6_xor1;
  wire [0:0] u_csamul_cska32_fa20_6_or0;
  wire [0:0] u_csamul_cska32_and21_6;
  wire [0:0] u_csamul_cska32_fa21_6_xor1;
  wire [0:0] u_csamul_cska32_fa21_6_or0;
  wire [0:0] u_csamul_cska32_and22_6;
  wire [0:0] u_csamul_cska32_fa22_6_xor1;
  wire [0:0] u_csamul_cska32_fa22_6_or0;
  wire [0:0] u_csamul_cska32_and23_6;
  wire [0:0] u_csamul_cska32_fa23_6_xor1;
  wire [0:0] u_csamul_cska32_fa23_6_or0;
  wire [0:0] u_csamul_cska32_and24_6;
  wire [0:0] u_csamul_cska32_fa24_6_xor1;
  wire [0:0] u_csamul_cska32_fa24_6_or0;
  wire [0:0] u_csamul_cska32_and25_6;
  wire [0:0] u_csamul_cska32_fa25_6_xor1;
  wire [0:0] u_csamul_cska32_fa25_6_or0;
  wire [0:0] u_csamul_cska32_and26_6;
  wire [0:0] u_csamul_cska32_fa26_6_xor1;
  wire [0:0] u_csamul_cska32_fa26_6_or0;
  wire [0:0] u_csamul_cska32_and27_6;
  wire [0:0] u_csamul_cska32_fa27_6_xor1;
  wire [0:0] u_csamul_cska32_fa27_6_or0;
  wire [0:0] u_csamul_cska32_and28_6;
  wire [0:0] u_csamul_cska32_fa28_6_xor1;
  wire [0:0] u_csamul_cska32_fa28_6_or0;
  wire [0:0] u_csamul_cska32_and29_6;
  wire [0:0] u_csamul_cska32_fa29_6_xor1;
  wire [0:0] u_csamul_cska32_fa29_6_or0;
  wire [0:0] u_csamul_cska32_and30_6;
  wire [0:0] u_csamul_cska32_fa30_6_xor1;
  wire [0:0] u_csamul_cska32_fa30_6_or0;
  wire [0:0] u_csamul_cska32_and31_6;
  wire [0:0] u_csamul_cska32_and0_7;
  wire [0:0] u_csamul_cska32_fa0_7_xor1;
  wire [0:0] u_csamul_cska32_fa0_7_or0;
  wire [0:0] u_csamul_cska32_and1_7;
  wire [0:0] u_csamul_cska32_fa1_7_xor1;
  wire [0:0] u_csamul_cska32_fa1_7_or0;
  wire [0:0] u_csamul_cska32_and2_7;
  wire [0:0] u_csamul_cska32_fa2_7_xor1;
  wire [0:0] u_csamul_cska32_fa2_7_or0;
  wire [0:0] u_csamul_cska32_and3_7;
  wire [0:0] u_csamul_cska32_fa3_7_xor1;
  wire [0:0] u_csamul_cska32_fa3_7_or0;
  wire [0:0] u_csamul_cska32_and4_7;
  wire [0:0] u_csamul_cska32_fa4_7_xor1;
  wire [0:0] u_csamul_cska32_fa4_7_or0;
  wire [0:0] u_csamul_cska32_and5_7;
  wire [0:0] u_csamul_cska32_fa5_7_xor1;
  wire [0:0] u_csamul_cska32_fa5_7_or0;
  wire [0:0] u_csamul_cska32_and6_7;
  wire [0:0] u_csamul_cska32_fa6_7_xor1;
  wire [0:0] u_csamul_cska32_fa6_7_or0;
  wire [0:0] u_csamul_cska32_and7_7;
  wire [0:0] u_csamul_cska32_fa7_7_xor1;
  wire [0:0] u_csamul_cska32_fa7_7_or0;
  wire [0:0] u_csamul_cska32_and8_7;
  wire [0:0] u_csamul_cska32_fa8_7_xor1;
  wire [0:0] u_csamul_cska32_fa8_7_or0;
  wire [0:0] u_csamul_cska32_and9_7;
  wire [0:0] u_csamul_cska32_fa9_7_xor1;
  wire [0:0] u_csamul_cska32_fa9_7_or0;
  wire [0:0] u_csamul_cska32_and10_7;
  wire [0:0] u_csamul_cska32_fa10_7_xor1;
  wire [0:0] u_csamul_cska32_fa10_7_or0;
  wire [0:0] u_csamul_cska32_and11_7;
  wire [0:0] u_csamul_cska32_fa11_7_xor1;
  wire [0:0] u_csamul_cska32_fa11_7_or0;
  wire [0:0] u_csamul_cska32_and12_7;
  wire [0:0] u_csamul_cska32_fa12_7_xor1;
  wire [0:0] u_csamul_cska32_fa12_7_or0;
  wire [0:0] u_csamul_cska32_and13_7;
  wire [0:0] u_csamul_cska32_fa13_7_xor1;
  wire [0:0] u_csamul_cska32_fa13_7_or0;
  wire [0:0] u_csamul_cska32_and14_7;
  wire [0:0] u_csamul_cska32_fa14_7_xor1;
  wire [0:0] u_csamul_cska32_fa14_7_or0;
  wire [0:0] u_csamul_cska32_and15_7;
  wire [0:0] u_csamul_cska32_fa15_7_xor1;
  wire [0:0] u_csamul_cska32_fa15_7_or0;
  wire [0:0] u_csamul_cska32_and16_7;
  wire [0:0] u_csamul_cska32_fa16_7_xor1;
  wire [0:0] u_csamul_cska32_fa16_7_or0;
  wire [0:0] u_csamul_cska32_and17_7;
  wire [0:0] u_csamul_cska32_fa17_7_xor1;
  wire [0:0] u_csamul_cska32_fa17_7_or0;
  wire [0:0] u_csamul_cska32_and18_7;
  wire [0:0] u_csamul_cska32_fa18_7_xor1;
  wire [0:0] u_csamul_cska32_fa18_7_or0;
  wire [0:0] u_csamul_cska32_and19_7;
  wire [0:0] u_csamul_cska32_fa19_7_xor1;
  wire [0:0] u_csamul_cska32_fa19_7_or0;
  wire [0:0] u_csamul_cska32_and20_7;
  wire [0:0] u_csamul_cska32_fa20_7_xor1;
  wire [0:0] u_csamul_cska32_fa20_7_or0;
  wire [0:0] u_csamul_cska32_and21_7;
  wire [0:0] u_csamul_cska32_fa21_7_xor1;
  wire [0:0] u_csamul_cska32_fa21_7_or0;
  wire [0:0] u_csamul_cska32_and22_7;
  wire [0:0] u_csamul_cska32_fa22_7_xor1;
  wire [0:0] u_csamul_cska32_fa22_7_or0;
  wire [0:0] u_csamul_cska32_and23_7;
  wire [0:0] u_csamul_cska32_fa23_7_xor1;
  wire [0:0] u_csamul_cska32_fa23_7_or0;
  wire [0:0] u_csamul_cska32_and24_7;
  wire [0:0] u_csamul_cska32_fa24_7_xor1;
  wire [0:0] u_csamul_cska32_fa24_7_or0;
  wire [0:0] u_csamul_cska32_and25_7;
  wire [0:0] u_csamul_cska32_fa25_7_xor1;
  wire [0:0] u_csamul_cska32_fa25_7_or0;
  wire [0:0] u_csamul_cska32_and26_7;
  wire [0:0] u_csamul_cska32_fa26_7_xor1;
  wire [0:0] u_csamul_cska32_fa26_7_or0;
  wire [0:0] u_csamul_cska32_and27_7;
  wire [0:0] u_csamul_cska32_fa27_7_xor1;
  wire [0:0] u_csamul_cska32_fa27_7_or0;
  wire [0:0] u_csamul_cska32_and28_7;
  wire [0:0] u_csamul_cska32_fa28_7_xor1;
  wire [0:0] u_csamul_cska32_fa28_7_or0;
  wire [0:0] u_csamul_cska32_and29_7;
  wire [0:0] u_csamul_cska32_fa29_7_xor1;
  wire [0:0] u_csamul_cska32_fa29_7_or0;
  wire [0:0] u_csamul_cska32_and30_7;
  wire [0:0] u_csamul_cska32_fa30_7_xor1;
  wire [0:0] u_csamul_cska32_fa30_7_or0;
  wire [0:0] u_csamul_cska32_and31_7;
  wire [0:0] u_csamul_cska32_and0_8;
  wire [0:0] u_csamul_cska32_fa0_8_xor1;
  wire [0:0] u_csamul_cska32_fa0_8_or0;
  wire [0:0] u_csamul_cska32_and1_8;
  wire [0:0] u_csamul_cska32_fa1_8_xor1;
  wire [0:0] u_csamul_cska32_fa1_8_or0;
  wire [0:0] u_csamul_cska32_and2_8;
  wire [0:0] u_csamul_cska32_fa2_8_xor1;
  wire [0:0] u_csamul_cska32_fa2_8_or0;
  wire [0:0] u_csamul_cska32_and3_8;
  wire [0:0] u_csamul_cska32_fa3_8_xor1;
  wire [0:0] u_csamul_cska32_fa3_8_or0;
  wire [0:0] u_csamul_cska32_and4_8;
  wire [0:0] u_csamul_cska32_fa4_8_xor1;
  wire [0:0] u_csamul_cska32_fa4_8_or0;
  wire [0:0] u_csamul_cska32_and5_8;
  wire [0:0] u_csamul_cska32_fa5_8_xor1;
  wire [0:0] u_csamul_cska32_fa5_8_or0;
  wire [0:0] u_csamul_cska32_and6_8;
  wire [0:0] u_csamul_cska32_fa6_8_xor1;
  wire [0:0] u_csamul_cska32_fa6_8_or0;
  wire [0:0] u_csamul_cska32_and7_8;
  wire [0:0] u_csamul_cska32_fa7_8_xor1;
  wire [0:0] u_csamul_cska32_fa7_8_or0;
  wire [0:0] u_csamul_cska32_and8_8;
  wire [0:0] u_csamul_cska32_fa8_8_xor1;
  wire [0:0] u_csamul_cska32_fa8_8_or0;
  wire [0:0] u_csamul_cska32_and9_8;
  wire [0:0] u_csamul_cska32_fa9_8_xor1;
  wire [0:0] u_csamul_cska32_fa9_8_or0;
  wire [0:0] u_csamul_cska32_and10_8;
  wire [0:0] u_csamul_cska32_fa10_8_xor1;
  wire [0:0] u_csamul_cska32_fa10_8_or0;
  wire [0:0] u_csamul_cska32_and11_8;
  wire [0:0] u_csamul_cska32_fa11_8_xor1;
  wire [0:0] u_csamul_cska32_fa11_8_or0;
  wire [0:0] u_csamul_cska32_and12_8;
  wire [0:0] u_csamul_cska32_fa12_8_xor1;
  wire [0:0] u_csamul_cska32_fa12_8_or0;
  wire [0:0] u_csamul_cska32_and13_8;
  wire [0:0] u_csamul_cska32_fa13_8_xor1;
  wire [0:0] u_csamul_cska32_fa13_8_or0;
  wire [0:0] u_csamul_cska32_and14_8;
  wire [0:0] u_csamul_cska32_fa14_8_xor1;
  wire [0:0] u_csamul_cska32_fa14_8_or0;
  wire [0:0] u_csamul_cska32_and15_8;
  wire [0:0] u_csamul_cska32_fa15_8_xor1;
  wire [0:0] u_csamul_cska32_fa15_8_or0;
  wire [0:0] u_csamul_cska32_and16_8;
  wire [0:0] u_csamul_cska32_fa16_8_xor1;
  wire [0:0] u_csamul_cska32_fa16_8_or0;
  wire [0:0] u_csamul_cska32_and17_8;
  wire [0:0] u_csamul_cska32_fa17_8_xor1;
  wire [0:0] u_csamul_cska32_fa17_8_or0;
  wire [0:0] u_csamul_cska32_and18_8;
  wire [0:0] u_csamul_cska32_fa18_8_xor1;
  wire [0:0] u_csamul_cska32_fa18_8_or0;
  wire [0:0] u_csamul_cska32_and19_8;
  wire [0:0] u_csamul_cska32_fa19_8_xor1;
  wire [0:0] u_csamul_cska32_fa19_8_or0;
  wire [0:0] u_csamul_cska32_and20_8;
  wire [0:0] u_csamul_cska32_fa20_8_xor1;
  wire [0:0] u_csamul_cska32_fa20_8_or0;
  wire [0:0] u_csamul_cska32_and21_8;
  wire [0:0] u_csamul_cska32_fa21_8_xor1;
  wire [0:0] u_csamul_cska32_fa21_8_or0;
  wire [0:0] u_csamul_cska32_and22_8;
  wire [0:0] u_csamul_cska32_fa22_8_xor1;
  wire [0:0] u_csamul_cska32_fa22_8_or0;
  wire [0:0] u_csamul_cska32_and23_8;
  wire [0:0] u_csamul_cska32_fa23_8_xor1;
  wire [0:0] u_csamul_cska32_fa23_8_or0;
  wire [0:0] u_csamul_cska32_and24_8;
  wire [0:0] u_csamul_cska32_fa24_8_xor1;
  wire [0:0] u_csamul_cska32_fa24_8_or0;
  wire [0:0] u_csamul_cska32_and25_8;
  wire [0:0] u_csamul_cska32_fa25_8_xor1;
  wire [0:0] u_csamul_cska32_fa25_8_or0;
  wire [0:0] u_csamul_cska32_and26_8;
  wire [0:0] u_csamul_cska32_fa26_8_xor1;
  wire [0:0] u_csamul_cska32_fa26_8_or0;
  wire [0:0] u_csamul_cska32_and27_8;
  wire [0:0] u_csamul_cska32_fa27_8_xor1;
  wire [0:0] u_csamul_cska32_fa27_8_or0;
  wire [0:0] u_csamul_cska32_and28_8;
  wire [0:0] u_csamul_cska32_fa28_8_xor1;
  wire [0:0] u_csamul_cska32_fa28_8_or0;
  wire [0:0] u_csamul_cska32_and29_8;
  wire [0:0] u_csamul_cska32_fa29_8_xor1;
  wire [0:0] u_csamul_cska32_fa29_8_or0;
  wire [0:0] u_csamul_cska32_and30_8;
  wire [0:0] u_csamul_cska32_fa30_8_xor1;
  wire [0:0] u_csamul_cska32_fa30_8_or0;
  wire [0:0] u_csamul_cska32_and31_8;
  wire [0:0] u_csamul_cska32_and0_9;
  wire [0:0] u_csamul_cska32_fa0_9_xor1;
  wire [0:0] u_csamul_cska32_fa0_9_or0;
  wire [0:0] u_csamul_cska32_and1_9;
  wire [0:0] u_csamul_cska32_fa1_9_xor1;
  wire [0:0] u_csamul_cska32_fa1_9_or0;
  wire [0:0] u_csamul_cska32_and2_9;
  wire [0:0] u_csamul_cska32_fa2_9_xor1;
  wire [0:0] u_csamul_cska32_fa2_9_or0;
  wire [0:0] u_csamul_cska32_and3_9;
  wire [0:0] u_csamul_cska32_fa3_9_xor1;
  wire [0:0] u_csamul_cska32_fa3_9_or0;
  wire [0:0] u_csamul_cska32_and4_9;
  wire [0:0] u_csamul_cska32_fa4_9_xor1;
  wire [0:0] u_csamul_cska32_fa4_9_or0;
  wire [0:0] u_csamul_cska32_and5_9;
  wire [0:0] u_csamul_cska32_fa5_9_xor1;
  wire [0:0] u_csamul_cska32_fa5_9_or0;
  wire [0:0] u_csamul_cska32_and6_9;
  wire [0:0] u_csamul_cska32_fa6_9_xor1;
  wire [0:0] u_csamul_cska32_fa6_9_or0;
  wire [0:0] u_csamul_cska32_and7_9;
  wire [0:0] u_csamul_cska32_fa7_9_xor1;
  wire [0:0] u_csamul_cska32_fa7_9_or0;
  wire [0:0] u_csamul_cska32_and8_9;
  wire [0:0] u_csamul_cska32_fa8_9_xor1;
  wire [0:0] u_csamul_cska32_fa8_9_or0;
  wire [0:0] u_csamul_cska32_and9_9;
  wire [0:0] u_csamul_cska32_fa9_9_xor1;
  wire [0:0] u_csamul_cska32_fa9_9_or0;
  wire [0:0] u_csamul_cska32_and10_9;
  wire [0:0] u_csamul_cska32_fa10_9_xor1;
  wire [0:0] u_csamul_cska32_fa10_9_or0;
  wire [0:0] u_csamul_cska32_and11_9;
  wire [0:0] u_csamul_cska32_fa11_9_xor1;
  wire [0:0] u_csamul_cska32_fa11_9_or0;
  wire [0:0] u_csamul_cska32_and12_9;
  wire [0:0] u_csamul_cska32_fa12_9_xor1;
  wire [0:0] u_csamul_cska32_fa12_9_or0;
  wire [0:0] u_csamul_cska32_and13_9;
  wire [0:0] u_csamul_cska32_fa13_9_xor1;
  wire [0:0] u_csamul_cska32_fa13_9_or0;
  wire [0:0] u_csamul_cska32_and14_9;
  wire [0:0] u_csamul_cska32_fa14_9_xor1;
  wire [0:0] u_csamul_cska32_fa14_9_or0;
  wire [0:0] u_csamul_cska32_and15_9;
  wire [0:0] u_csamul_cska32_fa15_9_xor1;
  wire [0:0] u_csamul_cska32_fa15_9_or0;
  wire [0:0] u_csamul_cska32_and16_9;
  wire [0:0] u_csamul_cska32_fa16_9_xor1;
  wire [0:0] u_csamul_cska32_fa16_9_or0;
  wire [0:0] u_csamul_cska32_and17_9;
  wire [0:0] u_csamul_cska32_fa17_9_xor1;
  wire [0:0] u_csamul_cska32_fa17_9_or0;
  wire [0:0] u_csamul_cska32_and18_9;
  wire [0:0] u_csamul_cska32_fa18_9_xor1;
  wire [0:0] u_csamul_cska32_fa18_9_or0;
  wire [0:0] u_csamul_cska32_and19_9;
  wire [0:0] u_csamul_cska32_fa19_9_xor1;
  wire [0:0] u_csamul_cska32_fa19_9_or0;
  wire [0:0] u_csamul_cska32_and20_9;
  wire [0:0] u_csamul_cska32_fa20_9_xor1;
  wire [0:0] u_csamul_cska32_fa20_9_or0;
  wire [0:0] u_csamul_cska32_and21_9;
  wire [0:0] u_csamul_cska32_fa21_9_xor1;
  wire [0:0] u_csamul_cska32_fa21_9_or0;
  wire [0:0] u_csamul_cska32_and22_9;
  wire [0:0] u_csamul_cska32_fa22_9_xor1;
  wire [0:0] u_csamul_cska32_fa22_9_or0;
  wire [0:0] u_csamul_cska32_and23_9;
  wire [0:0] u_csamul_cska32_fa23_9_xor1;
  wire [0:0] u_csamul_cska32_fa23_9_or0;
  wire [0:0] u_csamul_cska32_and24_9;
  wire [0:0] u_csamul_cska32_fa24_9_xor1;
  wire [0:0] u_csamul_cska32_fa24_9_or0;
  wire [0:0] u_csamul_cska32_and25_9;
  wire [0:0] u_csamul_cska32_fa25_9_xor1;
  wire [0:0] u_csamul_cska32_fa25_9_or0;
  wire [0:0] u_csamul_cska32_and26_9;
  wire [0:0] u_csamul_cska32_fa26_9_xor1;
  wire [0:0] u_csamul_cska32_fa26_9_or0;
  wire [0:0] u_csamul_cska32_and27_9;
  wire [0:0] u_csamul_cska32_fa27_9_xor1;
  wire [0:0] u_csamul_cska32_fa27_9_or0;
  wire [0:0] u_csamul_cska32_and28_9;
  wire [0:0] u_csamul_cska32_fa28_9_xor1;
  wire [0:0] u_csamul_cska32_fa28_9_or0;
  wire [0:0] u_csamul_cska32_and29_9;
  wire [0:0] u_csamul_cska32_fa29_9_xor1;
  wire [0:0] u_csamul_cska32_fa29_9_or0;
  wire [0:0] u_csamul_cska32_and30_9;
  wire [0:0] u_csamul_cska32_fa30_9_xor1;
  wire [0:0] u_csamul_cska32_fa30_9_or0;
  wire [0:0] u_csamul_cska32_and31_9;
  wire [0:0] u_csamul_cska32_and0_10;
  wire [0:0] u_csamul_cska32_fa0_10_xor1;
  wire [0:0] u_csamul_cska32_fa0_10_or0;
  wire [0:0] u_csamul_cska32_and1_10;
  wire [0:0] u_csamul_cska32_fa1_10_xor1;
  wire [0:0] u_csamul_cska32_fa1_10_or0;
  wire [0:0] u_csamul_cska32_and2_10;
  wire [0:0] u_csamul_cska32_fa2_10_xor1;
  wire [0:0] u_csamul_cska32_fa2_10_or0;
  wire [0:0] u_csamul_cska32_and3_10;
  wire [0:0] u_csamul_cska32_fa3_10_xor1;
  wire [0:0] u_csamul_cska32_fa3_10_or0;
  wire [0:0] u_csamul_cska32_and4_10;
  wire [0:0] u_csamul_cska32_fa4_10_xor1;
  wire [0:0] u_csamul_cska32_fa4_10_or0;
  wire [0:0] u_csamul_cska32_and5_10;
  wire [0:0] u_csamul_cska32_fa5_10_xor1;
  wire [0:0] u_csamul_cska32_fa5_10_or0;
  wire [0:0] u_csamul_cska32_and6_10;
  wire [0:0] u_csamul_cska32_fa6_10_xor1;
  wire [0:0] u_csamul_cska32_fa6_10_or0;
  wire [0:0] u_csamul_cska32_and7_10;
  wire [0:0] u_csamul_cska32_fa7_10_xor1;
  wire [0:0] u_csamul_cska32_fa7_10_or0;
  wire [0:0] u_csamul_cska32_and8_10;
  wire [0:0] u_csamul_cska32_fa8_10_xor1;
  wire [0:0] u_csamul_cska32_fa8_10_or0;
  wire [0:0] u_csamul_cska32_and9_10;
  wire [0:0] u_csamul_cska32_fa9_10_xor1;
  wire [0:0] u_csamul_cska32_fa9_10_or0;
  wire [0:0] u_csamul_cska32_and10_10;
  wire [0:0] u_csamul_cska32_fa10_10_xor1;
  wire [0:0] u_csamul_cska32_fa10_10_or0;
  wire [0:0] u_csamul_cska32_and11_10;
  wire [0:0] u_csamul_cska32_fa11_10_xor1;
  wire [0:0] u_csamul_cska32_fa11_10_or0;
  wire [0:0] u_csamul_cska32_and12_10;
  wire [0:0] u_csamul_cska32_fa12_10_xor1;
  wire [0:0] u_csamul_cska32_fa12_10_or0;
  wire [0:0] u_csamul_cska32_and13_10;
  wire [0:0] u_csamul_cska32_fa13_10_xor1;
  wire [0:0] u_csamul_cska32_fa13_10_or0;
  wire [0:0] u_csamul_cska32_and14_10;
  wire [0:0] u_csamul_cska32_fa14_10_xor1;
  wire [0:0] u_csamul_cska32_fa14_10_or0;
  wire [0:0] u_csamul_cska32_and15_10;
  wire [0:0] u_csamul_cska32_fa15_10_xor1;
  wire [0:0] u_csamul_cska32_fa15_10_or0;
  wire [0:0] u_csamul_cska32_and16_10;
  wire [0:0] u_csamul_cska32_fa16_10_xor1;
  wire [0:0] u_csamul_cska32_fa16_10_or0;
  wire [0:0] u_csamul_cska32_and17_10;
  wire [0:0] u_csamul_cska32_fa17_10_xor1;
  wire [0:0] u_csamul_cska32_fa17_10_or0;
  wire [0:0] u_csamul_cska32_and18_10;
  wire [0:0] u_csamul_cska32_fa18_10_xor1;
  wire [0:0] u_csamul_cska32_fa18_10_or0;
  wire [0:0] u_csamul_cska32_and19_10;
  wire [0:0] u_csamul_cska32_fa19_10_xor1;
  wire [0:0] u_csamul_cska32_fa19_10_or0;
  wire [0:0] u_csamul_cska32_and20_10;
  wire [0:0] u_csamul_cska32_fa20_10_xor1;
  wire [0:0] u_csamul_cska32_fa20_10_or0;
  wire [0:0] u_csamul_cska32_and21_10;
  wire [0:0] u_csamul_cska32_fa21_10_xor1;
  wire [0:0] u_csamul_cska32_fa21_10_or0;
  wire [0:0] u_csamul_cska32_and22_10;
  wire [0:0] u_csamul_cska32_fa22_10_xor1;
  wire [0:0] u_csamul_cska32_fa22_10_or0;
  wire [0:0] u_csamul_cska32_and23_10;
  wire [0:0] u_csamul_cska32_fa23_10_xor1;
  wire [0:0] u_csamul_cska32_fa23_10_or0;
  wire [0:0] u_csamul_cska32_and24_10;
  wire [0:0] u_csamul_cska32_fa24_10_xor1;
  wire [0:0] u_csamul_cska32_fa24_10_or0;
  wire [0:0] u_csamul_cska32_and25_10;
  wire [0:0] u_csamul_cska32_fa25_10_xor1;
  wire [0:0] u_csamul_cska32_fa25_10_or0;
  wire [0:0] u_csamul_cska32_and26_10;
  wire [0:0] u_csamul_cska32_fa26_10_xor1;
  wire [0:0] u_csamul_cska32_fa26_10_or0;
  wire [0:0] u_csamul_cska32_and27_10;
  wire [0:0] u_csamul_cska32_fa27_10_xor1;
  wire [0:0] u_csamul_cska32_fa27_10_or0;
  wire [0:0] u_csamul_cska32_and28_10;
  wire [0:0] u_csamul_cska32_fa28_10_xor1;
  wire [0:0] u_csamul_cska32_fa28_10_or0;
  wire [0:0] u_csamul_cska32_and29_10;
  wire [0:0] u_csamul_cska32_fa29_10_xor1;
  wire [0:0] u_csamul_cska32_fa29_10_or0;
  wire [0:0] u_csamul_cska32_and30_10;
  wire [0:0] u_csamul_cska32_fa30_10_xor1;
  wire [0:0] u_csamul_cska32_fa30_10_or0;
  wire [0:0] u_csamul_cska32_and31_10;
  wire [0:0] u_csamul_cska32_and0_11;
  wire [0:0] u_csamul_cska32_fa0_11_xor1;
  wire [0:0] u_csamul_cska32_fa0_11_or0;
  wire [0:0] u_csamul_cska32_and1_11;
  wire [0:0] u_csamul_cska32_fa1_11_xor1;
  wire [0:0] u_csamul_cska32_fa1_11_or0;
  wire [0:0] u_csamul_cska32_and2_11;
  wire [0:0] u_csamul_cska32_fa2_11_xor1;
  wire [0:0] u_csamul_cska32_fa2_11_or0;
  wire [0:0] u_csamul_cska32_and3_11;
  wire [0:0] u_csamul_cska32_fa3_11_xor1;
  wire [0:0] u_csamul_cska32_fa3_11_or0;
  wire [0:0] u_csamul_cska32_and4_11;
  wire [0:0] u_csamul_cska32_fa4_11_xor1;
  wire [0:0] u_csamul_cska32_fa4_11_or0;
  wire [0:0] u_csamul_cska32_and5_11;
  wire [0:0] u_csamul_cska32_fa5_11_xor1;
  wire [0:0] u_csamul_cska32_fa5_11_or0;
  wire [0:0] u_csamul_cska32_and6_11;
  wire [0:0] u_csamul_cska32_fa6_11_xor1;
  wire [0:0] u_csamul_cska32_fa6_11_or0;
  wire [0:0] u_csamul_cska32_and7_11;
  wire [0:0] u_csamul_cska32_fa7_11_xor1;
  wire [0:0] u_csamul_cska32_fa7_11_or0;
  wire [0:0] u_csamul_cska32_and8_11;
  wire [0:0] u_csamul_cska32_fa8_11_xor1;
  wire [0:0] u_csamul_cska32_fa8_11_or0;
  wire [0:0] u_csamul_cska32_and9_11;
  wire [0:0] u_csamul_cska32_fa9_11_xor1;
  wire [0:0] u_csamul_cska32_fa9_11_or0;
  wire [0:0] u_csamul_cska32_and10_11;
  wire [0:0] u_csamul_cska32_fa10_11_xor1;
  wire [0:0] u_csamul_cska32_fa10_11_or0;
  wire [0:0] u_csamul_cska32_and11_11;
  wire [0:0] u_csamul_cska32_fa11_11_xor1;
  wire [0:0] u_csamul_cska32_fa11_11_or0;
  wire [0:0] u_csamul_cska32_and12_11;
  wire [0:0] u_csamul_cska32_fa12_11_xor1;
  wire [0:0] u_csamul_cska32_fa12_11_or0;
  wire [0:0] u_csamul_cska32_and13_11;
  wire [0:0] u_csamul_cska32_fa13_11_xor1;
  wire [0:0] u_csamul_cska32_fa13_11_or0;
  wire [0:0] u_csamul_cska32_and14_11;
  wire [0:0] u_csamul_cska32_fa14_11_xor1;
  wire [0:0] u_csamul_cska32_fa14_11_or0;
  wire [0:0] u_csamul_cska32_and15_11;
  wire [0:0] u_csamul_cska32_fa15_11_xor1;
  wire [0:0] u_csamul_cska32_fa15_11_or0;
  wire [0:0] u_csamul_cska32_and16_11;
  wire [0:0] u_csamul_cska32_fa16_11_xor1;
  wire [0:0] u_csamul_cska32_fa16_11_or0;
  wire [0:0] u_csamul_cska32_and17_11;
  wire [0:0] u_csamul_cska32_fa17_11_xor1;
  wire [0:0] u_csamul_cska32_fa17_11_or0;
  wire [0:0] u_csamul_cska32_and18_11;
  wire [0:0] u_csamul_cska32_fa18_11_xor1;
  wire [0:0] u_csamul_cska32_fa18_11_or0;
  wire [0:0] u_csamul_cska32_and19_11;
  wire [0:0] u_csamul_cska32_fa19_11_xor1;
  wire [0:0] u_csamul_cska32_fa19_11_or0;
  wire [0:0] u_csamul_cska32_and20_11;
  wire [0:0] u_csamul_cska32_fa20_11_xor1;
  wire [0:0] u_csamul_cska32_fa20_11_or0;
  wire [0:0] u_csamul_cska32_and21_11;
  wire [0:0] u_csamul_cska32_fa21_11_xor1;
  wire [0:0] u_csamul_cska32_fa21_11_or0;
  wire [0:0] u_csamul_cska32_and22_11;
  wire [0:0] u_csamul_cska32_fa22_11_xor1;
  wire [0:0] u_csamul_cska32_fa22_11_or0;
  wire [0:0] u_csamul_cska32_and23_11;
  wire [0:0] u_csamul_cska32_fa23_11_xor1;
  wire [0:0] u_csamul_cska32_fa23_11_or0;
  wire [0:0] u_csamul_cska32_and24_11;
  wire [0:0] u_csamul_cska32_fa24_11_xor1;
  wire [0:0] u_csamul_cska32_fa24_11_or0;
  wire [0:0] u_csamul_cska32_and25_11;
  wire [0:0] u_csamul_cska32_fa25_11_xor1;
  wire [0:0] u_csamul_cska32_fa25_11_or0;
  wire [0:0] u_csamul_cska32_and26_11;
  wire [0:0] u_csamul_cska32_fa26_11_xor1;
  wire [0:0] u_csamul_cska32_fa26_11_or0;
  wire [0:0] u_csamul_cska32_and27_11;
  wire [0:0] u_csamul_cska32_fa27_11_xor1;
  wire [0:0] u_csamul_cska32_fa27_11_or0;
  wire [0:0] u_csamul_cska32_and28_11;
  wire [0:0] u_csamul_cska32_fa28_11_xor1;
  wire [0:0] u_csamul_cska32_fa28_11_or0;
  wire [0:0] u_csamul_cska32_and29_11;
  wire [0:0] u_csamul_cska32_fa29_11_xor1;
  wire [0:0] u_csamul_cska32_fa29_11_or0;
  wire [0:0] u_csamul_cska32_and30_11;
  wire [0:0] u_csamul_cska32_fa30_11_xor1;
  wire [0:0] u_csamul_cska32_fa30_11_or0;
  wire [0:0] u_csamul_cska32_and31_11;
  wire [0:0] u_csamul_cska32_and0_12;
  wire [0:0] u_csamul_cska32_fa0_12_xor1;
  wire [0:0] u_csamul_cska32_fa0_12_or0;
  wire [0:0] u_csamul_cska32_and1_12;
  wire [0:0] u_csamul_cska32_fa1_12_xor1;
  wire [0:0] u_csamul_cska32_fa1_12_or0;
  wire [0:0] u_csamul_cska32_and2_12;
  wire [0:0] u_csamul_cska32_fa2_12_xor1;
  wire [0:0] u_csamul_cska32_fa2_12_or0;
  wire [0:0] u_csamul_cska32_and3_12;
  wire [0:0] u_csamul_cska32_fa3_12_xor1;
  wire [0:0] u_csamul_cska32_fa3_12_or0;
  wire [0:0] u_csamul_cska32_and4_12;
  wire [0:0] u_csamul_cska32_fa4_12_xor1;
  wire [0:0] u_csamul_cska32_fa4_12_or0;
  wire [0:0] u_csamul_cska32_and5_12;
  wire [0:0] u_csamul_cska32_fa5_12_xor1;
  wire [0:0] u_csamul_cska32_fa5_12_or0;
  wire [0:0] u_csamul_cska32_and6_12;
  wire [0:0] u_csamul_cska32_fa6_12_xor1;
  wire [0:0] u_csamul_cska32_fa6_12_or0;
  wire [0:0] u_csamul_cska32_and7_12;
  wire [0:0] u_csamul_cska32_fa7_12_xor1;
  wire [0:0] u_csamul_cska32_fa7_12_or0;
  wire [0:0] u_csamul_cska32_and8_12;
  wire [0:0] u_csamul_cska32_fa8_12_xor1;
  wire [0:0] u_csamul_cska32_fa8_12_or0;
  wire [0:0] u_csamul_cska32_and9_12;
  wire [0:0] u_csamul_cska32_fa9_12_xor1;
  wire [0:0] u_csamul_cska32_fa9_12_or0;
  wire [0:0] u_csamul_cska32_and10_12;
  wire [0:0] u_csamul_cska32_fa10_12_xor1;
  wire [0:0] u_csamul_cska32_fa10_12_or0;
  wire [0:0] u_csamul_cska32_and11_12;
  wire [0:0] u_csamul_cska32_fa11_12_xor1;
  wire [0:0] u_csamul_cska32_fa11_12_or0;
  wire [0:0] u_csamul_cska32_and12_12;
  wire [0:0] u_csamul_cska32_fa12_12_xor1;
  wire [0:0] u_csamul_cska32_fa12_12_or0;
  wire [0:0] u_csamul_cska32_and13_12;
  wire [0:0] u_csamul_cska32_fa13_12_xor1;
  wire [0:0] u_csamul_cska32_fa13_12_or0;
  wire [0:0] u_csamul_cska32_and14_12;
  wire [0:0] u_csamul_cska32_fa14_12_xor1;
  wire [0:0] u_csamul_cska32_fa14_12_or0;
  wire [0:0] u_csamul_cska32_and15_12;
  wire [0:0] u_csamul_cska32_fa15_12_xor1;
  wire [0:0] u_csamul_cska32_fa15_12_or0;
  wire [0:0] u_csamul_cska32_and16_12;
  wire [0:0] u_csamul_cska32_fa16_12_xor1;
  wire [0:0] u_csamul_cska32_fa16_12_or0;
  wire [0:0] u_csamul_cska32_and17_12;
  wire [0:0] u_csamul_cska32_fa17_12_xor1;
  wire [0:0] u_csamul_cska32_fa17_12_or0;
  wire [0:0] u_csamul_cska32_and18_12;
  wire [0:0] u_csamul_cska32_fa18_12_xor1;
  wire [0:0] u_csamul_cska32_fa18_12_or0;
  wire [0:0] u_csamul_cska32_and19_12;
  wire [0:0] u_csamul_cska32_fa19_12_xor1;
  wire [0:0] u_csamul_cska32_fa19_12_or0;
  wire [0:0] u_csamul_cska32_and20_12;
  wire [0:0] u_csamul_cska32_fa20_12_xor1;
  wire [0:0] u_csamul_cska32_fa20_12_or0;
  wire [0:0] u_csamul_cska32_and21_12;
  wire [0:0] u_csamul_cska32_fa21_12_xor1;
  wire [0:0] u_csamul_cska32_fa21_12_or0;
  wire [0:0] u_csamul_cska32_and22_12;
  wire [0:0] u_csamul_cska32_fa22_12_xor1;
  wire [0:0] u_csamul_cska32_fa22_12_or0;
  wire [0:0] u_csamul_cska32_and23_12;
  wire [0:0] u_csamul_cska32_fa23_12_xor1;
  wire [0:0] u_csamul_cska32_fa23_12_or0;
  wire [0:0] u_csamul_cska32_and24_12;
  wire [0:0] u_csamul_cska32_fa24_12_xor1;
  wire [0:0] u_csamul_cska32_fa24_12_or0;
  wire [0:0] u_csamul_cska32_and25_12;
  wire [0:0] u_csamul_cska32_fa25_12_xor1;
  wire [0:0] u_csamul_cska32_fa25_12_or0;
  wire [0:0] u_csamul_cska32_and26_12;
  wire [0:0] u_csamul_cska32_fa26_12_xor1;
  wire [0:0] u_csamul_cska32_fa26_12_or0;
  wire [0:0] u_csamul_cska32_and27_12;
  wire [0:0] u_csamul_cska32_fa27_12_xor1;
  wire [0:0] u_csamul_cska32_fa27_12_or0;
  wire [0:0] u_csamul_cska32_and28_12;
  wire [0:0] u_csamul_cska32_fa28_12_xor1;
  wire [0:0] u_csamul_cska32_fa28_12_or0;
  wire [0:0] u_csamul_cska32_and29_12;
  wire [0:0] u_csamul_cska32_fa29_12_xor1;
  wire [0:0] u_csamul_cska32_fa29_12_or0;
  wire [0:0] u_csamul_cska32_and30_12;
  wire [0:0] u_csamul_cska32_fa30_12_xor1;
  wire [0:0] u_csamul_cska32_fa30_12_or0;
  wire [0:0] u_csamul_cska32_and31_12;
  wire [0:0] u_csamul_cska32_and0_13;
  wire [0:0] u_csamul_cska32_fa0_13_xor1;
  wire [0:0] u_csamul_cska32_fa0_13_or0;
  wire [0:0] u_csamul_cska32_and1_13;
  wire [0:0] u_csamul_cska32_fa1_13_xor1;
  wire [0:0] u_csamul_cska32_fa1_13_or0;
  wire [0:0] u_csamul_cska32_and2_13;
  wire [0:0] u_csamul_cska32_fa2_13_xor1;
  wire [0:0] u_csamul_cska32_fa2_13_or0;
  wire [0:0] u_csamul_cska32_and3_13;
  wire [0:0] u_csamul_cska32_fa3_13_xor1;
  wire [0:0] u_csamul_cska32_fa3_13_or0;
  wire [0:0] u_csamul_cska32_and4_13;
  wire [0:0] u_csamul_cska32_fa4_13_xor1;
  wire [0:0] u_csamul_cska32_fa4_13_or0;
  wire [0:0] u_csamul_cska32_and5_13;
  wire [0:0] u_csamul_cska32_fa5_13_xor1;
  wire [0:0] u_csamul_cska32_fa5_13_or0;
  wire [0:0] u_csamul_cska32_and6_13;
  wire [0:0] u_csamul_cska32_fa6_13_xor1;
  wire [0:0] u_csamul_cska32_fa6_13_or0;
  wire [0:0] u_csamul_cska32_and7_13;
  wire [0:0] u_csamul_cska32_fa7_13_xor1;
  wire [0:0] u_csamul_cska32_fa7_13_or0;
  wire [0:0] u_csamul_cska32_and8_13;
  wire [0:0] u_csamul_cska32_fa8_13_xor1;
  wire [0:0] u_csamul_cska32_fa8_13_or0;
  wire [0:0] u_csamul_cska32_and9_13;
  wire [0:0] u_csamul_cska32_fa9_13_xor1;
  wire [0:0] u_csamul_cska32_fa9_13_or0;
  wire [0:0] u_csamul_cska32_and10_13;
  wire [0:0] u_csamul_cska32_fa10_13_xor1;
  wire [0:0] u_csamul_cska32_fa10_13_or0;
  wire [0:0] u_csamul_cska32_and11_13;
  wire [0:0] u_csamul_cska32_fa11_13_xor1;
  wire [0:0] u_csamul_cska32_fa11_13_or0;
  wire [0:0] u_csamul_cska32_and12_13;
  wire [0:0] u_csamul_cska32_fa12_13_xor1;
  wire [0:0] u_csamul_cska32_fa12_13_or0;
  wire [0:0] u_csamul_cska32_and13_13;
  wire [0:0] u_csamul_cska32_fa13_13_xor1;
  wire [0:0] u_csamul_cska32_fa13_13_or0;
  wire [0:0] u_csamul_cska32_and14_13;
  wire [0:0] u_csamul_cska32_fa14_13_xor1;
  wire [0:0] u_csamul_cska32_fa14_13_or0;
  wire [0:0] u_csamul_cska32_and15_13;
  wire [0:0] u_csamul_cska32_fa15_13_xor1;
  wire [0:0] u_csamul_cska32_fa15_13_or0;
  wire [0:0] u_csamul_cska32_and16_13;
  wire [0:0] u_csamul_cska32_fa16_13_xor1;
  wire [0:0] u_csamul_cska32_fa16_13_or0;
  wire [0:0] u_csamul_cska32_and17_13;
  wire [0:0] u_csamul_cska32_fa17_13_xor1;
  wire [0:0] u_csamul_cska32_fa17_13_or0;
  wire [0:0] u_csamul_cska32_and18_13;
  wire [0:0] u_csamul_cska32_fa18_13_xor1;
  wire [0:0] u_csamul_cska32_fa18_13_or0;
  wire [0:0] u_csamul_cska32_and19_13;
  wire [0:0] u_csamul_cska32_fa19_13_xor1;
  wire [0:0] u_csamul_cska32_fa19_13_or0;
  wire [0:0] u_csamul_cska32_and20_13;
  wire [0:0] u_csamul_cska32_fa20_13_xor1;
  wire [0:0] u_csamul_cska32_fa20_13_or0;
  wire [0:0] u_csamul_cska32_and21_13;
  wire [0:0] u_csamul_cska32_fa21_13_xor1;
  wire [0:0] u_csamul_cska32_fa21_13_or0;
  wire [0:0] u_csamul_cska32_and22_13;
  wire [0:0] u_csamul_cska32_fa22_13_xor1;
  wire [0:0] u_csamul_cska32_fa22_13_or0;
  wire [0:0] u_csamul_cska32_and23_13;
  wire [0:0] u_csamul_cska32_fa23_13_xor1;
  wire [0:0] u_csamul_cska32_fa23_13_or0;
  wire [0:0] u_csamul_cska32_and24_13;
  wire [0:0] u_csamul_cska32_fa24_13_xor1;
  wire [0:0] u_csamul_cska32_fa24_13_or0;
  wire [0:0] u_csamul_cska32_and25_13;
  wire [0:0] u_csamul_cska32_fa25_13_xor1;
  wire [0:0] u_csamul_cska32_fa25_13_or0;
  wire [0:0] u_csamul_cska32_and26_13;
  wire [0:0] u_csamul_cska32_fa26_13_xor1;
  wire [0:0] u_csamul_cska32_fa26_13_or0;
  wire [0:0] u_csamul_cska32_and27_13;
  wire [0:0] u_csamul_cska32_fa27_13_xor1;
  wire [0:0] u_csamul_cska32_fa27_13_or0;
  wire [0:0] u_csamul_cska32_and28_13;
  wire [0:0] u_csamul_cska32_fa28_13_xor1;
  wire [0:0] u_csamul_cska32_fa28_13_or0;
  wire [0:0] u_csamul_cska32_and29_13;
  wire [0:0] u_csamul_cska32_fa29_13_xor1;
  wire [0:0] u_csamul_cska32_fa29_13_or0;
  wire [0:0] u_csamul_cska32_and30_13;
  wire [0:0] u_csamul_cska32_fa30_13_xor1;
  wire [0:0] u_csamul_cska32_fa30_13_or0;
  wire [0:0] u_csamul_cska32_and31_13;
  wire [0:0] u_csamul_cska32_and0_14;
  wire [0:0] u_csamul_cska32_fa0_14_xor1;
  wire [0:0] u_csamul_cska32_fa0_14_or0;
  wire [0:0] u_csamul_cska32_and1_14;
  wire [0:0] u_csamul_cska32_fa1_14_xor1;
  wire [0:0] u_csamul_cska32_fa1_14_or0;
  wire [0:0] u_csamul_cska32_and2_14;
  wire [0:0] u_csamul_cska32_fa2_14_xor1;
  wire [0:0] u_csamul_cska32_fa2_14_or0;
  wire [0:0] u_csamul_cska32_and3_14;
  wire [0:0] u_csamul_cska32_fa3_14_xor1;
  wire [0:0] u_csamul_cska32_fa3_14_or0;
  wire [0:0] u_csamul_cska32_and4_14;
  wire [0:0] u_csamul_cska32_fa4_14_xor1;
  wire [0:0] u_csamul_cska32_fa4_14_or0;
  wire [0:0] u_csamul_cska32_and5_14;
  wire [0:0] u_csamul_cska32_fa5_14_xor1;
  wire [0:0] u_csamul_cska32_fa5_14_or0;
  wire [0:0] u_csamul_cska32_and6_14;
  wire [0:0] u_csamul_cska32_fa6_14_xor1;
  wire [0:0] u_csamul_cska32_fa6_14_or0;
  wire [0:0] u_csamul_cska32_and7_14;
  wire [0:0] u_csamul_cska32_fa7_14_xor1;
  wire [0:0] u_csamul_cska32_fa7_14_or0;
  wire [0:0] u_csamul_cska32_and8_14;
  wire [0:0] u_csamul_cska32_fa8_14_xor1;
  wire [0:0] u_csamul_cska32_fa8_14_or0;
  wire [0:0] u_csamul_cska32_and9_14;
  wire [0:0] u_csamul_cska32_fa9_14_xor1;
  wire [0:0] u_csamul_cska32_fa9_14_or0;
  wire [0:0] u_csamul_cska32_and10_14;
  wire [0:0] u_csamul_cska32_fa10_14_xor1;
  wire [0:0] u_csamul_cska32_fa10_14_or0;
  wire [0:0] u_csamul_cska32_and11_14;
  wire [0:0] u_csamul_cska32_fa11_14_xor1;
  wire [0:0] u_csamul_cska32_fa11_14_or0;
  wire [0:0] u_csamul_cska32_and12_14;
  wire [0:0] u_csamul_cska32_fa12_14_xor1;
  wire [0:0] u_csamul_cska32_fa12_14_or0;
  wire [0:0] u_csamul_cska32_and13_14;
  wire [0:0] u_csamul_cska32_fa13_14_xor1;
  wire [0:0] u_csamul_cska32_fa13_14_or0;
  wire [0:0] u_csamul_cska32_and14_14;
  wire [0:0] u_csamul_cska32_fa14_14_xor1;
  wire [0:0] u_csamul_cska32_fa14_14_or0;
  wire [0:0] u_csamul_cska32_and15_14;
  wire [0:0] u_csamul_cska32_fa15_14_xor1;
  wire [0:0] u_csamul_cska32_fa15_14_or0;
  wire [0:0] u_csamul_cska32_and16_14;
  wire [0:0] u_csamul_cska32_fa16_14_xor1;
  wire [0:0] u_csamul_cska32_fa16_14_or0;
  wire [0:0] u_csamul_cska32_and17_14;
  wire [0:0] u_csamul_cska32_fa17_14_xor1;
  wire [0:0] u_csamul_cska32_fa17_14_or0;
  wire [0:0] u_csamul_cska32_and18_14;
  wire [0:0] u_csamul_cska32_fa18_14_xor1;
  wire [0:0] u_csamul_cska32_fa18_14_or0;
  wire [0:0] u_csamul_cska32_and19_14;
  wire [0:0] u_csamul_cska32_fa19_14_xor1;
  wire [0:0] u_csamul_cska32_fa19_14_or0;
  wire [0:0] u_csamul_cska32_and20_14;
  wire [0:0] u_csamul_cska32_fa20_14_xor1;
  wire [0:0] u_csamul_cska32_fa20_14_or0;
  wire [0:0] u_csamul_cska32_and21_14;
  wire [0:0] u_csamul_cska32_fa21_14_xor1;
  wire [0:0] u_csamul_cska32_fa21_14_or0;
  wire [0:0] u_csamul_cska32_and22_14;
  wire [0:0] u_csamul_cska32_fa22_14_xor1;
  wire [0:0] u_csamul_cska32_fa22_14_or0;
  wire [0:0] u_csamul_cska32_and23_14;
  wire [0:0] u_csamul_cska32_fa23_14_xor1;
  wire [0:0] u_csamul_cska32_fa23_14_or0;
  wire [0:0] u_csamul_cska32_and24_14;
  wire [0:0] u_csamul_cska32_fa24_14_xor1;
  wire [0:0] u_csamul_cska32_fa24_14_or0;
  wire [0:0] u_csamul_cska32_and25_14;
  wire [0:0] u_csamul_cska32_fa25_14_xor1;
  wire [0:0] u_csamul_cska32_fa25_14_or0;
  wire [0:0] u_csamul_cska32_and26_14;
  wire [0:0] u_csamul_cska32_fa26_14_xor1;
  wire [0:0] u_csamul_cska32_fa26_14_or0;
  wire [0:0] u_csamul_cska32_and27_14;
  wire [0:0] u_csamul_cska32_fa27_14_xor1;
  wire [0:0] u_csamul_cska32_fa27_14_or0;
  wire [0:0] u_csamul_cska32_and28_14;
  wire [0:0] u_csamul_cska32_fa28_14_xor1;
  wire [0:0] u_csamul_cska32_fa28_14_or0;
  wire [0:0] u_csamul_cska32_and29_14;
  wire [0:0] u_csamul_cska32_fa29_14_xor1;
  wire [0:0] u_csamul_cska32_fa29_14_or0;
  wire [0:0] u_csamul_cska32_and30_14;
  wire [0:0] u_csamul_cska32_fa30_14_xor1;
  wire [0:0] u_csamul_cska32_fa30_14_or0;
  wire [0:0] u_csamul_cska32_and31_14;
  wire [0:0] u_csamul_cska32_and0_15;
  wire [0:0] u_csamul_cska32_fa0_15_xor1;
  wire [0:0] u_csamul_cska32_fa0_15_or0;
  wire [0:0] u_csamul_cska32_and1_15;
  wire [0:0] u_csamul_cska32_fa1_15_xor1;
  wire [0:0] u_csamul_cska32_fa1_15_or0;
  wire [0:0] u_csamul_cska32_and2_15;
  wire [0:0] u_csamul_cska32_fa2_15_xor1;
  wire [0:0] u_csamul_cska32_fa2_15_or0;
  wire [0:0] u_csamul_cska32_and3_15;
  wire [0:0] u_csamul_cska32_fa3_15_xor1;
  wire [0:0] u_csamul_cska32_fa3_15_or0;
  wire [0:0] u_csamul_cska32_and4_15;
  wire [0:0] u_csamul_cska32_fa4_15_xor1;
  wire [0:0] u_csamul_cska32_fa4_15_or0;
  wire [0:0] u_csamul_cska32_and5_15;
  wire [0:0] u_csamul_cska32_fa5_15_xor1;
  wire [0:0] u_csamul_cska32_fa5_15_or0;
  wire [0:0] u_csamul_cska32_and6_15;
  wire [0:0] u_csamul_cska32_fa6_15_xor1;
  wire [0:0] u_csamul_cska32_fa6_15_or0;
  wire [0:0] u_csamul_cska32_and7_15;
  wire [0:0] u_csamul_cska32_fa7_15_xor1;
  wire [0:0] u_csamul_cska32_fa7_15_or0;
  wire [0:0] u_csamul_cska32_and8_15;
  wire [0:0] u_csamul_cska32_fa8_15_xor1;
  wire [0:0] u_csamul_cska32_fa8_15_or0;
  wire [0:0] u_csamul_cska32_and9_15;
  wire [0:0] u_csamul_cska32_fa9_15_xor1;
  wire [0:0] u_csamul_cska32_fa9_15_or0;
  wire [0:0] u_csamul_cska32_and10_15;
  wire [0:0] u_csamul_cska32_fa10_15_xor1;
  wire [0:0] u_csamul_cska32_fa10_15_or0;
  wire [0:0] u_csamul_cska32_and11_15;
  wire [0:0] u_csamul_cska32_fa11_15_xor1;
  wire [0:0] u_csamul_cska32_fa11_15_or0;
  wire [0:0] u_csamul_cska32_and12_15;
  wire [0:0] u_csamul_cska32_fa12_15_xor1;
  wire [0:0] u_csamul_cska32_fa12_15_or0;
  wire [0:0] u_csamul_cska32_and13_15;
  wire [0:0] u_csamul_cska32_fa13_15_xor1;
  wire [0:0] u_csamul_cska32_fa13_15_or0;
  wire [0:0] u_csamul_cska32_and14_15;
  wire [0:0] u_csamul_cska32_fa14_15_xor1;
  wire [0:0] u_csamul_cska32_fa14_15_or0;
  wire [0:0] u_csamul_cska32_and15_15;
  wire [0:0] u_csamul_cska32_fa15_15_xor1;
  wire [0:0] u_csamul_cska32_fa15_15_or0;
  wire [0:0] u_csamul_cska32_and16_15;
  wire [0:0] u_csamul_cska32_fa16_15_xor1;
  wire [0:0] u_csamul_cska32_fa16_15_or0;
  wire [0:0] u_csamul_cska32_and17_15;
  wire [0:0] u_csamul_cska32_fa17_15_xor1;
  wire [0:0] u_csamul_cska32_fa17_15_or0;
  wire [0:0] u_csamul_cska32_and18_15;
  wire [0:0] u_csamul_cska32_fa18_15_xor1;
  wire [0:0] u_csamul_cska32_fa18_15_or0;
  wire [0:0] u_csamul_cska32_and19_15;
  wire [0:0] u_csamul_cska32_fa19_15_xor1;
  wire [0:0] u_csamul_cska32_fa19_15_or0;
  wire [0:0] u_csamul_cska32_and20_15;
  wire [0:0] u_csamul_cska32_fa20_15_xor1;
  wire [0:0] u_csamul_cska32_fa20_15_or0;
  wire [0:0] u_csamul_cska32_and21_15;
  wire [0:0] u_csamul_cska32_fa21_15_xor1;
  wire [0:0] u_csamul_cska32_fa21_15_or0;
  wire [0:0] u_csamul_cska32_and22_15;
  wire [0:0] u_csamul_cska32_fa22_15_xor1;
  wire [0:0] u_csamul_cska32_fa22_15_or0;
  wire [0:0] u_csamul_cska32_and23_15;
  wire [0:0] u_csamul_cska32_fa23_15_xor1;
  wire [0:0] u_csamul_cska32_fa23_15_or0;
  wire [0:0] u_csamul_cska32_and24_15;
  wire [0:0] u_csamul_cska32_fa24_15_xor1;
  wire [0:0] u_csamul_cska32_fa24_15_or0;
  wire [0:0] u_csamul_cska32_and25_15;
  wire [0:0] u_csamul_cska32_fa25_15_xor1;
  wire [0:0] u_csamul_cska32_fa25_15_or0;
  wire [0:0] u_csamul_cska32_and26_15;
  wire [0:0] u_csamul_cska32_fa26_15_xor1;
  wire [0:0] u_csamul_cska32_fa26_15_or0;
  wire [0:0] u_csamul_cska32_and27_15;
  wire [0:0] u_csamul_cska32_fa27_15_xor1;
  wire [0:0] u_csamul_cska32_fa27_15_or0;
  wire [0:0] u_csamul_cska32_and28_15;
  wire [0:0] u_csamul_cska32_fa28_15_xor1;
  wire [0:0] u_csamul_cska32_fa28_15_or0;
  wire [0:0] u_csamul_cska32_and29_15;
  wire [0:0] u_csamul_cska32_fa29_15_xor1;
  wire [0:0] u_csamul_cska32_fa29_15_or0;
  wire [0:0] u_csamul_cska32_and30_15;
  wire [0:0] u_csamul_cska32_fa30_15_xor1;
  wire [0:0] u_csamul_cska32_fa30_15_or0;
  wire [0:0] u_csamul_cska32_and31_15;
  wire [0:0] u_csamul_cska32_and0_16;
  wire [0:0] u_csamul_cska32_fa0_16_xor1;
  wire [0:0] u_csamul_cska32_fa0_16_or0;
  wire [0:0] u_csamul_cska32_and1_16;
  wire [0:0] u_csamul_cska32_fa1_16_xor1;
  wire [0:0] u_csamul_cska32_fa1_16_or0;
  wire [0:0] u_csamul_cska32_and2_16;
  wire [0:0] u_csamul_cska32_fa2_16_xor1;
  wire [0:0] u_csamul_cska32_fa2_16_or0;
  wire [0:0] u_csamul_cska32_and3_16;
  wire [0:0] u_csamul_cska32_fa3_16_xor1;
  wire [0:0] u_csamul_cska32_fa3_16_or0;
  wire [0:0] u_csamul_cska32_and4_16;
  wire [0:0] u_csamul_cska32_fa4_16_xor1;
  wire [0:0] u_csamul_cska32_fa4_16_or0;
  wire [0:0] u_csamul_cska32_and5_16;
  wire [0:0] u_csamul_cska32_fa5_16_xor1;
  wire [0:0] u_csamul_cska32_fa5_16_or0;
  wire [0:0] u_csamul_cska32_and6_16;
  wire [0:0] u_csamul_cska32_fa6_16_xor1;
  wire [0:0] u_csamul_cska32_fa6_16_or0;
  wire [0:0] u_csamul_cska32_and7_16;
  wire [0:0] u_csamul_cska32_fa7_16_xor1;
  wire [0:0] u_csamul_cska32_fa7_16_or0;
  wire [0:0] u_csamul_cska32_and8_16;
  wire [0:0] u_csamul_cska32_fa8_16_xor1;
  wire [0:0] u_csamul_cska32_fa8_16_or0;
  wire [0:0] u_csamul_cska32_and9_16;
  wire [0:0] u_csamul_cska32_fa9_16_xor1;
  wire [0:0] u_csamul_cska32_fa9_16_or0;
  wire [0:0] u_csamul_cska32_and10_16;
  wire [0:0] u_csamul_cska32_fa10_16_xor1;
  wire [0:0] u_csamul_cska32_fa10_16_or0;
  wire [0:0] u_csamul_cska32_and11_16;
  wire [0:0] u_csamul_cska32_fa11_16_xor1;
  wire [0:0] u_csamul_cska32_fa11_16_or0;
  wire [0:0] u_csamul_cska32_and12_16;
  wire [0:0] u_csamul_cska32_fa12_16_xor1;
  wire [0:0] u_csamul_cska32_fa12_16_or0;
  wire [0:0] u_csamul_cska32_and13_16;
  wire [0:0] u_csamul_cska32_fa13_16_xor1;
  wire [0:0] u_csamul_cska32_fa13_16_or0;
  wire [0:0] u_csamul_cska32_and14_16;
  wire [0:0] u_csamul_cska32_fa14_16_xor1;
  wire [0:0] u_csamul_cska32_fa14_16_or0;
  wire [0:0] u_csamul_cska32_and15_16;
  wire [0:0] u_csamul_cska32_fa15_16_xor1;
  wire [0:0] u_csamul_cska32_fa15_16_or0;
  wire [0:0] u_csamul_cska32_and16_16;
  wire [0:0] u_csamul_cska32_fa16_16_xor1;
  wire [0:0] u_csamul_cska32_fa16_16_or0;
  wire [0:0] u_csamul_cska32_and17_16;
  wire [0:0] u_csamul_cska32_fa17_16_xor1;
  wire [0:0] u_csamul_cska32_fa17_16_or0;
  wire [0:0] u_csamul_cska32_and18_16;
  wire [0:0] u_csamul_cska32_fa18_16_xor1;
  wire [0:0] u_csamul_cska32_fa18_16_or0;
  wire [0:0] u_csamul_cska32_and19_16;
  wire [0:0] u_csamul_cska32_fa19_16_xor1;
  wire [0:0] u_csamul_cska32_fa19_16_or0;
  wire [0:0] u_csamul_cska32_and20_16;
  wire [0:0] u_csamul_cska32_fa20_16_xor1;
  wire [0:0] u_csamul_cska32_fa20_16_or0;
  wire [0:0] u_csamul_cska32_and21_16;
  wire [0:0] u_csamul_cska32_fa21_16_xor1;
  wire [0:0] u_csamul_cska32_fa21_16_or0;
  wire [0:0] u_csamul_cska32_and22_16;
  wire [0:0] u_csamul_cska32_fa22_16_xor1;
  wire [0:0] u_csamul_cska32_fa22_16_or0;
  wire [0:0] u_csamul_cska32_and23_16;
  wire [0:0] u_csamul_cska32_fa23_16_xor1;
  wire [0:0] u_csamul_cska32_fa23_16_or0;
  wire [0:0] u_csamul_cska32_and24_16;
  wire [0:0] u_csamul_cska32_fa24_16_xor1;
  wire [0:0] u_csamul_cska32_fa24_16_or0;
  wire [0:0] u_csamul_cska32_and25_16;
  wire [0:0] u_csamul_cska32_fa25_16_xor1;
  wire [0:0] u_csamul_cska32_fa25_16_or0;
  wire [0:0] u_csamul_cska32_and26_16;
  wire [0:0] u_csamul_cska32_fa26_16_xor1;
  wire [0:0] u_csamul_cska32_fa26_16_or0;
  wire [0:0] u_csamul_cska32_and27_16;
  wire [0:0] u_csamul_cska32_fa27_16_xor1;
  wire [0:0] u_csamul_cska32_fa27_16_or0;
  wire [0:0] u_csamul_cska32_and28_16;
  wire [0:0] u_csamul_cska32_fa28_16_xor1;
  wire [0:0] u_csamul_cska32_fa28_16_or0;
  wire [0:0] u_csamul_cska32_and29_16;
  wire [0:0] u_csamul_cska32_fa29_16_xor1;
  wire [0:0] u_csamul_cska32_fa29_16_or0;
  wire [0:0] u_csamul_cska32_and30_16;
  wire [0:0] u_csamul_cska32_fa30_16_xor1;
  wire [0:0] u_csamul_cska32_fa30_16_or0;
  wire [0:0] u_csamul_cska32_and31_16;
  wire [0:0] u_csamul_cska32_and0_17;
  wire [0:0] u_csamul_cska32_fa0_17_xor1;
  wire [0:0] u_csamul_cska32_fa0_17_or0;
  wire [0:0] u_csamul_cska32_and1_17;
  wire [0:0] u_csamul_cska32_fa1_17_xor1;
  wire [0:0] u_csamul_cska32_fa1_17_or0;
  wire [0:0] u_csamul_cska32_and2_17;
  wire [0:0] u_csamul_cska32_fa2_17_xor1;
  wire [0:0] u_csamul_cska32_fa2_17_or0;
  wire [0:0] u_csamul_cska32_and3_17;
  wire [0:0] u_csamul_cska32_fa3_17_xor1;
  wire [0:0] u_csamul_cska32_fa3_17_or0;
  wire [0:0] u_csamul_cska32_and4_17;
  wire [0:0] u_csamul_cska32_fa4_17_xor1;
  wire [0:0] u_csamul_cska32_fa4_17_or0;
  wire [0:0] u_csamul_cska32_and5_17;
  wire [0:0] u_csamul_cska32_fa5_17_xor1;
  wire [0:0] u_csamul_cska32_fa5_17_or0;
  wire [0:0] u_csamul_cska32_and6_17;
  wire [0:0] u_csamul_cska32_fa6_17_xor1;
  wire [0:0] u_csamul_cska32_fa6_17_or0;
  wire [0:0] u_csamul_cska32_and7_17;
  wire [0:0] u_csamul_cska32_fa7_17_xor1;
  wire [0:0] u_csamul_cska32_fa7_17_or0;
  wire [0:0] u_csamul_cska32_and8_17;
  wire [0:0] u_csamul_cska32_fa8_17_xor1;
  wire [0:0] u_csamul_cska32_fa8_17_or0;
  wire [0:0] u_csamul_cska32_and9_17;
  wire [0:0] u_csamul_cska32_fa9_17_xor1;
  wire [0:0] u_csamul_cska32_fa9_17_or0;
  wire [0:0] u_csamul_cska32_and10_17;
  wire [0:0] u_csamul_cska32_fa10_17_xor1;
  wire [0:0] u_csamul_cska32_fa10_17_or0;
  wire [0:0] u_csamul_cska32_and11_17;
  wire [0:0] u_csamul_cska32_fa11_17_xor1;
  wire [0:0] u_csamul_cska32_fa11_17_or0;
  wire [0:0] u_csamul_cska32_and12_17;
  wire [0:0] u_csamul_cska32_fa12_17_xor1;
  wire [0:0] u_csamul_cska32_fa12_17_or0;
  wire [0:0] u_csamul_cska32_and13_17;
  wire [0:0] u_csamul_cska32_fa13_17_xor1;
  wire [0:0] u_csamul_cska32_fa13_17_or0;
  wire [0:0] u_csamul_cska32_and14_17;
  wire [0:0] u_csamul_cska32_fa14_17_xor1;
  wire [0:0] u_csamul_cska32_fa14_17_or0;
  wire [0:0] u_csamul_cska32_and15_17;
  wire [0:0] u_csamul_cska32_fa15_17_xor1;
  wire [0:0] u_csamul_cska32_fa15_17_or0;
  wire [0:0] u_csamul_cska32_and16_17;
  wire [0:0] u_csamul_cska32_fa16_17_xor1;
  wire [0:0] u_csamul_cska32_fa16_17_or0;
  wire [0:0] u_csamul_cska32_and17_17;
  wire [0:0] u_csamul_cska32_fa17_17_xor1;
  wire [0:0] u_csamul_cska32_fa17_17_or0;
  wire [0:0] u_csamul_cska32_and18_17;
  wire [0:0] u_csamul_cska32_fa18_17_xor1;
  wire [0:0] u_csamul_cska32_fa18_17_or0;
  wire [0:0] u_csamul_cska32_and19_17;
  wire [0:0] u_csamul_cska32_fa19_17_xor1;
  wire [0:0] u_csamul_cska32_fa19_17_or0;
  wire [0:0] u_csamul_cska32_and20_17;
  wire [0:0] u_csamul_cska32_fa20_17_xor1;
  wire [0:0] u_csamul_cska32_fa20_17_or0;
  wire [0:0] u_csamul_cska32_and21_17;
  wire [0:0] u_csamul_cska32_fa21_17_xor1;
  wire [0:0] u_csamul_cska32_fa21_17_or0;
  wire [0:0] u_csamul_cska32_and22_17;
  wire [0:0] u_csamul_cska32_fa22_17_xor1;
  wire [0:0] u_csamul_cska32_fa22_17_or0;
  wire [0:0] u_csamul_cska32_and23_17;
  wire [0:0] u_csamul_cska32_fa23_17_xor1;
  wire [0:0] u_csamul_cska32_fa23_17_or0;
  wire [0:0] u_csamul_cska32_and24_17;
  wire [0:0] u_csamul_cska32_fa24_17_xor1;
  wire [0:0] u_csamul_cska32_fa24_17_or0;
  wire [0:0] u_csamul_cska32_and25_17;
  wire [0:0] u_csamul_cska32_fa25_17_xor1;
  wire [0:0] u_csamul_cska32_fa25_17_or0;
  wire [0:0] u_csamul_cska32_and26_17;
  wire [0:0] u_csamul_cska32_fa26_17_xor1;
  wire [0:0] u_csamul_cska32_fa26_17_or0;
  wire [0:0] u_csamul_cska32_and27_17;
  wire [0:0] u_csamul_cska32_fa27_17_xor1;
  wire [0:0] u_csamul_cska32_fa27_17_or0;
  wire [0:0] u_csamul_cska32_and28_17;
  wire [0:0] u_csamul_cska32_fa28_17_xor1;
  wire [0:0] u_csamul_cska32_fa28_17_or0;
  wire [0:0] u_csamul_cska32_and29_17;
  wire [0:0] u_csamul_cska32_fa29_17_xor1;
  wire [0:0] u_csamul_cska32_fa29_17_or0;
  wire [0:0] u_csamul_cska32_and30_17;
  wire [0:0] u_csamul_cska32_fa30_17_xor1;
  wire [0:0] u_csamul_cska32_fa30_17_or0;
  wire [0:0] u_csamul_cska32_and31_17;
  wire [0:0] u_csamul_cska32_and0_18;
  wire [0:0] u_csamul_cska32_fa0_18_xor1;
  wire [0:0] u_csamul_cska32_fa0_18_or0;
  wire [0:0] u_csamul_cska32_and1_18;
  wire [0:0] u_csamul_cska32_fa1_18_xor1;
  wire [0:0] u_csamul_cska32_fa1_18_or0;
  wire [0:0] u_csamul_cska32_and2_18;
  wire [0:0] u_csamul_cska32_fa2_18_xor1;
  wire [0:0] u_csamul_cska32_fa2_18_or0;
  wire [0:0] u_csamul_cska32_and3_18;
  wire [0:0] u_csamul_cska32_fa3_18_xor1;
  wire [0:0] u_csamul_cska32_fa3_18_or0;
  wire [0:0] u_csamul_cska32_and4_18;
  wire [0:0] u_csamul_cska32_fa4_18_xor1;
  wire [0:0] u_csamul_cska32_fa4_18_or0;
  wire [0:0] u_csamul_cska32_and5_18;
  wire [0:0] u_csamul_cska32_fa5_18_xor1;
  wire [0:0] u_csamul_cska32_fa5_18_or0;
  wire [0:0] u_csamul_cska32_and6_18;
  wire [0:0] u_csamul_cska32_fa6_18_xor1;
  wire [0:0] u_csamul_cska32_fa6_18_or0;
  wire [0:0] u_csamul_cska32_and7_18;
  wire [0:0] u_csamul_cska32_fa7_18_xor1;
  wire [0:0] u_csamul_cska32_fa7_18_or0;
  wire [0:0] u_csamul_cska32_and8_18;
  wire [0:0] u_csamul_cska32_fa8_18_xor1;
  wire [0:0] u_csamul_cska32_fa8_18_or0;
  wire [0:0] u_csamul_cska32_and9_18;
  wire [0:0] u_csamul_cska32_fa9_18_xor1;
  wire [0:0] u_csamul_cska32_fa9_18_or0;
  wire [0:0] u_csamul_cska32_and10_18;
  wire [0:0] u_csamul_cska32_fa10_18_xor1;
  wire [0:0] u_csamul_cska32_fa10_18_or0;
  wire [0:0] u_csamul_cska32_and11_18;
  wire [0:0] u_csamul_cska32_fa11_18_xor1;
  wire [0:0] u_csamul_cska32_fa11_18_or0;
  wire [0:0] u_csamul_cska32_and12_18;
  wire [0:0] u_csamul_cska32_fa12_18_xor1;
  wire [0:0] u_csamul_cska32_fa12_18_or0;
  wire [0:0] u_csamul_cska32_and13_18;
  wire [0:0] u_csamul_cska32_fa13_18_xor1;
  wire [0:0] u_csamul_cska32_fa13_18_or0;
  wire [0:0] u_csamul_cska32_and14_18;
  wire [0:0] u_csamul_cska32_fa14_18_xor1;
  wire [0:0] u_csamul_cska32_fa14_18_or0;
  wire [0:0] u_csamul_cska32_and15_18;
  wire [0:0] u_csamul_cska32_fa15_18_xor1;
  wire [0:0] u_csamul_cska32_fa15_18_or0;
  wire [0:0] u_csamul_cska32_and16_18;
  wire [0:0] u_csamul_cska32_fa16_18_xor1;
  wire [0:0] u_csamul_cska32_fa16_18_or0;
  wire [0:0] u_csamul_cska32_and17_18;
  wire [0:0] u_csamul_cska32_fa17_18_xor1;
  wire [0:0] u_csamul_cska32_fa17_18_or0;
  wire [0:0] u_csamul_cska32_and18_18;
  wire [0:0] u_csamul_cska32_fa18_18_xor1;
  wire [0:0] u_csamul_cska32_fa18_18_or0;
  wire [0:0] u_csamul_cska32_and19_18;
  wire [0:0] u_csamul_cska32_fa19_18_xor1;
  wire [0:0] u_csamul_cska32_fa19_18_or0;
  wire [0:0] u_csamul_cska32_and20_18;
  wire [0:0] u_csamul_cska32_fa20_18_xor1;
  wire [0:0] u_csamul_cska32_fa20_18_or0;
  wire [0:0] u_csamul_cska32_and21_18;
  wire [0:0] u_csamul_cska32_fa21_18_xor1;
  wire [0:0] u_csamul_cska32_fa21_18_or0;
  wire [0:0] u_csamul_cska32_and22_18;
  wire [0:0] u_csamul_cska32_fa22_18_xor1;
  wire [0:0] u_csamul_cska32_fa22_18_or0;
  wire [0:0] u_csamul_cska32_and23_18;
  wire [0:0] u_csamul_cska32_fa23_18_xor1;
  wire [0:0] u_csamul_cska32_fa23_18_or0;
  wire [0:0] u_csamul_cska32_and24_18;
  wire [0:0] u_csamul_cska32_fa24_18_xor1;
  wire [0:0] u_csamul_cska32_fa24_18_or0;
  wire [0:0] u_csamul_cska32_and25_18;
  wire [0:0] u_csamul_cska32_fa25_18_xor1;
  wire [0:0] u_csamul_cska32_fa25_18_or0;
  wire [0:0] u_csamul_cska32_and26_18;
  wire [0:0] u_csamul_cska32_fa26_18_xor1;
  wire [0:0] u_csamul_cska32_fa26_18_or0;
  wire [0:0] u_csamul_cska32_and27_18;
  wire [0:0] u_csamul_cska32_fa27_18_xor1;
  wire [0:0] u_csamul_cska32_fa27_18_or0;
  wire [0:0] u_csamul_cska32_and28_18;
  wire [0:0] u_csamul_cska32_fa28_18_xor1;
  wire [0:0] u_csamul_cska32_fa28_18_or0;
  wire [0:0] u_csamul_cska32_and29_18;
  wire [0:0] u_csamul_cska32_fa29_18_xor1;
  wire [0:0] u_csamul_cska32_fa29_18_or0;
  wire [0:0] u_csamul_cska32_and30_18;
  wire [0:0] u_csamul_cska32_fa30_18_xor1;
  wire [0:0] u_csamul_cska32_fa30_18_or0;
  wire [0:0] u_csamul_cska32_and31_18;
  wire [0:0] u_csamul_cska32_and0_19;
  wire [0:0] u_csamul_cska32_fa0_19_xor1;
  wire [0:0] u_csamul_cska32_fa0_19_or0;
  wire [0:0] u_csamul_cska32_and1_19;
  wire [0:0] u_csamul_cska32_fa1_19_xor1;
  wire [0:0] u_csamul_cska32_fa1_19_or0;
  wire [0:0] u_csamul_cska32_and2_19;
  wire [0:0] u_csamul_cska32_fa2_19_xor1;
  wire [0:0] u_csamul_cska32_fa2_19_or0;
  wire [0:0] u_csamul_cska32_and3_19;
  wire [0:0] u_csamul_cska32_fa3_19_xor1;
  wire [0:0] u_csamul_cska32_fa3_19_or0;
  wire [0:0] u_csamul_cska32_and4_19;
  wire [0:0] u_csamul_cska32_fa4_19_xor1;
  wire [0:0] u_csamul_cska32_fa4_19_or0;
  wire [0:0] u_csamul_cska32_and5_19;
  wire [0:0] u_csamul_cska32_fa5_19_xor1;
  wire [0:0] u_csamul_cska32_fa5_19_or0;
  wire [0:0] u_csamul_cska32_and6_19;
  wire [0:0] u_csamul_cska32_fa6_19_xor1;
  wire [0:0] u_csamul_cska32_fa6_19_or0;
  wire [0:0] u_csamul_cska32_and7_19;
  wire [0:0] u_csamul_cska32_fa7_19_xor1;
  wire [0:0] u_csamul_cska32_fa7_19_or0;
  wire [0:0] u_csamul_cska32_and8_19;
  wire [0:0] u_csamul_cska32_fa8_19_xor1;
  wire [0:0] u_csamul_cska32_fa8_19_or0;
  wire [0:0] u_csamul_cska32_and9_19;
  wire [0:0] u_csamul_cska32_fa9_19_xor1;
  wire [0:0] u_csamul_cska32_fa9_19_or0;
  wire [0:0] u_csamul_cska32_and10_19;
  wire [0:0] u_csamul_cska32_fa10_19_xor1;
  wire [0:0] u_csamul_cska32_fa10_19_or0;
  wire [0:0] u_csamul_cska32_and11_19;
  wire [0:0] u_csamul_cska32_fa11_19_xor1;
  wire [0:0] u_csamul_cska32_fa11_19_or0;
  wire [0:0] u_csamul_cska32_and12_19;
  wire [0:0] u_csamul_cska32_fa12_19_xor1;
  wire [0:0] u_csamul_cska32_fa12_19_or0;
  wire [0:0] u_csamul_cska32_and13_19;
  wire [0:0] u_csamul_cska32_fa13_19_xor1;
  wire [0:0] u_csamul_cska32_fa13_19_or0;
  wire [0:0] u_csamul_cska32_and14_19;
  wire [0:0] u_csamul_cska32_fa14_19_xor1;
  wire [0:0] u_csamul_cska32_fa14_19_or0;
  wire [0:0] u_csamul_cska32_and15_19;
  wire [0:0] u_csamul_cska32_fa15_19_xor1;
  wire [0:0] u_csamul_cska32_fa15_19_or0;
  wire [0:0] u_csamul_cska32_and16_19;
  wire [0:0] u_csamul_cska32_fa16_19_xor1;
  wire [0:0] u_csamul_cska32_fa16_19_or0;
  wire [0:0] u_csamul_cska32_and17_19;
  wire [0:0] u_csamul_cska32_fa17_19_xor1;
  wire [0:0] u_csamul_cska32_fa17_19_or0;
  wire [0:0] u_csamul_cska32_and18_19;
  wire [0:0] u_csamul_cska32_fa18_19_xor1;
  wire [0:0] u_csamul_cska32_fa18_19_or0;
  wire [0:0] u_csamul_cska32_and19_19;
  wire [0:0] u_csamul_cska32_fa19_19_xor1;
  wire [0:0] u_csamul_cska32_fa19_19_or0;
  wire [0:0] u_csamul_cska32_and20_19;
  wire [0:0] u_csamul_cska32_fa20_19_xor1;
  wire [0:0] u_csamul_cska32_fa20_19_or0;
  wire [0:0] u_csamul_cska32_and21_19;
  wire [0:0] u_csamul_cska32_fa21_19_xor1;
  wire [0:0] u_csamul_cska32_fa21_19_or0;
  wire [0:0] u_csamul_cska32_and22_19;
  wire [0:0] u_csamul_cska32_fa22_19_xor1;
  wire [0:0] u_csamul_cska32_fa22_19_or0;
  wire [0:0] u_csamul_cska32_and23_19;
  wire [0:0] u_csamul_cska32_fa23_19_xor1;
  wire [0:0] u_csamul_cska32_fa23_19_or0;
  wire [0:0] u_csamul_cska32_and24_19;
  wire [0:0] u_csamul_cska32_fa24_19_xor1;
  wire [0:0] u_csamul_cska32_fa24_19_or0;
  wire [0:0] u_csamul_cska32_and25_19;
  wire [0:0] u_csamul_cska32_fa25_19_xor1;
  wire [0:0] u_csamul_cska32_fa25_19_or0;
  wire [0:0] u_csamul_cska32_and26_19;
  wire [0:0] u_csamul_cska32_fa26_19_xor1;
  wire [0:0] u_csamul_cska32_fa26_19_or0;
  wire [0:0] u_csamul_cska32_and27_19;
  wire [0:0] u_csamul_cska32_fa27_19_xor1;
  wire [0:0] u_csamul_cska32_fa27_19_or0;
  wire [0:0] u_csamul_cska32_and28_19;
  wire [0:0] u_csamul_cska32_fa28_19_xor1;
  wire [0:0] u_csamul_cska32_fa28_19_or0;
  wire [0:0] u_csamul_cska32_and29_19;
  wire [0:0] u_csamul_cska32_fa29_19_xor1;
  wire [0:0] u_csamul_cska32_fa29_19_or0;
  wire [0:0] u_csamul_cska32_and30_19;
  wire [0:0] u_csamul_cska32_fa30_19_xor1;
  wire [0:0] u_csamul_cska32_fa30_19_or0;
  wire [0:0] u_csamul_cska32_and31_19;
  wire [0:0] u_csamul_cska32_and0_20;
  wire [0:0] u_csamul_cska32_fa0_20_xor1;
  wire [0:0] u_csamul_cska32_fa0_20_or0;
  wire [0:0] u_csamul_cska32_and1_20;
  wire [0:0] u_csamul_cska32_fa1_20_xor1;
  wire [0:0] u_csamul_cska32_fa1_20_or0;
  wire [0:0] u_csamul_cska32_and2_20;
  wire [0:0] u_csamul_cska32_fa2_20_xor1;
  wire [0:0] u_csamul_cska32_fa2_20_or0;
  wire [0:0] u_csamul_cska32_and3_20;
  wire [0:0] u_csamul_cska32_fa3_20_xor1;
  wire [0:0] u_csamul_cska32_fa3_20_or0;
  wire [0:0] u_csamul_cska32_and4_20;
  wire [0:0] u_csamul_cska32_fa4_20_xor1;
  wire [0:0] u_csamul_cska32_fa4_20_or0;
  wire [0:0] u_csamul_cska32_and5_20;
  wire [0:0] u_csamul_cska32_fa5_20_xor1;
  wire [0:0] u_csamul_cska32_fa5_20_or0;
  wire [0:0] u_csamul_cska32_and6_20;
  wire [0:0] u_csamul_cska32_fa6_20_xor1;
  wire [0:0] u_csamul_cska32_fa6_20_or0;
  wire [0:0] u_csamul_cska32_and7_20;
  wire [0:0] u_csamul_cska32_fa7_20_xor1;
  wire [0:0] u_csamul_cska32_fa7_20_or0;
  wire [0:0] u_csamul_cska32_and8_20;
  wire [0:0] u_csamul_cska32_fa8_20_xor1;
  wire [0:0] u_csamul_cska32_fa8_20_or0;
  wire [0:0] u_csamul_cska32_and9_20;
  wire [0:0] u_csamul_cska32_fa9_20_xor1;
  wire [0:0] u_csamul_cska32_fa9_20_or0;
  wire [0:0] u_csamul_cska32_and10_20;
  wire [0:0] u_csamul_cska32_fa10_20_xor1;
  wire [0:0] u_csamul_cska32_fa10_20_or0;
  wire [0:0] u_csamul_cska32_and11_20;
  wire [0:0] u_csamul_cska32_fa11_20_xor1;
  wire [0:0] u_csamul_cska32_fa11_20_or0;
  wire [0:0] u_csamul_cska32_and12_20;
  wire [0:0] u_csamul_cska32_fa12_20_xor1;
  wire [0:0] u_csamul_cska32_fa12_20_or0;
  wire [0:0] u_csamul_cska32_and13_20;
  wire [0:0] u_csamul_cska32_fa13_20_xor1;
  wire [0:0] u_csamul_cska32_fa13_20_or0;
  wire [0:0] u_csamul_cska32_and14_20;
  wire [0:0] u_csamul_cska32_fa14_20_xor1;
  wire [0:0] u_csamul_cska32_fa14_20_or0;
  wire [0:0] u_csamul_cska32_and15_20;
  wire [0:0] u_csamul_cska32_fa15_20_xor1;
  wire [0:0] u_csamul_cska32_fa15_20_or0;
  wire [0:0] u_csamul_cska32_and16_20;
  wire [0:0] u_csamul_cska32_fa16_20_xor1;
  wire [0:0] u_csamul_cska32_fa16_20_or0;
  wire [0:0] u_csamul_cska32_and17_20;
  wire [0:0] u_csamul_cska32_fa17_20_xor1;
  wire [0:0] u_csamul_cska32_fa17_20_or0;
  wire [0:0] u_csamul_cska32_and18_20;
  wire [0:0] u_csamul_cska32_fa18_20_xor1;
  wire [0:0] u_csamul_cska32_fa18_20_or0;
  wire [0:0] u_csamul_cska32_and19_20;
  wire [0:0] u_csamul_cska32_fa19_20_xor1;
  wire [0:0] u_csamul_cska32_fa19_20_or0;
  wire [0:0] u_csamul_cska32_and20_20;
  wire [0:0] u_csamul_cska32_fa20_20_xor1;
  wire [0:0] u_csamul_cska32_fa20_20_or0;
  wire [0:0] u_csamul_cska32_and21_20;
  wire [0:0] u_csamul_cska32_fa21_20_xor1;
  wire [0:0] u_csamul_cska32_fa21_20_or0;
  wire [0:0] u_csamul_cska32_and22_20;
  wire [0:0] u_csamul_cska32_fa22_20_xor1;
  wire [0:0] u_csamul_cska32_fa22_20_or0;
  wire [0:0] u_csamul_cska32_and23_20;
  wire [0:0] u_csamul_cska32_fa23_20_xor1;
  wire [0:0] u_csamul_cska32_fa23_20_or0;
  wire [0:0] u_csamul_cska32_and24_20;
  wire [0:0] u_csamul_cska32_fa24_20_xor1;
  wire [0:0] u_csamul_cska32_fa24_20_or0;
  wire [0:0] u_csamul_cska32_and25_20;
  wire [0:0] u_csamul_cska32_fa25_20_xor1;
  wire [0:0] u_csamul_cska32_fa25_20_or0;
  wire [0:0] u_csamul_cska32_and26_20;
  wire [0:0] u_csamul_cska32_fa26_20_xor1;
  wire [0:0] u_csamul_cska32_fa26_20_or0;
  wire [0:0] u_csamul_cska32_and27_20;
  wire [0:0] u_csamul_cska32_fa27_20_xor1;
  wire [0:0] u_csamul_cska32_fa27_20_or0;
  wire [0:0] u_csamul_cska32_and28_20;
  wire [0:0] u_csamul_cska32_fa28_20_xor1;
  wire [0:0] u_csamul_cska32_fa28_20_or0;
  wire [0:0] u_csamul_cska32_and29_20;
  wire [0:0] u_csamul_cska32_fa29_20_xor1;
  wire [0:0] u_csamul_cska32_fa29_20_or0;
  wire [0:0] u_csamul_cska32_and30_20;
  wire [0:0] u_csamul_cska32_fa30_20_xor1;
  wire [0:0] u_csamul_cska32_fa30_20_or0;
  wire [0:0] u_csamul_cska32_and31_20;
  wire [0:0] u_csamul_cska32_and0_21;
  wire [0:0] u_csamul_cska32_fa0_21_xor1;
  wire [0:0] u_csamul_cska32_fa0_21_or0;
  wire [0:0] u_csamul_cska32_and1_21;
  wire [0:0] u_csamul_cska32_fa1_21_xor1;
  wire [0:0] u_csamul_cska32_fa1_21_or0;
  wire [0:0] u_csamul_cska32_and2_21;
  wire [0:0] u_csamul_cska32_fa2_21_xor1;
  wire [0:0] u_csamul_cska32_fa2_21_or0;
  wire [0:0] u_csamul_cska32_and3_21;
  wire [0:0] u_csamul_cska32_fa3_21_xor1;
  wire [0:0] u_csamul_cska32_fa3_21_or0;
  wire [0:0] u_csamul_cska32_and4_21;
  wire [0:0] u_csamul_cska32_fa4_21_xor1;
  wire [0:0] u_csamul_cska32_fa4_21_or0;
  wire [0:0] u_csamul_cska32_and5_21;
  wire [0:0] u_csamul_cska32_fa5_21_xor1;
  wire [0:0] u_csamul_cska32_fa5_21_or0;
  wire [0:0] u_csamul_cska32_and6_21;
  wire [0:0] u_csamul_cska32_fa6_21_xor1;
  wire [0:0] u_csamul_cska32_fa6_21_or0;
  wire [0:0] u_csamul_cska32_and7_21;
  wire [0:0] u_csamul_cska32_fa7_21_xor1;
  wire [0:0] u_csamul_cska32_fa7_21_or0;
  wire [0:0] u_csamul_cska32_and8_21;
  wire [0:0] u_csamul_cska32_fa8_21_xor1;
  wire [0:0] u_csamul_cska32_fa8_21_or0;
  wire [0:0] u_csamul_cska32_and9_21;
  wire [0:0] u_csamul_cska32_fa9_21_xor1;
  wire [0:0] u_csamul_cska32_fa9_21_or0;
  wire [0:0] u_csamul_cska32_and10_21;
  wire [0:0] u_csamul_cska32_fa10_21_xor1;
  wire [0:0] u_csamul_cska32_fa10_21_or0;
  wire [0:0] u_csamul_cska32_and11_21;
  wire [0:0] u_csamul_cska32_fa11_21_xor1;
  wire [0:0] u_csamul_cska32_fa11_21_or0;
  wire [0:0] u_csamul_cska32_and12_21;
  wire [0:0] u_csamul_cska32_fa12_21_xor1;
  wire [0:0] u_csamul_cska32_fa12_21_or0;
  wire [0:0] u_csamul_cska32_and13_21;
  wire [0:0] u_csamul_cska32_fa13_21_xor1;
  wire [0:0] u_csamul_cska32_fa13_21_or0;
  wire [0:0] u_csamul_cska32_and14_21;
  wire [0:0] u_csamul_cska32_fa14_21_xor1;
  wire [0:0] u_csamul_cska32_fa14_21_or0;
  wire [0:0] u_csamul_cska32_and15_21;
  wire [0:0] u_csamul_cska32_fa15_21_xor1;
  wire [0:0] u_csamul_cska32_fa15_21_or0;
  wire [0:0] u_csamul_cska32_and16_21;
  wire [0:0] u_csamul_cska32_fa16_21_xor1;
  wire [0:0] u_csamul_cska32_fa16_21_or0;
  wire [0:0] u_csamul_cska32_and17_21;
  wire [0:0] u_csamul_cska32_fa17_21_xor1;
  wire [0:0] u_csamul_cska32_fa17_21_or0;
  wire [0:0] u_csamul_cska32_and18_21;
  wire [0:0] u_csamul_cska32_fa18_21_xor1;
  wire [0:0] u_csamul_cska32_fa18_21_or0;
  wire [0:0] u_csamul_cska32_and19_21;
  wire [0:0] u_csamul_cska32_fa19_21_xor1;
  wire [0:0] u_csamul_cska32_fa19_21_or0;
  wire [0:0] u_csamul_cska32_and20_21;
  wire [0:0] u_csamul_cska32_fa20_21_xor1;
  wire [0:0] u_csamul_cska32_fa20_21_or0;
  wire [0:0] u_csamul_cska32_and21_21;
  wire [0:0] u_csamul_cska32_fa21_21_xor1;
  wire [0:0] u_csamul_cska32_fa21_21_or0;
  wire [0:0] u_csamul_cska32_and22_21;
  wire [0:0] u_csamul_cska32_fa22_21_xor1;
  wire [0:0] u_csamul_cska32_fa22_21_or0;
  wire [0:0] u_csamul_cska32_and23_21;
  wire [0:0] u_csamul_cska32_fa23_21_xor1;
  wire [0:0] u_csamul_cska32_fa23_21_or0;
  wire [0:0] u_csamul_cska32_and24_21;
  wire [0:0] u_csamul_cska32_fa24_21_xor1;
  wire [0:0] u_csamul_cska32_fa24_21_or0;
  wire [0:0] u_csamul_cska32_and25_21;
  wire [0:0] u_csamul_cska32_fa25_21_xor1;
  wire [0:0] u_csamul_cska32_fa25_21_or0;
  wire [0:0] u_csamul_cska32_and26_21;
  wire [0:0] u_csamul_cska32_fa26_21_xor1;
  wire [0:0] u_csamul_cska32_fa26_21_or0;
  wire [0:0] u_csamul_cska32_and27_21;
  wire [0:0] u_csamul_cska32_fa27_21_xor1;
  wire [0:0] u_csamul_cska32_fa27_21_or0;
  wire [0:0] u_csamul_cska32_and28_21;
  wire [0:0] u_csamul_cska32_fa28_21_xor1;
  wire [0:0] u_csamul_cska32_fa28_21_or0;
  wire [0:0] u_csamul_cska32_and29_21;
  wire [0:0] u_csamul_cska32_fa29_21_xor1;
  wire [0:0] u_csamul_cska32_fa29_21_or0;
  wire [0:0] u_csamul_cska32_and30_21;
  wire [0:0] u_csamul_cska32_fa30_21_xor1;
  wire [0:0] u_csamul_cska32_fa30_21_or0;
  wire [0:0] u_csamul_cska32_and31_21;
  wire [0:0] u_csamul_cska32_and0_22;
  wire [0:0] u_csamul_cska32_fa0_22_xor1;
  wire [0:0] u_csamul_cska32_fa0_22_or0;
  wire [0:0] u_csamul_cska32_and1_22;
  wire [0:0] u_csamul_cska32_fa1_22_xor1;
  wire [0:0] u_csamul_cska32_fa1_22_or0;
  wire [0:0] u_csamul_cska32_and2_22;
  wire [0:0] u_csamul_cska32_fa2_22_xor1;
  wire [0:0] u_csamul_cska32_fa2_22_or0;
  wire [0:0] u_csamul_cska32_and3_22;
  wire [0:0] u_csamul_cska32_fa3_22_xor1;
  wire [0:0] u_csamul_cska32_fa3_22_or0;
  wire [0:0] u_csamul_cska32_and4_22;
  wire [0:0] u_csamul_cska32_fa4_22_xor1;
  wire [0:0] u_csamul_cska32_fa4_22_or0;
  wire [0:0] u_csamul_cska32_and5_22;
  wire [0:0] u_csamul_cska32_fa5_22_xor1;
  wire [0:0] u_csamul_cska32_fa5_22_or0;
  wire [0:0] u_csamul_cska32_and6_22;
  wire [0:0] u_csamul_cska32_fa6_22_xor1;
  wire [0:0] u_csamul_cska32_fa6_22_or0;
  wire [0:0] u_csamul_cska32_and7_22;
  wire [0:0] u_csamul_cska32_fa7_22_xor1;
  wire [0:0] u_csamul_cska32_fa7_22_or0;
  wire [0:0] u_csamul_cska32_and8_22;
  wire [0:0] u_csamul_cska32_fa8_22_xor1;
  wire [0:0] u_csamul_cska32_fa8_22_or0;
  wire [0:0] u_csamul_cska32_and9_22;
  wire [0:0] u_csamul_cska32_fa9_22_xor1;
  wire [0:0] u_csamul_cska32_fa9_22_or0;
  wire [0:0] u_csamul_cska32_and10_22;
  wire [0:0] u_csamul_cska32_fa10_22_xor1;
  wire [0:0] u_csamul_cska32_fa10_22_or0;
  wire [0:0] u_csamul_cska32_and11_22;
  wire [0:0] u_csamul_cska32_fa11_22_xor1;
  wire [0:0] u_csamul_cska32_fa11_22_or0;
  wire [0:0] u_csamul_cska32_and12_22;
  wire [0:0] u_csamul_cska32_fa12_22_xor1;
  wire [0:0] u_csamul_cska32_fa12_22_or0;
  wire [0:0] u_csamul_cska32_and13_22;
  wire [0:0] u_csamul_cska32_fa13_22_xor1;
  wire [0:0] u_csamul_cska32_fa13_22_or0;
  wire [0:0] u_csamul_cska32_and14_22;
  wire [0:0] u_csamul_cska32_fa14_22_xor1;
  wire [0:0] u_csamul_cska32_fa14_22_or0;
  wire [0:0] u_csamul_cska32_and15_22;
  wire [0:0] u_csamul_cska32_fa15_22_xor1;
  wire [0:0] u_csamul_cska32_fa15_22_or0;
  wire [0:0] u_csamul_cska32_and16_22;
  wire [0:0] u_csamul_cska32_fa16_22_xor1;
  wire [0:0] u_csamul_cska32_fa16_22_or0;
  wire [0:0] u_csamul_cska32_and17_22;
  wire [0:0] u_csamul_cska32_fa17_22_xor1;
  wire [0:0] u_csamul_cska32_fa17_22_or0;
  wire [0:0] u_csamul_cska32_and18_22;
  wire [0:0] u_csamul_cska32_fa18_22_xor1;
  wire [0:0] u_csamul_cska32_fa18_22_or0;
  wire [0:0] u_csamul_cska32_and19_22;
  wire [0:0] u_csamul_cska32_fa19_22_xor1;
  wire [0:0] u_csamul_cska32_fa19_22_or0;
  wire [0:0] u_csamul_cska32_and20_22;
  wire [0:0] u_csamul_cska32_fa20_22_xor1;
  wire [0:0] u_csamul_cska32_fa20_22_or0;
  wire [0:0] u_csamul_cska32_and21_22;
  wire [0:0] u_csamul_cska32_fa21_22_xor1;
  wire [0:0] u_csamul_cska32_fa21_22_or0;
  wire [0:0] u_csamul_cska32_and22_22;
  wire [0:0] u_csamul_cska32_fa22_22_xor1;
  wire [0:0] u_csamul_cska32_fa22_22_or0;
  wire [0:0] u_csamul_cska32_and23_22;
  wire [0:0] u_csamul_cska32_fa23_22_xor1;
  wire [0:0] u_csamul_cska32_fa23_22_or0;
  wire [0:0] u_csamul_cska32_and24_22;
  wire [0:0] u_csamul_cska32_fa24_22_xor1;
  wire [0:0] u_csamul_cska32_fa24_22_or0;
  wire [0:0] u_csamul_cska32_and25_22;
  wire [0:0] u_csamul_cska32_fa25_22_xor1;
  wire [0:0] u_csamul_cska32_fa25_22_or0;
  wire [0:0] u_csamul_cska32_and26_22;
  wire [0:0] u_csamul_cska32_fa26_22_xor1;
  wire [0:0] u_csamul_cska32_fa26_22_or0;
  wire [0:0] u_csamul_cska32_and27_22;
  wire [0:0] u_csamul_cska32_fa27_22_xor1;
  wire [0:0] u_csamul_cska32_fa27_22_or0;
  wire [0:0] u_csamul_cska32_and28_22;
  wire [0:0] u_csamul_cska32_fa28_22_xor1;
  wire [0:0] u_csamul_cska32_fa28_22_or0;
  wire [0:0] u_csamul_cska32_and29_22;
  wire [0:0] u_csamul_cska32_fa29_22_xor1;
  wire [0:0] u_csamul_cska32_fa29_22_or0;
  wire [0:0] u_csamul_cska32_and30_22;
  wire [0:0] u_csamul_cska32_fa30_22_xor1;
  wire [0:0] u_csamul_cska32_fa30_22_or0;
  wire [0:0] u_csamul_cska32_and31_22;
  wire [0:0] u_csamul_cska32_and0_23;
  wire [0:0] u_csamul_cska32_fa0_23_xor1;
  wire [0:0] u_csamul_cska32_fa0_23_or0;
  wire [0:0] u_csamul_cska32_and1_23;
  wire [0:0] u_csamul_cska32_fa1_23_xor1;
  wire [0:0] u_csamul_cska32_fa1_23_or0;
  wire [0:0] u_csamul_cska32_and2_23;
  wire [0:0] u_csamul_cska32_fa2_23_xor1;
  wire [0:0] u_csamul_cska32_fa2_23_or0;
  wire [0:0] u_csamul_cska32_and3_23;
  wire [0:0] u_csamul_cska32_fa3_23_xor1;
  wire [0:0] u_csamul_cska32_fa3_23_or0;
  wire [0:0] u_csamul_cska32_and4_23;
  wire [0:0] u_csamul_cska32_fa4_23_xor1;
  wire [0:0] u_csamul_cska32_fa4_23_or0;
  wire [0:0] u_csamul_cska32_and5_23;
  wire [0:0] u_csamul_cska32_fa5_23_xor1;
  wire [0:0] u_csamul_cska32_fa5_23_or0;
  wire [0:0] u_csamul_cska32_and6_23;
  wire [0:0] u_csamul_cska32_fa6_23_xor1;
  wire [0:0] u_csamul_cska32_fa6_23_or0;
  wire [0:0] u_csamul_cska32_and7_23;
  wire [0:0] u_csamul_cska32_fa7_23_xor1;
  wire [0:0] u_csamul_cska32_fa7_23_or0;
  wire [0:0] u_csamul_cska32_and8_23;
  wire [0:0] u_csamul_cska32_fa8_23_xor1;
  wire [0:0] u_csamul_cska32_fa8_23_or0;
  wire [0:0] u_csamul_cska32_and9_23;
  wire [0:0] u_csamul_cska32_fa9_23_xor1;
  wire [0:0] u_csamul_cska32_fa9_23_or0;
  wire [0:0] u_csamul_cska32_and10_23;
  wire [0:0] u_csamul_cska32_fa10_23_xor1;
  wire [0:0] u_csamul_cska32_fa10_23_or0;
  wire [0:0] u_csamul_cska32_and11_23;
  wire [0:0] u_csamul_cska32_fa11_23_xor1;
  wire [0:0] u_csamul_cska32_fa11_23_or0;
  wire [0:0] u_csamul_cska32_and12_23;
  wire [0:0] u_csamul_cska32_fa12_23_xor1;
  wire [0:0] u_csamul_cska32_fa12_23_or0;
  wire [0:0] u_csamul_cska32_and13_23;
  wire [0:0] u_csamul_cska32_fa13_23_xor1;
  wire [0:0] u_csamul_cska32_fa13_23_or0;
  wire [0:0] u_csamul_cska32_and14_23;
  wire [0:0] u_csamul_cska32_fa14_23_xor1;
  wire [0:0] u_csamul_cska32_fa14_23_or0;
  wire [0:0] u_csamul_cska32_and15_23;
  wire [0:0] u_csamul_cska32_fa15_23_xor1;
  wire [0:0] u_csamul_cska32_fa15_23_or0;
  wire [0:0] u_csamul_cska32_and16_23;
  wire [0:0] u_csamul_cska32_fa16_23_xor1;
  wire [0:0] u_csamul_cska32_fa16_23_or0;
  wire [0:0] u_csamul_cska32_and17_23;
  wire [0:0] u_csamul_cska32_fa17_23_xor1;
  wire [0:0] u_csamul_cska32_fa17_23_or0;
  wire [0:0] u_csamul_cska32_and18_23;
  wire [0:0] u_csamul_cska32_fa18_23_xor1;
  wire [0:0] u_csamul_cska32_fa18_23_or0;
  wire [0:0] u_csamul_cska32_and19_23;
  wire [0:0] u_csamul_cska32_fa19_23_xor1;
  wire [0:0] u_csamul_cska32_fa19_23_or0;
  wire [0:0] u_csamul_cska32_and20_23;
  wire [0:0] u_csamul_cska32_fa20_23_xor1;
  wire [0:0] u_csamul_cska32_fa20_23_or0;
  wire [0:0] u_csamul_cska32_and21_23;
  wire [0:0] u_csamul_cska32_fa21_23_xor1;
  wire [0:0] u_csamul_cska32_fa21_23_or0;
  wire [0:0] u_csamul_cska32_and22_23;
  wire [0:0] u_csamul_cska32_fa22_23_xor1;
  wire [0:0] u_csamul_cska32_fa22_23_or0;
  wire [0:0] u_csamul_cska32_and23_23;
  wire [0:0] u_csamul_cska32_fa23_23_xor1;
  wire [0:0] u_csamul_cska32_fa23_23_or0;
  wire [0:0] u_csamul_cska32_and24_23;
  wire [0:0] u_csamul_cska32_fa24_23_xor1;
  wire [0:0] u_csamul_cska32_fa24_23_or0;
  wire [0:0] u_csamul_cska32_and25_23;
  wire [0:0] u_csamul_cska32_fa25_23_xor1;
  wire [0:0] u_csamul_cska32_fa25_23_or0;
  wire [0:0] u_csamul_cska32_and26_23;
  wire [0:0] u_csamul_cska32_fa26_23_xor1;
  wire [0:0] u_csamul_cska32_fa26_23_or0;
  wire [0:0] u_csamul_cska32_and27_23;
  wire [0:0] u_csamul_cska32_fa27_23_xor1;
  wire [0:0] u_csamul_cska32_fa27_23_or0;
  wire [0:0] u_csamul_cska32_and28_23;
  wire [0:0] u_csamul_cska32_fa28_23_xor1;
  wire [0:0] u_csamul_cska32_fa28_23_or0;
  wire [0:0] u_csamul_cska32_and29_23;
  wire [0:0] u_csamul_cska32_fa29_23_xor1;
  wire [0:0] u_csamul_cska32_fa29_23_or0;
  wire [0:0] u_csamul_cska32_and30_23;
  wire [0:0] u_csamul_cska32_fa30_23_xor1;
  wire [0:0] u_csamul_cska32_fa30_23_or0;
  wire [0:0] u_csamul_cska32_and31_23;
  wire [0:0] u_csamul_cska32_and0_24;
  wire [0:0] u_csamul_cska32_fa0_24_xor1;
  wire [0:0] u_csamul_cska32_fa0_24_or0;
  wire [0:0] u_csamul_cska32_and1_24;
  wire [0:0] u_csamul_cska32_fa1_24_xor1;
  wire [0:0] u_csamul_cska32_fa1_24_or0;
  wire [0:0] u_csamul_cska32_and2_24;
  wire [0:0] u_csamul_cska32_fa2_24_xor1;
  wire [0:0] u_csamul_cska32_fa2_24_or0;
  wire [0:0] u_csamul_cska32_and3_24;
  wire [0:0] u_csamul_cska32_fa3_24_xor1;
  wire [0:0] u_csamul_cska32_fa3_24_or0;
  wire [0:0] u_csamul_cska32_and4_24;
  wire [0:0] u_csamul_cska32_fa4_24_xor1;
  wire [0:0] u_csamul_cska32_fa4_24_or0;
  wire [0:0] u_csamul_cska32_and5_24;
  wire [0:0] u_csamul_cska32_fa5_24_xor1;
  wire [0:0] u_csamul_cska32_fa5_24_or0;
  wire [0:0] u_csamul_cska32_and6_24;
  wire [0:0] u_csamul_cska32_fa6_24_xor1;
  wire [0:0] u_csamul_cska32_fa6_24_or0;
  wire [0:0] u_csamul_cska32_and7_24;
  wire [0:0] u_csamul_cska32_fa7_24_xor1;
  wire [0:0] u_csamul_cska32_fa7_24_or0;
  wire [0:0] u_csamul_cska32_and8_24;
  wire [0:0] u_csamul_cska32_fa8_24_xor1;
  wire [0:0] u_csamul_cska32_fa8_24_or0;
  wire [0:0] u_csamul_cska32_and9_24;
  wire [0:0] u_csamul_cska32_fa9_24_xor1;
  wire [0:0] u_csamul_cska32_fa9_24_or0;
  wire [0:0] u_csamul_cska32_and10_24;
  wire [0:0] u_csamul_cska32_fa10_24_xor1;
  wire [0:0] u_csamul_cska32_fa10_24_or0;
  wire [0:0] u_csamul_cska32_and11_24;
  wire [0:0] u_csamul_cska32_fa11_24_xor1;
  wire [0:0] u_csamul_cska32_fa11_24_or0;
  wire [0:0] u_csamul_cska32_and12_24;
  wire [0:0] u_csamul_cska32_fa12_24_xor1;
  wire [0:0] u_csamul_cska32_fa12_24_or0;
  wire [0:0] u_csamul_cska32_and13_24;
  wire [0:0] u_csamul_cska32_fa13_24_xor1;
  wire [0:0] u_csamul_cska32_fa13_24_or0;
  wire [0:0] u_csamul_cska32_and14_24;
  wire [0:0] u_csamul_cska32_fa14_24_xor1;
  wire [0:0] u_csamul_cska32_fa14_24_or0;
  wire [0:0] u_csamul_cska32_and15_24;
  wire [0:0] u_csamul_cska32_fa15_24_xor1;
  wire [0:0] u_csamul_cska32_fa15_24_or0;
  wire [0:0] u_csamul_cska32_and16_24;
  wire [0:0] u_csamul_cska32_fa16_24_xor1;
  wire [0:0] u_csamul_cska32_fa16_24_or0;
  wire [0:0] u_csamul_cska32_and17_24;
  wire [0:0] u_csamul_cska32_fa17_24_xor1;
  wire [0:0] u_csamul_cska32_fa17_24_or0;
  wire [0:0] u_csamul_cska32_and18_24;
  wire [0:0] u_csamul_cska32_fa18_24_xor1;
  wire [0:0] u_csamul_cska32_fa18_24_or0;
  wire [0:0] u_csamul_cska32_and19_24;
  wire [0:0] u_csamul_cska32_fa19_24_xor1;
  wire [0:0] u_csamul_cska32_fa19_24_or0;
  wire [0:0] u_csamul_cska32_and20_24;
  wire [0:0] u_csamul_cska32_fa20_24_xor1;
  wire [0:0] u_csamul_cska32_fa20_24_or0;
  wire [0:0] u_csamul_cska32_and21_24;
  wire [0:0] u_csamul_cska32_fa21_24_xor1;
  wire [0:0] u_csamul_cska32_fa21_24_or0;
  wire [0:0] u_csamul_cska32_and22_24;
  wire [0:0] u_csamul_cska32_fa22_24_xor1;
  wire [0:0] u_csamul_cska32_fa22_24_or0;
  wire [0:0] u_csamul_cska32_and23_24;
  wire [0:0] u_csamul_cska32_fa23_24_xor1;
  wire [0:0] u_csamul_cska32_fa23_24_or0;
  wire [0:0] u_csamul_cska32_and24_24;
  wire [0:0] u_csamul_cska32_fa24_24_xor1;
  wire [0:0] u_csamul_cska32_fa24_24_or0;
  wire [0:0] u_csamul_cska32_and25_24;
  wire [0:0] u_csamul_cska32_fa25_24_xor1;
  wire [0:0] u_csamul_cska32_fa25_24_or0;
  wire [0:0] u_csamul_cska32_and26_24;
  wire [0:0] u_csamul_cska32_fa26_24_xor1;
  wire [0:0] u_csamul_cska32_fa26_24_or0;
  wire [0:0] u_csamul_cska32_and27_24;
  wire [0:0] u_csamul_cska32_fa27_24_xor1;
  wire [0:0] u_csamul_cska32_fa27_24_or0;
  wire [0:0] u_csamul_cska32_and28_24;
  wire [0:0] u_csamul_cska32_fa28_24_xor1;
  wire [0:0] u_csamul_cska32_fa28_24_or0;
  wire [0:0] u_csamul_cska32_and29_24;
  wire [0:0] u_csamul_cska32_fa29_24_xor1;
  wire [0:0] u_csamul_cska32_fa29_24_or0;
  wire [0:0] u_csamul_cska32_and30_24;
  wire [0:0] u_csamul_cska32_fa30_24_xor1;
  wire [0:0] u_csamul_cska32_fa30_24_or0;
  wire [0:0] u_csamul_cska32_and31_24;
  wire [0:0] u_csamul_cska32_and0_25;
  wire [0:0] u_csamul_cska32_fa0_25_xor1;
  wire [0:0] u_csamul_cska32_fa0_25_or0;
  wire [0:0] u_csamul_cska32_and1_25;
  wire [0:0] u_csamul_cska32_fa1_25_xor1;
  wire [0:0] u_csamul_cska32_fa1_25_or0;
  wire [0:0] u_csamul_cska32_and2_25;
  wire [0:0] u_csamul_cska32_fa2_25_xor1;
  wire [0:0] u_csamul_cska32_fa2_25_or0;
  wire [0:0] u_csamul_cska32_and3_25;
  wire [0:0] u_csamul_cska32_fa3_25_xor1;
  wire [0:0] u_csamul_cska32_fa3_25_or0;
  wire [0:0] u_csamul_cska32_and4_25;
  wire [0:0] u_csamul_cska32_fa4_25_xor1;
  wire [0:0] u_csamul_cska32_fa4_25_or0;
  wire [0:0] u_csamul_cska32_and5_25;
  wire [0:0] u_csamul_cska32_fa5_25_xor1;
  wire [0:0] u_csamul_cska32_fa5_25_or0;
  wire [0:0] u_csamul_cska32_and6_25;
  wire [0:0] u_csamul_cska32_fa6_25_xor1;
  wire [0:0] u_csamul_cska32_fa6_25_or0;
  wire [0:0] u_csamul_cska32_and7_25;
  wire [0:0] u_csamul_cska32_fa7_25_xor1;
  wire [0:0] u_csamul_cska32_fa7_25_or0;
  wire [0:0] u_csamul_cska32_and8_25;
  wire [0:0] u_csamul_cska32_fa8_25_xor1;
  wire [0:0] u_csamul_cska32_fa8_25_or0;
  wire [0:0] u_csamul_cska32_and9_25;
  wire [0:0] u_csamul_cska32_fa9_25_xor1;
  wire [0:0] u_csamul_cska32_fa9_25_or0;
  wire [0:0] u_csamul_cska32_and10_25;
  wire [0:0] u_csamul_cska32_fa10_25_xor1;
  wire [0:0] u_csamul_cska32_fa10_25_or0;
  wire [0:0] u_csamul_cska32_and11_25;
  wire [0:0] u_csamul_cska32_fa11_25_xor1;
  wire [0:0] u_csamul_cska32_fa11_25_or0;
  wire [0:0] u_csamul_cska32_and12_25;
  wire [0:0] u_csamul_cska32_fa12_25_xor1;
  wire [0:0] u_csamul_cska32_fa12_25_or0;
  wire [0:0] u_csamul_cska32_and13_25;
  wire [0:0] u_csamul_cska32_fa13_25_xor1;
  wire [0:0] u_csamul_cska32_fa13_25_or0;
  wire [0:0] u_csamul_cska32_and14_25;
  wire [0:0] u_csamul_cska32_fa14_25_xor1;
  wire [0:0] u_csamul_cska32_fa14_25_or0;
  wire [0:0] u_csamul_cska32_and15_25;
  wire [0:0] u_csamul_cska32_fa15_25_xor1;
  wire [0:0] u_csamul_cska32_fa15_25_or0;
  wire [0:0] u_csamul_cska32_and16_25;
  wire [0:0] u_csamul_cska32_fa16_25_xor1;
  wire [0:0] u_csamul_cska32_fa16_25_or0;
  wire [0:0] u_csamul_cska32_and17_25;
  wire [0:0] u_csamul_cska32_fa17_25_xor1;
  wire [0:0] u_csamul_cska32_fa17_25_or0;
  wire [0:0] u_csamul_cska32_and18_25;
  wire [0:0] u_csamul_cska32_fa18_25_xor1;
  wire [0:0] u_csamul_cska32_fa18_25_or0;
  wire [0:0] u_csamul_cska32_and19_25;
  wire [0:0] u_csamul_cska32_fa19_25_xor1;
  wire [0:0] u_csamul_cska32_fa19_25_or0;
  wire [0:0] u_csamul_cska32_and20_25;
  wire [0:0] u_csamul_cska32_fa20_25_xor1;
  wire [0:0] u_csamul_cska32_fa20_25_or0;
  wire [0:0] u_csamul_cska32_and21_25;
  wire [0:0] u_csamul_cska32_fa21_25_xor1;
  wire [0:0] u_csamul_cska32_fa21_25_or0;
  wire [0:0] u_csamul_cska32_and22_25;
  wire [0:0] u_csamul_cska32_fa22_25_xor1;
  wire [0:0] u_csamul_cska32_fa22_25_or0;
  wire [0:0] u_csamul_cska32_and23_25;
  wire [0:0] u_csamul_cska32_fa23_25_xor1;
  wire [0:0] u_csamul_cska32_fa23_25_or0;
  wire [0:0] u_csamul_cska32_and24_25;
  wire [0:0] u_csamul_cska32_fa24_25_xor1;
  wire [0:0] u_csamul_cska32_fa24_25_or0;
  wire [0:0] u_csamul_cska32_and25_25;
  wire [0:0] u_csamul_cska32_fa25_25_xor1;
  wire [0:0] u_csamul_cska32_fa25_25_or0;
  wire [0:0] u_csamul_cska32_and26_25;
  wire [0:0] u_csamul_cska32_fa26_25_xor1;
  wire [0:0] u_csamul_cska32_fa26_25_or0;
  wire [0:0] u_csamul_cska32_and27_25;
  wire [0:0] u_csamul_cska32_fa27_25_xor1;
  wire [0:0] u_csamul_cska32_fa27_25_or0;
  wire [0:0] u_csamul_cska32_and28_25;
  wire [0:0] u_csamul_cska32_fa28_25_xor1;
  wire [0:0] u_csamul_cska32_fa28_25_or0;
  wire [0:0] u_csamul_cska32_and29_25;
  wire [0:0] u_csamul_cska32_fa29_25_xor1;
  wire [0:0] u_csamul_cska32_fa29_25_or0;
  wire [0:0] u_csamul_cska32_and30_25;
  wire [0:0] u_csamul_cska32_fa30_25_xor1;
  wire [0:0] u_csamul_cska32_fa30_25_or0;
  wire [0:0] u_csamul_cska32_and31_25;
  wire [0:0] u_csamul_cska32_and0_26;
  wire [0:0] u_csamul_cska32_fa0_26_xor1;
  wire [0:0] u_csamul_cska32_fa0_26_or0;
  wire [0:0] u_csamul_cska32_and1_26;
  wire [0:0] u_csamul_cska32_fa1_26_xor1;
  wire [0:0] u_csamul_cska32_fa1_26_or0;
  wire [0:0] u_csamul_cska32_and2_26;
  wire [0:0] u_csamul_cska32_fa2_26_xor1;
  wire [0:0] u_csamul_cska32_fa2_26_or0;
  wire [0:0] u_csamul_cska32_and3_26;
  wire [0:0] u_csamul_cska32_fa3_26_xor1;
  wire [0:0] u_csamul_cska32_fa3_26_or0;
  wire [0:0] u_csamul_cska32_and4_26;
  wire [0:0] u_csamul_cska32_fa4_26_xor1;
  wire [0:0] u_csamul_cska32_fa4_26_or0;
  wire [0:0] u_csamul_cska32_and5_26;
  wire [0:0] u_csamul_cska32_fa5_26_xor1;
  wire [0:0] u_csamul_cska32_fa5_26_or0;
  wire [0:0] u_csamul_cska32_and6_26;
  wire [0:0] u_csamul_cska32_fa6_26_xor1;
  wire [0:0] u_csamul_cska32_fa6_26_or0;
  wire [0:0] u_csamul_cska32_and7_26;
  wire [0:0] u_csamul_cska32_fa7_26_xor1;
  wire [0:0] u_csamul_cska32_fa7_26_or0;
  wire [0:0] u_csamul_cska32_and8_26;
  wire [0:0] u_csamul_cska32_fa8_26_xor1;
  wire [0:0] u_csamul_cska32_fa8_26_or0;
  wire [0:0] u_csamul_cska32_and9_26;
  wire [0:0] u_csamul_cska32_fa9_26_xor1;
  wire [0:0] u_csamul_cska32_fa9_26_or0;
  wire [0:0] u_csamul_cska32_and10_26;
  wire [0:0] u_csamul_cska32_fa10_26_xor1;
  wire [0:0] u_csamul_cska32_fa10_26_or0;
  wire [0:0] u_csamul_cska32_and11_26;
  wire [0:0] u_csamul_cska32_fa11_26_xor1;
  wire [0:0] u_csamul_cska32_fa11_26_or0;
  wire [0:0] u_csamul_cska32_and12_26;
  wire [0:0] u_csamul_cska32_fa12_26_xor1;
  wire [0:0] u_csamul_cska32_fa12_26_or0;
  wire [0:0] u_csamul_cska32_and13_26;
  wire [0:0] u_csamul_cska32_fa13_26_xor1;
  wire [0:0] u_csamul_cska32_fa13_26_or0;
  wire [0:0] u_csamul_cska32_and14_26;
  wire [0:0] u_csamul_cska32_fa14_26_xor1;
  wire [0:0] u_csamul_cska32_fa14_26_or0;
  wire [0:0] u_csamul_cska32_and15_26;
  wire [0:0] u_csamul_cska32_fa15_26_xor1;
  wire [0:0] u_csamul_cska32_fa15_26_or0;
  wire [0:0] u_csamul_cska32_and16_26;
  wire [0:0] u_csamul_cska32_fa16_26_xor1;
  wire [0:0] u_csamul_cska32_fa16_26_or0;
  wire [0:0] u_csamul_cska32_and17_26;
  wire [0:0] u_csamul_cska32_fa17_26_xor1;
  wire [0:0] u_csamul_cska32_fa17_26_or0;
  wire [0:0] u_csamul_cska32_and18_26;
  wire [0:0] u_csamul_cska32_fa18_26_xor1;
  wire [0:0] u_csamul_cska32_fa18_26_or0;
  wire [0:0] u_csamul_cska32_and19_26;
  wire [0:0] u_csamul_cska32_fa19_26_xor1;
  wire [0:0] u_csamul_cska32_fa19_26_or0;
  wire [0:0] u_csamul_cska32_and20_26;
  wire [0:0] u_csamul_cska32_fa20_26_xor1;
  wire [0:0] u_csamul_cska32_fa20_26_or0;
  wire [0:0] u_csamul_cska32_and21_26;
  wire [0:0] u_csamul_cska32_fa21_26_xor1;
  wire [0:0] u_csamul_cska32_fa21_26_or0;
  wire [0:0] u_csamul_cska32_and22_26;
  wire [0:0] u_csamul_cska32_fa22_26_xor1;
  wire [0:0] u_csamul_cska32_fa22_26_or0;
  wire [0:0] u_csamul_cska32_and23_26;
  wire [0:0] u_csamul_cska32_fa23_26_xor1;
  wire [0:0] u_csamul_cska32_fa23_26_or0;
  wire [0:0] u_csamul_cska32_and24_26;
  wire [0:0] u_csamul_cska32_fa24_26_xor1;
  wire [0:0] u_csamul_cska32_fa24_26_or0;
  wire [0:0] u_csamul_cska32_and25_26;
  wire [0:0] u_csamul_cska32_fa25_26_xor1;
  wire [0:0] u_csamul_cska32_fa25_26_or0;
  wire [0:0] u_csamul_cska32_and26_26;
  wire [0:0] u_csamul_cska32_fa26_26_xor1;
  wire [0:0] u_csamul_cska32_fa26_26_or0;
  wire [0:0] u_csamul_cska32_and27_26;
  wire [0:0] u_csamul_cska32_fa27_26_xor1;
  wire [0:0] u_csamul_cska32_fa27_26_or0;
  wire [0:0] u_csamul_cska32_and28_26;
  wire [0:0] u_csamul_cska32_fa28_26_xor1;
  wire [0:0] u_csamul_cska32_fa28_26_or0;
  wire [0:0] u_csamul_cska32_and29_26;
  wire [0:0] u_csamul_cska32_fa29_26_xor1;
  wire [0:0] u_csamul_cska32_fa29_26_or0;
  wire [0:0] u_csamul_cska32_and30_26;
  wire [0:0] u_csamul_cska32_fa30_26_xor1;
  wire [0:0] u_csamul_cska32_fa30_26_or0;
  wire [0:0] u_csamul_cska32_and31_26;
  wire [0:0] u_csamul_cska32_and0_27;
  wire [0:0] u_csamul_cska32_fa0_27_xor1;
  wire [0:0] u_csamul_cska32_fa0_27_or0;
  wire [0:0] u_csamul_cska32_and1_27;
  wire [0:0] u_csamul_cska32_fa1_27_xor1;
  wire [0:0] u_csamul_cska32_fa1_27_or0;
  wire [0:0] u_csamul_cska32_and2_27;
  wire [0:0] u_csamul_cska32_fa2_27_xor1;
  wire [0:0] u_csamul_cska32_fa2_27_or0;
  wire [0:0] u_csamul_cska32_and3_27;
  wire [0:0] u_csamul_cska32_fa3_27_xor1;
  wire [0:0] u_csamul_cska32_fa3_27_or0;
  wire [0:0] u_csamul_cska32_and4_27;
  wire [0:0] u_csamul_cska32_fa4_27_xor1;
  wire [0:0] u_csamul_cska32_fa4_27_or0;
  wire [0:0] u_csamul_cska32_and5_27;
  wire [0:0] u_csamul_cska32_fa5_27_xor1;
  wire [0:0] u_csamul_cska32_fa5_27_or0;
  wire [0:0] u_csamul_cska32_and6_27;
  wire [0:0] u_csamul_cska32_fa6_27_xor1;
  wire [0:0] u_csamul_cska32_fa6_27_or0;
  wire [0:0] u_csamul_cska32_and7_27;
  wire [0:0] u_csamul_cska32_fa7_27_xor1;
  wire [0:0] u_csamul_cska32_fa7_27_or0;
  wire [0:0] u_csamul_cska32_and8_27;
  wire [0:0] u_csamul_cska32_fa8_27_xor1;
  wire [0:0] u_csamul_cska32_fa8_27_or0;
  wire [0:0] u_csamul_cska32_and9_27;
  wire [0:0] u_csamul_cska32_fa9_27_xor1;
  wire [0:0] u_csamul_cska32_fa9_27_or0;
  wire [0:0] u_csamul_cska32_and10_27;
  wire [0:0] u_csamul_cska32_fa10_27_xor1;
  wire [0:0] u_csamul_cska32_fa10_27_or0;
  wire [0:0] u_csamul_cska32_and11_27;
  wire [0:0] u_csamul_cska32_fa11_27_xor1;
  wire [0:0] u_csamul_cska32_fa11_27_or0;
  wire [0:0] u_csamul_cska32_and12_27;
  wire [0:0] u_csamul_cska32_fa12_27_xor1;
  wire [0:0] u_csamul_cska32_fa12_27_or0;
  wire [0:0] u_csamul_cska32_and13_27;
  wire [0:0] u_csamul_cska32_fa13_27_xor1;
  wire [0:0] u_csamul_cska32_fa13_27_or0;
  wire [0:0] u_csamul_cska32_and14_27;
  wire [0:0] u_csamul_cska32_fa14_27_xor1;
  wire [0:0] u_csamul_cska32_fa14_27_or0;
  wire [0:0] u_csamul_cska32_and15_27;
  wire [0:0] u_csamul_cska32_fa15_27_xor1;
  wire [0:0] u_csamul_cska32_fa15_27_or0;
  wire [0:0] u_csamul_cska32_and16_27;
  wire [0:0] u_csamul_cska32_fa16_27_xor1;
  wire [0:0] u_csamul_cska32_fa16_27_or0;
  wire [0:0] u_csamul_cska32_and17_27;
  wire [0:0] u_csamul_cska32_fa17_27_xor1;
  wire [0:0] u_csamul_cska32_fa17_27_or0;
  wire [0:0] u_csamul_cska32_and18_27;
  wire [0:0] u_csamul_cska32_fa18_27_xor1;
  wire [0:0] u_csamul_cska32_fa18_27_or0;
  wire [0:0] u_csamul_cska32_and19_27;
  wire [0:0] u_csamul_cska32_fa19_27_xor1;
  wire [0:0] u_csamul_cska32_fa19_27_or0;
  wire [0:0] u_csamul_cska32_and20_27;
  wire [0:0] u_csamul_cska32_fa20_27_xor1;
  wire [0:0] u_csamul_cska32_fa20_27_or0;
  wire [0:0] u_csamul_cska32_and21_27;
  wire [0:0] u_csamul_cska32_fa21_27_xor1;
  wire [0:0] u_csamul_cska32_fa21_27_or0;
  wire [0:0] u_csamul_cska32_and22_27;
  wire [0:0] u_csamul_cska32_fa22_27_xor1;
  wire [0:0] u_csamul_cska32_fa22_27_or0;
  wire [0:0] u_csamul_cska32_and23_27;
  wire [0:0] u_csamul_cska32_fa23_27_xor1;
  wire [0:0] u_csamul_cska32_fa23_27_or0;
  wire [0:0] u_csamul_cska32_and24_27;
  wire [0:0] u_csamul_cska32_fa24_27_xor1;
  wire [0:0] u_csamul_cska32_fa24_27_or0;
  wire [0:0] u_csamul_cska32_and25_27;
  wire [0:0] u_csamul_cska32_fa25_27_xor1;
  wire [0:0] u_csamul_cska32_fa25_27_or0;
  wire [0:0] u_csamul_cska32_and26_27;
  wire [0:0] u_csamul_cska32_fa26_27_xor1;
  wire [0:0] u_csamul_cska32_fa26_27_or0;
  wire [0:0] u_csamul_cska32_and27_27;
  wire [0:0] u_csamul_cska32_fa27_27_xor1;
  wire [0:0] u_csamul_cska32_fa27_27_or0;
  wire [0:0] u_csamul_cska32_and28_27;
  wire [0:0] u_csamul_cska32_fa28_27_xor1;
  wire [0:0] u_csamul_cska32_fa28_27_or0;
  wire [0:0] u_csamul_cska32_and29_27;
  wire [0:0] u_csamul_cska32_fa29_27_xor1;
  wire [0:0] u_csamul_cska32_fa29_27_or0;
  wire [0:0] u_csamul_cska32_and30_27;
  wire [0:0] u_csamul_cska32_fa30_27_xor1;
  wire [0:0] u_csamul_cska32_fa30_27_or0;
  wire [0:0] u_csamul_cska32_and31_27;
  wire [0:0] u_csamul_cska32_and0_28;
  wire [0:0] u_csamul_cska32_fa0_28_xor1;
  wire [0:0] u_csamul_cska32_fa0_28_or0;
  wire [0:0] u_csamul_cska32_and1_28;
  wire [0:0] u_csamul_cska32_fa1_28_xor1;
  wire [0:0] u_csamul_cska32_fa1_28_or0;
  wire [0:0] u_csamul_cska32_and2_28;
  wire [0:0] u_csamul_cska32_fa2_28_xor1;
  wire [0:0] u_csamul_cska32_fa2_28_or0;
  wire [0:0] u_csamul_cska32_and3_28;
  wire [0:0] u_csamul_cska32_fa3_28_xor1;
  wire [0:0] u_csamul_cska32_fa3_28_or0;
  wire [0:0] u_csamul_cska32_and4_28;
  wire [0:0] u_csamul_cska32_fa4_28_xor1;
  wire [0:0] u_csamul_cska32_fa4_28_or0;
  wire [0:0] u_csamul_cska32_and5_28;
  wire [0:0] u_csamul_cska32_fa5_28_xor1;
  wire [0:0] u_csamul_cska32_fa5_28_or0;
  wire [0:0] u_csamul_cska32_and6_28;
  wire [0:0] u_csamul_cska32_fa6_28_xor1;
  wire [0:0] u_csamul_cska32_fa6_28_or0;
  wire [0:0] u_csamul_cska32_and7_28;
  wire [0:0] u_csamul_cska32_fa7_28_xor1;
  wire [0:0] u_csamul_cska32_fa7_28_or0;
  wire [0:0] u_csamul_cska32_and8_28;
  wire [0:0] u_csamul_cska32_fa8_28_xor1;
  wire [0:0] u_csamul_cska32_fa8_28_or0;
  wire [0:0] u_csamul_cska32_and9_28;
  wire [0:0] u_csamul_cska32_fa9_28_xor1;
  wire [0:0] u_csamul_cska32_fa9_28_or0;
  wire [0:0] u_csamul_cska32_and10_28;
  wire [0:0] u_csamul_cska32_fa10_28_xor1;
  wire [0:0] u_csamul_cska32_fa10_28_or0;
  wire [0:0] u_csamul_cska32_and11_28;
  wire [0:0] u_csamul_cska32_fa11_28_xor1;
  wire [0:0] u_csamul_cska32_fa11_28_or0;
  wire [0:0] u_csamul_cska32_and12_28;
  wire [0:0] u_csamul_cska32_fa12_28_xor1;
  wire [0:0] u_csamul_cska32_fa12_28_or0;
  wire [0:0] u_csamul_cska32_and13_28;
  wire [0:0] u_csamul_cska32_fa13_28_xor1;
  wire [0:0] u_csamul_cska32_fa13_28_or0;
  wire [0:0] u_csamul_cska32_and14_28;
  wire [0:0] u_csamul_cska32_fa14_28_xor1;
  wire [0:0] u_csamul_cska32_fa14_28_or0;
  wire [0:0] u_csamul_cska32_and15_28;
  wire [0:0] u_csamul_cska32_fa15_28_xor1;
  wire [0:0] u_csamul_cska32_fa15_28_or0;
  wire [0:0] u_csamul_cska32_and16_28;
  wire [0:0] u_csamul_cska32_fa16_28_xor1;
  wire [0:0] u_csamul_cska32_fa16_28_or0;
  wire [0:0] u_csamul_cska32_and17_28;
  wire [0:0] u_csamul_cska32_fa17_28_xor1;
  wire [0:0] u_csamul_cska32_fa17_28_or0;
  wire [0:0] u_csamul_cska32_and18_28;
  wire [0:0] u_csamul_cska32_fa18_28_xor1;
  wire [0:0] u_csamul_cska32_fa18_28_or0;
  wire [0:0] u_csamul_cska32_and19_28;
  wire [0:0] u_csamul_cska32_fa19_28_xor1;
  wire [0:0] u_csamul_cska32_fa19_28_or0;
  wire [0:0] u_csamul_cska32_and20_28;
  wire [0:0] u_csamul_cska32_fa20_28_xor1;
  wire [0:0] u_csamul_cska32_fa20_28_or0;
  wire [0:0] u_csamul_cska32_and21_28;
  wire [0:0] u_csamul_cska32_fa21_28_xor1;
  wire [0:0] u_csamul_cska32_fa21_28_or0;
  wire [0:0] u_csamul_cska32_and22_28;
  wire [0:0] u_csamul_cska32_fa22_28_xor1;
  wire [0:0] u_csamul_cska32_fa22_28_or0;
  wire [0:0] u_csamul_cska32_and23_28;
  wire [0:0] u_csamul_cska32_fa23_28_xor1;
  wire [0:0] u_csamul_cska32_fa23_28_or0;
  wire [0:0] u_csamul_cska32_and24_28;
  wire [0:0] u_csamul_cska32_fa24_28_xor1;
  wire [0:0] u_csamul_cska32_fa24_28_or0;
  wire [0:0] u_csamul_cska32_and25_28;
  wire [0:0] u_csamul_cska32_fa25_28_xor1;
  wire [0:0] u_csamul_cska32_fa25_28_or0;
  wire [0:0] u_csamul_cska32_and26_28;
  wire [0:0] u_csamul_cska32_fa26_28_xor1;
  wire [0:0] u_csamul_cska32_fa26_28_or0;
  wire [0:0] u_csamul_cska32_and27_28;
  wire [0:0] u_csamul_cska32_fa27_28_xor1;
  wire [0:0] u_csamul_cska32_fa27_28_or0;
  wire [0:0] u_csamul_cska32_and28_28;
  wire [0:0] u_csamul_cska32_fa28_28_xor1;
  wire [0:0] u_csamul_cska32_fa28_28_or0;
  wire [0:0] u_csamul_cska32_and29_28;
  wire [0:0] u_csamul_cska32_fa29_28_xor1;
  wire [0:0] u_csamul_cska32_fa29_28_or0;
  wire [0:0] u_csamul_cska32_and30_28;
  wire [0:0] u_csamul_cska32_fa30_28_xor1;
  wire [0:0] u_csamul_cska32_fa30_28_or0;
  wire [0:0] u_csamul_cska32_and31_28;
  wire [0:0] u_csamul_cska32_and0_29;
  wire [0:0] u_csamul_cska32_fa0_29_xor1;
  wire [0:0] u_csamul_cska32_fa0_29_or0;
  wire [0:0] u_csamul_cska32_and1_29;
  wire [0:0] u_csamul_cska32_fa1_29_xor1;
  wire [0:0] u_csamul_cska32_fa1_29_or0;
  wire [0:0] u_csamul_cska32_and2_29;
  wire [0:0] u_csamul_cska32_fa2_29_xor1;
  wire [0:0] u_csamul_cska32_fa2_29_or0;
  wire [0:0] u_csamul_cska32_and3_29;
  wire [0:0] u_csamul_cska32_fa3_29_xor1;
  wire [0:0] u_csamul_cska32_fa3_29_or0;
  wire [0:0] u_csamul_cska32_and4_29;
  wire [0:0] u_csamul_cska32_fa4_29_xor1;
  wire [0:0] u_csamul_cska32_fa4_29_or0;
  wire [0:0] u_csamul_cska32_and5_29;
  wire [0:0] u_csamul_cska32_fa5_29_xor1;
  wire [0:0] u_csamul_cska32_fa5_29_or0;
  wire [0:0] u_csamul_cska32_and6_29;
  wire [0:0] u_csamul_cska32_fa6_29_xor1;
  wire [0:0] u_csamul_cska32_fa6_29_or0;
  wire [0:0] u_csamul_cska32_and7_29;
  wire [0:0] u_csamul_cska32_fa7_29_xor1;
  wire [0:0] u_csamul_cska32_fa7_29_or0;
  wire [0:0] u_csamul_cska32_and8_29;
  wire [0:0] u_csamul_cska32_fa8_29_xor1;
  wire [0:0] u_csamul_cska32_fa8_29_or0;
  wire [0:0] u_csamul_cska32_and9_29;
  wire [0:0] u_csamul_cska32_fa9_29_xor1;
  wire [0:0] u_csamul_cska32_fa9_29_or0;
  wire [0:0] u_csamul_cska32_and10_29;
  wire [0:0] u_csamul_cska32_fa10_29_xor1;
  wire [0:0] u_csamul_cska32_fa10_29_or0;
  wire [0:0] u_csamul_cska32_and11_29;
  wire [0:0] u_csamul_cska32_fa11_29_xor1;
  wire [0:0] u_csamul_cska32_fa11_29_or0;
  wire [0:0] u_csamul_cska32_and12_29;
  wire [0:0] u_csamul_cska32_fa12_29_xor1;
  wire [0:0] u_csamul_cska32_fa12_29_or0;
  wire [0:0] u_csamul_cska32_and13_29;
  wire [0:0] u_csamul_cska32_fa13_29_xor1;
  wire [0:0] u_csamul_cska32_fa13_29_or0;
  wire [0:0] u_csamul_cska32_and14_29;
  wire [0:0] u_csamul_cska32_fa14_29_xor1;
  wire [0:0] u_csamul_cska32_fa14_29_or0;
  wire [0:0] u_csamul_cska32_and15_29;
  wire [0:0] u_csamul_cska32_fa15_29_xor1;
  wire [0:0] u_csamul_cska32_fa15_29_or0;
  wire [0:0] u_csamul_cska32_and16_29;
  wire [0:0] u_csamul_cska32_fa16_29_xor1;
  wire [0:0] u_csamul_cska32_fa16_29_or0;
  wire [0:0] u_csamul_cska32_and17_29;
  wire [0:0] u_csamul_cska32_fa17_29_xor1;
  wire [0:0] u_csamul_cska32_fa17_29_or0;
  wire [0:0] u_csamul_cska32_and18_29;
  wire [0:0] u_csamul_cska32_fa18_29_xor1;
  wire [0:0] u_csamul_cska32_fa18_29_or0;
  wire [0:0] u_csamul_cska32_and19_29;
  wire [0:0] u_csamul_cska32_fa19_29_xor1;
  wire [0:0] u_csamul_cska32_fa19_29_or0;
  wire [0:0] u_csamul_cska32_and20_29;
  wire [0:0] u_csamul_cska32_fa20_29_xor1;
  wire [0:0] u_csamul_cska32_fa20_29_or0;
  wire [0:0] u_csamul_cska32_and21_29;
  wire [0:0] u_csamul_cska32_fa21_29_xor1;
  wire [0:0] u_csamul_cska32_fa21_29_or0;
  wire [0:0] u_csamul_cska32_and22_29;
  wire [0:0] u_csamul_cska32_fa22_29_xor1;
  wire [0:0] u_csamul_cska32_fa22_29_or0;
  wire [0:0] u_csamul_cska32_and23_29;
  wire [0:0] u_csamul_cska32_fa23_29_xor1;
  wire [0:0] u_csamul_cska32_fa23_29_or0;
  wire [0:0] u_csamul_cska32_and24_29;
  wire [0:0] u_csamul_cska32_fa24_29_xor1;
  wire [0:0] u_csamul_cska32_fa24_29_or0;
  wire [0:0] u_csamul_cska32_and25_29;
  wire [0:0] u_csamul_cska32_fa25_29_xor1;
  wire [0:0] u_csamul_cska32_fa25_29_or0;
  wire [0:0] u_csamul_cska32_and26_29;
  wire [0:0] u_csamul_cska32_fa26_29_xor1;
  wire [0:0] u_csamul_cska32_fa26_29_or0;
  wire [0:0] u_csamul_cska32_and27_29;
  wire [0:0] u_csamul_cska32_fa27_29_xor1;
  wire [0:0] u_csamul_cska32_fa27_29_or0;
  wire [0:0] u_csamul_cska32_and28_29;
  wire [0:0] u_csamul_cska32_fa28_29_xor1;
  wire [0:0] u_csamul_cska32_fa28_29_or0;
  wire [0:0] u_csamul_cska32_and29_29;
  wire [0:0] u_csamul_cska32_fa29_29_xor1;
  wire [0:0] u_csamul_cska32_fa29_29_or0;
  wire [0:0] u_csamul_cska32_and30_29;
  wire [0:0] u_csamul_cska32_fa30_29_xor1;
  wire [0:0] u_csamul_cska32_fa30_29_or0;
  wire [0:0] u_csamul_cska32_and31_29;
  wire [0:0] u_csamul_cska32_and0_30;
  wire [0:0] u_csamul_cska32_fa0_30_xor1;
  wire [0:0] u_csamul_cska32_fa0_30_or0;
  wire [0:0] u_csamul_cska32_and1_30;
  wire [0:0] u_csamul_cska32_fa1_30_xor1;
  wire [0:0] u_csamul_cska32_fa1_30_or0;
  wire [0:0] u_csamul_cska32_and2_30;
  wire [0:0] u_csamul_cska32_fa2_30_xor1;
  wire [0:0] u_csamul_cska32_fa2_30_or0;
  wire [0:0] u_csamul_cska32_and3_30;
  wire [0:0] u_csamul_cska32_fa3_30_xor1;
  wire [0:0] u_csamul_cska32_fa3_30_or0;
  wire [0:0] u_csamul_cska32_and4_30;
  wire [0:0] u_csamul_cska32_fa4_30_xor1;
  wire [0:0] u_csamul_cska32_fa4_30_or0;
  wire [0:0] u_csamul_cska32_and5_30;
  wire [0:0] u_csamul_cska32_fa5_30_xor1;
  wire [0:0] u_csamul_cska32_fa5_30_or0;
  wire [0:0] u_csamul_cska32_and6_30;
  wire [0:0] u_csamul_cska32_fa6_30_xor1;
  wire [0:0] u_csamul_cska32_fa6_30_or0;
  wire [0:0] u_csamul_cska32_and7_30;
  wire [0:0] u_csamul_cska32_fa7_30_xor1;
  wire [0:0] u_csamul_cska32_fa7_30_or0;
  wire [0:0] u_csamul_cska32_and8_30;
  wire [0:0] u_csamul_cska32_fa8_30_xor1;
  wire [0:0] u_csamul_cska32_fa8_30_or0;
  wire [0:0] u_csamul_cska32_and9_30;
  wire [0:0] u_csamul_cska32_fa9_30_xor1;
  wire [0:0] u_csamul_cska32_fa9_30_or0;
  wire [0:0] u_csamul_cska32_and10_30;
  wire [0:0] u_csamul_cska32_fa10_30_xor1;
  wire [0:0] u_csamul_cska32_fa10_30_or0;
  wire [0:0] u_csamul_cska32_and11_30;
  wire [0:0] u_csamul_cska32_fa11_30_xor1;
  wire [0:0] u_csamul_cska32_fa11_30_or0;
  wire [0:0] u_csamul_cska32_and12_30;
  wire [0:0] u_csamul_cska32_fa12_30_xor1;
  wire [0:0] u_csamul_cska32_fa12_30_or0;
  wire [0:0] u_csamul_cska32_and13_30;
  wire [0:0] u_csamul_cska32_fa13_30_xor1;
  wire [0:0] u_csamul_cska32_fa13_30_or0;
  wire [0:0] u_csamul_cska32_and14_30;
  wire [0:0] u_csamul_cska32_fa14_30_xor1;
  wire [0:0] u_csamul_cska32_fa14_30_or0;
  wire [0:0] u_csamul_cska32_and15_30;
  wire [0:0] u_csamul_cska32_fa15_30_xor1;
  wire [0:0] u_csamul_cska32_fa15_30_or0;
  wire [0:0] u_csamul_cska32_and16_30;
  wire [0:0] u_csamul_cska32_fa16_30_xor1;
  wire [0:0] u_csamul_cska32_fa16_30_or0;
  wire [0:0] u_csamul_cska32_and17_30;
  wire [0:0] u_csamul_cska32_fa17_30_xor1;
  wire [0:0] u_csamul_cska32_fa17_30_or0;
  wire [0:0] u_csamul_cska32_and18_30;
  wire [0:0] u_csamul_cska32_fa18_30_xor1;
  wire [0:0] u_csamul_cska32_fa18_30_or0;
  wire [0:0] u_csamul_cska32_and19_30;
  wire [0:0] u_csamul_cska32_fa19_30_xor1;
  wire [0:0] u_csamul_cska32_fa19_30_or0;
  wire [0:0] u_csamul_cska32_and20_30;
  wire [0:0] u_csamul_cska32_fa20_30_xor1;
  wire [0:0] u_csamul_cska32_fa20_30_or0;
  wire [0:0] u_csamul_cska32_and21_30;
  wire [0:0] u_csamul_cska32_fa21_30_xor1;
  wire [0:0] u_csamul_cska32_fa21_30_or0;
  wire [0:0] u_csamul_cska32_and22_30;
  wire [0:0] u_csamul_cska32_fa22_30_xor1;
  wire [0:0] u_csamul_cska32_fa22_30_or0;
  wire [0:0] u_csamul_cska32_and23_30;
  wire [0:0] u_csamul_cska32_fa23_30_xor1;
  wire [0:0] u_csamul_cska32_fa23_30_or0;
  wire [0:0] u_csamul_cska32_and24_30;
  wire [0:0] u_csamul_cska32_fa24_30_xor1;
  wire [0:0] u_csamul_cska32_fa24_30_or0;
  wire [0:0] u_csamul_cska32_and25_30;
  wire [0:0] u_csamul_cska32_fa25_30_xor1;
  wire [0:0] u_csamul_cska32_fa25_30_or0;
  wire [0:0] u_csamul_cska32_and26_30;
  wire [0:0] u_csamul_cska32_fa26_30_xor1;
  wire [0:0] u_csamul_cska32_fa26_30_or0;
  wire [0:0] u_csamul_cska32_and27_30;
  wire [0:0] u_csamul_cska32_fa27_30_xor1;
  wire [0:0] u_csamul_cska32_fa27_30_or0;
  wire [0:0] u_csamul_cska32_and28_30;
  wire [0:0] u_csamul_cska32_fa28_30_xor1;
  wire [0:0] u_csamul_cska32_fa28_30_or0;
  wire [0:0] u_csamul_cska32_and29_30;
  wire [0:0] u_csamul_cska32_fa29_30_xor1;
  wire [0:0] u_csamul_cska32_fa29_30_or0;
  wire [0:0] u_csamul_cska32_and30_30;
  wire [0:0] u_csamul_cska32_fa30_30_xor1;
  wire [0:0] u_csamul_cska32_fa30_30_or0;
  wire [0:0] u_csamul_cska32_and31_30;
  wire [0:0] u_csamul_cska32_and0_31;
  wire [0:0] u_csamul_cska32_fa0_31_xor1;
  wire [0:0] u_csamul_cska32_fa0_31_or0;
  wire [0:0] u_csamul_cska32_and1_31;
  wire [0:0] u_csamul_cska32_fa1_31_xor1;
  wire [0:0] u_csamul_cska32_fa1_31_or0;
  wire [0:0] u_csamul_cska32_and2_31;
  wire [0:0] u_csamul_cska32_fa2_31_xor1;
  wire [0:0] u_csamul_cska32_fa2_31_or0;
  wire [0:0] u_csamul_cska32_and3_31;
  wire [0:0] u_csamul_cska32_fa3_31_xor1;
  wire [0:0] u_csamul_cska32_fa3_31_or0;
  wire [0:0] u_csamul_cska32_and4_31;
  wire [0:0] u_csamul_cska32_fa4_31_xor1;
  wire [0:0] u_csamul_cska32_fa4_31_or0;
  wire [0:0] u_csamul_cska32_and5_31;
  wire [0:0] u_csamul_cska32_fa5_31_xor1;
  wire [0:0] u_csamul_cska32_fa5_31_or0;
  wire [0:0] u_csamul_cska32_and6_31;
  wire [0:0] u_csamul_cska32_fa6_31_xor1;
  wire [0:0] u_csamul_cska32_fa6_31_or0;
  wire [0:0] u_csamul_cska32_and7_31;
  wire [0:0] u_csamul_cska32_fa7_31_xor1;
  wire [0:0] u_csamul_cska32_fa7_31_or0;
  wire [0:0] u_csamul_cska32_and8_31;
  wire [0:0] u_csamul_cska32_fa8_31_xor1;
  wire [0:0] u_csamul_cska32_fa8_31_or0;
  wire [0:0] u_csamul_cska32_and9_31;
  wire [0:0] u_csamul_cska32_fa9_31_xor1;
  wire [0:0] u_csamul_cska32_fa9_31_or0;
  wire [0:0] u_csamul_cska32_and10_31;
  wire [0:0] u_csamul_cska32_fa10_31_xor1;
  wire [0:0] u_csamul_cska32_fa10_31_or0;
  wire [0:0] u_csamul_cska32_and11_31;
  wire [0:0] u_csamul_cska32_fa11_31_xor1;
  wire [0:0] u_csamul_cska32_fa11_31_or0;
  wire [0:0] u_csamul_cska32_and12_31;
  wire [0:0] u_csamul_cska32_fa12_31_xor1;
  wire [0:0] u_csamul_cska32_fa12_31_or0;
  wire [0:0] u_csamul_cska32_and13_31;
  wire [0:0] u_csamul_cska32_fa13_31_xor1;
  wire [0:0] u_csamul_cska32_fa13_31_or0;
  wire [0:0] u_csamul_cska32_and14_31;
  wire [0:0] u_csamul_cska32_fa14_31_xor1;
  wire [0:0] u_csamul_cska32_fa14_31_or0;
  wire [0:0] u_csamul_cska32_and15_31;
  wire [0:0] u_csamul_cska32_fa15_31_xor1;
  wire [0:0] u_csamul_cska32_fa15_31_or0;
  wire [0:0] u_csamul_cska32_and16_31;
  wire [0:0] u_csamul_cska32_fa16_31_xor1;
  wire [0:0] u_csamul_cska32_fa16_31_or0;
  wire [0:0] u_csamul_cska32_and17_31;
  wire [0:0] u_csamul_cska32_fa17_31_xor1;
  wire [0:0] u_csamul_cska32_fa17_31_or0;
  wire [0:0] u_csamul_cska32_and18_31;
  wire [0:0] u_csamul_cska32_fa18_31_xor1;
  wire [0:0] u_csamul_cska32_fa18_31_or0;
  wire [0:0] u_csamul_cska32_and19_31;
  wire [0:0] u_csamul_cska32_fa19_31_xor1;
  wire [0:0] u_csamul_cska32_fa19_31_or0;
  wire [0:0] u_csamul_cska32_and20_31;
  wire [0:0] u_csamul_cska32_fa20_31_xor1;
  wire [0:0] u_csamul_cska32_fa20_31_or0;
  wire [0:0] u_csamul_cska32_and21_31;
  wire [0:0] u_csamul_cska32_fa21_31_xor1;
  wire [0:0] u_csamul_cska32_fa21_31_or0;
  wire [0:0] u_csamul_cska32_and22_31;
  wire [0:0] u_csamul_cska32_fa22_31_xor1;
  wire [0:0] u_csamul_cska32_fa22_31_or0;
  wire [0:0] u_csamul_cska32_and23_31;
  wire [0:0] u_csamul_cska32_fa23_31_xor1;
  wire [0:0] u_csamul_cska32_fa23_31_or0;
  wire [0:0] u_csamul_cska32_and24_31;
  wire [0:0] u_csamul_cska32_fa24_31_xor1;
  wire [0:0] u_csamul_cska32_fa24_31_or0;
  wire [0:0] u_csamul_cska32_and25_31;
  wire [0:0] u_csamul_cska32_fa25_31_xor1;
  wire [0:0] u_csamul_cska32_fa25_31_or0;
  wire [0:0] u_csamul_cska32_and26_31;
  wire [0:0] u_csamul_cska32_fa26_31_xor1;
  wire [0:0] u_csamul_cska32_fa26_31_or0;
  wire [0:0] u_csamul_cska32_and27_31;
  wire [0:0] u_csamul_cska32_fa27_31_xor1;
  wire [0:0] u_csamul_cska32_fa27_31_or0;
  wire [0:0] u_csamul_cska32_and28_31;
  wire [0:0] u_csamul_cska32_fa28_31_xor1;
  wire [0:0] u_csamul_cska32_fa28_31_or0;
  wire [0:0] u_csamul_cska32_and29_31;
  wire [0:0] u_csamul_cska32_fa29_31_xor1;
  wire [0:0] u_csamul_cska32_fa29_31_or0;
  wire [0:0] u_csamul_cska32_and30_31;
  wire [0:0] u_csamul_cska32_fa30_31_xor1;
  wire [0:0] u_csamul_cska32_fa30_31_or0;
  wire [0:0] u_csamul_cska32_and31_31;
  wire [31:0] u_csamul_cska32_u_cska32_a;
  wire [31:0] u_csamul_cska32_u_cska32_b;
  wire [32:0] u_csamul_cska32_u_cska32_out;

  and_gate and_gate_u_csamul_cska32_and0_0(.a(a[0]), .b(b[0]), .out(u_csamul_cska32_and0_0));
  and_gate and_gate_u_csamul_cska32_and1_0(.a(a[1]), .b(b[0]), .out(u_csamul_cska32_and1_0));
  and_gate and_gate_u_csamul_cska32_and2_0(.a(a[2]), .b(b[0]), .out(u_csamul_cska32_and2_0));
  and_gate and_gate_u_csamul_cska32_and3_0(.a(a[3]), .b(b[0]), .out(u_csamul_cska32_and3_0));
  and_gate and_gate_u_csamul_cska32_and4_0(.a(a[4]), .b(b[0]), .out(u_csamul_cska32_and4_0));
  and_gate and_gate_u_csamul_cska32_and5_0(.a(a[5]), .b(b[0]), .out(u_csamul_cska32_and5_0));
  and_gate and_gate_u_csamul_cska32_and6_0(.a(a[6]), .b(b[0]), .out(u_csamul_cska32_and6_0));
  and_gate and_gate_u_csamul_cska32_and7_0(.a(a[7]), .b(b[0]), .out(u_csamul_cska32_and7_0));
  and_gate and_gate_u_csamul_cska32_and8_0(.a(a[8]), .b(b[0]), .out(u_csamul_cska32_and8_0));
  and_gate and_gate_u_csamul_cska32_and9_0(.a(a[9]), .b(b[0]), .out(u_csamul_cska32_and9_0));
  and_gate and_gate_u_csamul_cska32_and10_0(.a(a[10]), .b(b[0]), .out(u_csamul_cska32_and10_0));
  and_gate and_gate_u_csamul_cska32_and11_0(.a(a[11]), .b(b[0]), .out(u_csamul_cska32_and11_0));
  and_gate and_gate_u_csamul_cska32_and12_0(.a(a[12]), .b(b[0]), .out(u_csamul_cska32_and12_0));
  and_gate and_gate_u_csamul_cska32_and13_0(.a(a[13]), .b(b[0]), .out(u_csamul_cska32_and13_0));
  and_gate and_gate_u_csamul_cska32_and14_0(.a(a[14]), .b(b[0]), .out(u_csamul_cska32_and14_0));
  and_gate and_gate_u_csamul_cska32_and15_0(.a(a[15]), .b(b[0]), .out(u_csamul_cska32_and15_0));
  and_gate and_gate_u_csamul_cska32_and16_0(.a(a[16]), .b(b[0]), .out(u_csamul_cska32_and16_0));
  and_gate and_gate_u_csamul_cska32_and17_0(.a(a[17]), .b(b[0]), .out(u_csamul_cska32_and17_0));
  and_gate and_gate_u_csamul_cska32_and18_0(.a(a[18]), .b(b[0]), .out(u_csamul_cska32_and18_0));
  and_gate and_gate_u_csamul_cska32_and19_0(.a(a[19]), .b(b[0]), .out(u_csamul_cska32_and19_0));
  and_gate and_gate_u_csamul_cska32_and20_0(.a(a[20]), .b(b[0]), .out(u_csamul_cska32_and20_0));
  and_gate and_gate_u_csamul_cska32_and21_0(.a(a[21]), .b(b[0]), .out(u_csamul_cska32_and21_0));
  and_gate and_gate_u_csamul_cska32_and22_0(.a(a[22]), .b(b[0]), .out(u_csamul_cska32_and22_0));
  and_gate and_gate_u_csamul_cska32_and23_0(.a(a[23]), .b(b[0]), .out(u_csamul_cska32_and23_0));
  and_gate and_gate_u_csamul_cska32_and24_0(.a(a[24]), .b(b[0]), .out(u_csamul_cska32_and24_0));
  and_gate and_gate_u_csamul_cska32_and25_0(.a(a[25]), .b(b[0]), .out(u_csamul_cska32_and25_0));
  and_gate and_gate_u_csamul_cska32_and26_0(.a(a[26]), .b(b[0]), .out(u_csamul_cska32_and26_0));
  and_gate and_gate_u_csamul_cska32_and27_0(.a(a[27]), .b(b[0]), .out(u_csamul_cska32_and27_0));
  and_gate and_gate_u_csamul_cska32_and28_0(.a(a[28]), .b(b[0]), .out(u_csamul_cska32_and28_0));
  and_gate and_gate_u_csamul_cska32_and29_0(.a(a[29]), .b(b[0]), .out(u_csamul_cska32_and29_0));
  and_gate and_gate_u_csamul_cska32_and30_0(.a(a[30]), .b(b[0]), .out(u_csamul_cska32_and30_0));
  and_gate and_gate_u_csamul_cska32_and31_0(.a(a[31]), .b(b[0]), .out(u_csamul_cska32_and31_0));
  and_gate and_gate_u_csamul_cska32_and0_1(.a(a[0]), .b(b[1]), .out(u_csamul_cska32_and0_1));
  ha ha_u_csamul_cska32_ha0_1_out(.a(u_csamul_cska32_and0_1[0]), .b(u_csamul_cska32_and1_0[0]), .ha_xor0(u_csamul_cska32_ha0_1_xor0), .ha_and0(u_csamul_cska32_ha0_1_and0));
  and_gate and_gate_u_csamul_cska32_and1_1(.a(a[1]), .b(b[1]), .out(u_csamul_cska32_and1_1));
  ha ha_u_csamul_cska32_ha1_1_out(.a(u_csamul_cska32_and1_1[0]), .b(u_csamul_cska32_and2_0[0]), .ha_xor0(u_csamul_cska32_ha1_1_xor0), .ha_and0(u_csamul_cska32_ha1_1_and0));
  and_gate and_gate_u_csamul_cska32_and2_1(.a(a[2]), .b(b[1]), .out(u_csamul_cska32_and2_1));
  ha ha_u_csamul_cska32_ha2_1_out(.a(u_csamul_cska32_and2_1[0]), .b(u_csamul_cska32_and3_0[0]), .ha_xor0(u_csamul_cska32_ha2_1_xor0), .ha_and0(u_csamul_cska32_ha2_1_and0));
  and_gate and_gate_u_csamul_cska32_and3_1(.a(a[3]), .b(b[1]), .out(u_csamul_cska32_and3_1));
  ha ha_u_csamul_cska32_ha3_1_out(.a(u_csamul_cska32_and3_1[0]), .b(u_csamul_cska32_and4_0[0]), .ha_xor0(u_csamul_cska32_ha3_1_xor0), .ha_and0(u_csamul_cska32_ha3_1_and0));
  and_gate and_gate_u_csamul_cska32_and4_1(.a(a[4]), .b(b[1]), .out(u_csamul_cska32_and4_1));
  ha ha_u_csamul_cska32_ha4_1_out(.a(u_csamul_cska32_and4_1[0]), .b(u_csamul_cska32_and5_0[0]), .ha_xor0(u_csamul_cska32_ha4_1_xor0), .ha_and0(u_csamul_cska32_ha4_1_and0));
  and_gate and_gate_u_csamul_cska32_and5_1(.a(a[5]), .b(b[1]), .out(u_csamul_cska32_and5_1));
  ha ha_u_csamul_cska32_ha5_1_out(.a(u_csamul_cska32_and5_1[0]), .b(u_csamul_cska32_and6_0[0]), .ha_xor0(u_csamul_cska32_ha5_1_xor0), .ha_and0(u_csamul_cska32_ha5_1_and0));
  and_gate and_gate_u_csamul_cska32_and6_1(.a(a[6]), .b(b[1]), .out(u_csamul_cska32_and6_1));
  ha ha_u_csamul_cska32_ha6_1_out(.a(u_csamul_cska32_and6_1[0]), .b(u_csamul_cska32_and7_0[0]), .ha_xor0(u_csamul_cska32_ha6_1_xor0), .ha_and0(u_csamul_cska32_ha6_1_and0));
  and_gate and_gate_u_csamul_cska32_and7_1(.a(a[7]), .b(b[1]), .out(u_csamul_cska32_and7_1));
  ha ha_u_csamul_cska32_ha7_1_out(.a(u_csamul_cska32_and7_1[0]), .b(u_csamul_cska32_and8_0[0]), .ha_xor0(u_csamul_cska32_ha7_1_xor0), .ha_and0(u_csamul_cska32_ha7_1_and0));
  and_gate and_gate_u_csamul_cska32_and8_1(.a(a[8]), .b(b[1]), .out(u_csamul_cska32_and8_1));
  ha ha_u_csamul_cska32_ha8_1_out(.a(u_csamul_cska32_and8_1[0]), .b(u_csamul_cska32_and9_0[0]), .ha_xor0(u_csamul_cska32_ha8_1_xor0), .ha_and0(u_csamul_cska32_ha8_1_and0));
  and_gate and_gate_u_csamul_cska32_and9_1(.a(a[9]), .b(b[1]), .out(u_csamul_cska32_and9_1));
  ha ha_u_csamul_cska32_ha9_1_out(.a(u_csamul_cska32_and9_1[0]), .b(u_csamul_cska32_and10_0[0]), .ha_xor0(u_csamul_cska32_ha9_1_xor0), .ha_and0(u_csamul_cska32_ha9_1_and0));
  and_gate and_gate_u_csamul_cska32_and10_1(.a(a[10]), .b(b[1]), .out(u_csamul_cska32_and10_1));
  ha ha_u_csamul_cska32_ha10_1_out(.a(u_csamul_cska32_and10_1[0]), .b(u_csamul_cska32_and11_0[0]), .ha_xor0(u_csamul_cska32_ha10_1_xor0), .ha_and0(u_csamul_cska32_ha10_1_and0));
  and_gate and_gate_u_csamul_cska32_and11_1(.a(a[11]), .b(b[1]), .out(u_csamul_cska32_and11_1));
  ha ha_u_csamul_cska32_ha11_1_out(.a(u_csamul_cska32_and11_1[0]), .b(u_csamul_cska32_and12_0[0]), .ha_xor0(u_csamul_cska32_ha11_1_xor0), .ha_and0(u_csamul_cska32_ha11_1_and0));
  and_gate and_gate_u_csamul_cska32_and12_1(.a(a[12]), .b(b[1]), .out(u_csamul_cska32_and12_1));
  ha ha_u_csamul_cska32_ha12_1_out(.a(u_csamul_cska32_and12_1[0]), .b(u_csamul_cska32_and13_0[0]), .ha_xor0(u_csamul_cska32_ha12_1_xor0), .ha_and0(u_csamul_cska32_ha12_1_and0));
  and_gate and_gate_u_csamul_cska32_and13_1(.a(a[13]), .b(b[1]), .out(u_csamul_cska32_and13_1));
  ha ha_u_csamul_cska32_ha13_1_out(.a(u_csamul_cska32_and13_1[0]), .b(u_csamul_cska32_and14_0[0]), .ha_xor0(u_csamul_cska32_ha13_1_xor0), .ha_and0(u_csamul_cska32_ha13_1_and0));
  and_gate and_gate_u_csamul_cska32_and14_1(.a(a[14]), .b(b[1]), .out(u_csamul_cska32_and14_1));
  ha ha_u_csamul_cska32_ha14_1_out(.a(u_csamul_cska32_and14_1[0]), .b(u_csamul_cska32_and15_0[0]), .ha_xor0(u_csamul_cska32_ha14_1_xor0), .ha_and0(u_csamul_cska32_ha14_1_and0));
  and_gate and_gate_u_csamul_cska32_and15_1(.a(a[15]), .b(b[1]), .out(u_csamul_cska32_and15_1));
  ha ha_u_csamul_cska32_ha15_1_out(.a(u_csamul_cska32_and15_1[0]), .b(u_csamul_cska32_and16_0[0]), .ha_xor0(u_csamul_cska32_ha15_1_xor0), .ha_and0(u_csamul_cska32_ha15_1_and0));
  and_gate and_gate_u_csamul_cska32_and16_1(.a(a[16]), .b(b[1]), .out(u_csamul_cska32_and16_1));
  ha ha_u_csamul_cska32_ha16_1_out(.a(u_csamul_cska32_and16_1[0]), .b(u_csamul_cska32_and17_0[0]), .ha_xor0(u_csamul_cska32_ha16_1_xor0), .ha_and0(u_csamul_cska32_ha16_1_and0));
  and_gate and_gate_u_csamul_cska32_and17_1(.a(a[17]), .b(b[1]), .out(u_csamul_cska32_and17_1));
  ha ha_u_csamul_cska32_ha17_1_out(.a(u_csamul_cska32_and17_1[0]), .b(u_csamul_cska32_and18_0[0]), .ha_xor0(u_csamul_cska32_ha17_1_xor0), .ha_and0(u_csamul_cska32_ha17_1_and0));
  and_gate and_gate_u_csamul_cska32_and18_1(.a(a[18]), .b(b[1]), .out(u_csamul_cska32_and18_1));
  ha ha_u_csamul_cska32_ha18_1_out(.a(u_csamul_cska32_and18_1[0]), .b(u_csamul_cska32_and19_0[0]), .ha_xor0(u_csamul_cska32_ha18_1_xor0), .ha_and0(u_csamul_cska32_ha18_1_and0));
  and_gate and_gate_u_csamul_cska32_and19_1(.a(a[19]), .b(b[1]), .out(u_csamul_cska32_and19_1));
  ha ha_u_csamul_cska32_ha19_1_out(.a(u_csamul_cska32_and19_1[0]), .b(u_csamul_cska32_and20_0[0]), .ha_xor0(u_csamul_cska32_ha19_1_xor0), .ha_and0(u_csamul_cska32_ha19_1_and0));
  and_gate and_gate_u_csamul_cska32_and20_1(.a(a[20]), .b(b[1]), .out(u_csamul_cska32_and20_1));
  ha ha_u_csamul_cska32_ha20_1_out(.a(u_csamul_cska32_and20_1[0]), .b(u_csamul_cska32_and21_0[0]), .ha_xor0(u_csamul_cska32_ha20_1_xor0), .ha_and0(u_csamul_cska32_ha20_1_and0));
  and_gate and_gate_u_csamul_cska32_and21_1(.a(a[21]), .b(b[1]), .out(u_csamul_cska32_and21_1));
  ha ha_u_csamul_cska32_ha21_1_out(.a(u_csamul_cska32_and21_1[0]), .b(u_csamul_cska32_and22_0[0]), .ha_xor0(u_csamul_cska32_ha21_1_xor0), .ha_and0(u_csamul_cska32_ha21_1_and0));
  and_gate and_gate_u_csamul_cska32_and22_1(.a(a[22]), .b(b[1]), .out(u_csamul_cska32_and22_1));
  ha ha_u_csamul_cska32_ha22_1_out(.a(u_csamul_cska32_and22_1[0]), .b(u_csamul_cska32_and23_0[0]), .ha_xor0(u_csamul_cska32_ha22_1_xor0), .ha_and0(u_csamul_cska32_ha22_1_and0));
  and_gate and_gate_u_csamul_cska32_and23_1(.a(a[23]), .b(b[1]), .out(u_csamul_cska32_and23_1));
  ha ha_u_csamul_cska32_ha23_1_out(.a(u_csamul_cska32_and23_1[0]), .b(u_csamul_cska32_and24_0[0]), .ha_xor0(u_csamul_cska32_ha23_1_xor0), .ha_and0(u_csamul_cska32_ha23_1_and0));
  and_gate and_gate_u_csamul_cska32_and24_1(.a(a[24]), .b(b[1]), .out(u_csamul_cska32_and24_1));
  ha ha_u_csamul_cska32_ha24_1_out(.a(u_csamul_cska32_and24_1[0]), .b(u_csamul_cska32_and25_0[0]), .ha_xor0(u_csamul_cska32_ha24_1_xor0), .ha_and0(u_csamul_cska32_ha24_1_and0));
  and_gate and_gate_u_csamul_cska32_and25_1(.a(a[25]), .b(b[1]), .out(u_csamul_cska32_and25_1));
  ha ha_u_csamul_cska32_ha25_1_out(.a(u_csamul_cska32_and25_1[0]), .b(u_csamul_cska32_and26_0[0]), .ha_xor0(u_csamul_cska32_ha25_1_xor0), .ha_and0(u_csamul_cska32_ha25_1_and0));
  and_gate and_gate_u_csamul_cska32_and26_1(.a(a[26]), .b(b[1]), .out(u_csamul_cska32_and26_1));
  ha ha_u_csamul_cska32_ha26_1_out(.a(u_csamul_cska32_and26_1[0]), .b(u_csamul_cska32_and27_0[0]), .ha_xor0(u_csamul_cska32_ha26_1_xor0), .ha_and0(u_csamul_cska32_ha26_1_and0));
  and_gate and_gate_u_csamul_cska32_and27_1(.a(a[27]), .b(b[1]), .out(u_csamul_cska32_and27_1));
  ha ha_u_csamul_cska32_ha27_1_out(.a(u_csamul_cska32_and27_1[0]), .b(u_csamul_cska32_and28_0[0]), .ha_xor0(u_csamul_cska32_ha27_1_xor0), .ha_and0(u_csamul_cska32_ha27_1_and0));
  and_gate and_gate_u_csamul_cska32_and28_1(.a(a[28]), .b(b[1]), .out(u_csamul_cska32_and28_1));
  ha ha_u_csamul_cska32_ha28_1_out(.a(u_csamul_cska32_and28_1[0]), .b(u_csamul_cska32_and29_0[0]), .ha_xor0(u_csamul_cska32_ha28_1_xor0), .ha_and0(u_csamul_cska32_ha28_1_and0));
  and_gate and_gate_u_csamul_cska32_and29_1(.a(a[29]), .b(b[1]), .out(u_csamul_cska32_and29_1));
  ha ha_u_csamul_cska32_ha29_1_out(.a(u_csamul_cska32_and29_1[0]), .b(u_csamul_cska32_and30_0[0]), .ha_xor0(u_csamul_cska32_ha29_1_xor0), .ha_and0(u_csamul_cska32_ha29_1_and0));
  and_gate and_gate_u_csamul_cska32_and30_1(.a(a[30]), .b(b[1]), .out(u_csamul_cska32_and30_1));
  ha ha_u_csamul_cska32_ha30_1_out(.a(u_csamul_cska32_and30_1[0]), .b(u_csamul_cska32_and31_0[0]), .ha_xor0(u_csamul_cska32_ha30_1_xor0), .ha_and0(u_csamul_cska32_ha30_1_and0));
  and_gate and_gate_u_csamul_cska32_and31_1(.a(a[31]), .b(b[1]), .out(u_csamul_cska32_and31_1));
  and_gate and_gate_u_csamul_cska32_and0_2(.a(a[0]), .b(b[2]), .out(u_csamul_cska32_and0_2));
  fa fa_u_csamul_cska32_fa0_2_out(.a(u_csamul_cska32_and0_2[0]), .b(u_csamul_cska32_ha1_1_xor0[0]), .cin(u_csamul_cska32_ha0_1_and0[0]), .fa_xor1(u_csamul_cska32_fa0_2_xor1), .fa_or0(u_csamul_cska32_fa0_2_or0));
  and_gate and_gate_u_csamul_cska32_and1_2(.a(a[1]), .b(b[2]), .out(u_csamul_cska32_and1_2));
  fa fa_u_csamul_cska32_fa1_2_out(.a(u_csamul_cska32_and1_2[0]), .b(u_csamul_cska32_ha2_1_xor0[0]), .cin(u_csamul_cska32_ha1_1_and0[0]), .fa_xor1(u_csamul_cska32_fa1_2_xor1), .fa_or0(u_csamul_cska32_fa1_2_or0));
  and_gate and_gate_u_csamul_cska32_and2_2(.a(a[2]), .b(b[2]), .out(u_csamul_cska32_and2_2));
  fa fa_u_csamul_cska32_fa2_2_out(.a(u_csamul_cska32_and2_2[0]), .b(u_csamul_cska32_ha3_1_xor0[0]), .cin(u_csamul_cska32_ha2_1_and0[0]), .fa_xor1(u_csamul_cska32_fa2_2_xor1), .fa_or0(u_csamul_cska32_fa2_2_or0));
  and_gate and_gate_u_csamul_cska32_and3_2(.a(a[3]), .b(b[2]), .out(u_csamul_cska32_and3_2));
  fa fa_u_csamul_cska32_fa3_2_out(.a(u_csamul_cska32_and3_2[0]), .b(u_csamul_cska32_ha4_1_xor0[0]), .cin(u_csamul_cska32_ha3_1_and0[0]), .fa_xor1(u_csamul_cska32_fa3_2_xor1), .fa_or0(u_csamul_cska32_fa3_2_or0));
  and_gate and_gate_u_csamul_cska32_and4_2(.a(a[4]), .b(b[2]), .out(u_csamul_cska32_and4_2));
  fa fa_u_csamul_cska32_fa4_2_out(.a(u_csamul_cska32_and4_2[0]), .b(u_csamul_cska32_ha5_1_xor0[0]), .cin(u_csamul_cska32_ha4_1_and0[0]), .fa_xor1(u_csamul_cska32_fa4_2_xor1), .fa_or0(u_csamul_cska32_fa4_2_or0));
  and_gate and_gate_u_csamul_cska32_and5_2(.a(a[5]), .b(b[2]), .out(u_csamul_cska32_and5_2));
  fa fa_u_csamul_cska32_fa5_2_out(.a(u_csamul_cska32_and5_2[0]), .b(u_csamul_cska32_ha6_1_xor0[0]), .cin(u_csamul_cska32_ha5_1_and0[0]), .fa_xor1(u_csamul_cska32_fa5_2_xor1), .fa_or0(u_csamul_cska32_fa5_2_or0));
  and_gate and_gate_u_csamul_cska32_and6_2(.a(a[6]), .b(b[2]), .out(u_csamul_cska32_and6_2));
  fa fa_u_csamul_cska32_fa6_2_out(.a(u_csamul_cska32_and6_2[0]), .b(u_csamul_cska32_ha7_1_xor0[0]), .cin(u_csamul_cska32_ha6_1_and0[0]), .fa_xor1(u_csamul_cska32_fa6_2_xor1), .fa_or0(u_csamul_cska32_fa6_2_or0));
  and_gate and_gate_u_csamul_cska32_and7_2(.a(a[7]), .b(b[2]), .out(u_csamul_cska32_and7_2));
  fa fa_u_csamul_cska32_fa7_2_out(.a(u_csamul_cska32_and7_2[0]), .b(u_csamul_cska32_ha8_1_xor0[0]), .cin(u_csamul_cska32_ha7_1_and0[0]), .fa_xor1(u_csamul_cska32_fa7_2_xor1), .fa_or0(u_csamul_cska32_fa7_2_or0));
  and_gate and_gate_u_csamul_cska32_and8_2(.a(a[8]), .b(b[2]), .out(u_csamul_cska32_and8_2));
  fa fa_u_csamul_cska32_fa8_2_out(.a(u_csamul_cska32_and8_2[0]), .b(u_csamul_cska32_ha9_1_xor0[0]), .cin(u_csamul_cska32_ha8_1_and0[0]), .fa_xor1(u_csamul_cska32_fa8_2_xor1), .fa_or0(u_csamul_cska32_fa8_2_or0));
  and_gate and_gate_u_csamul_cska32_and9_2(.a(a[9]), .b(b[2]), .out(u_csamul_cska32_and9_2));
  fa fa_u_csamul_cska32_fa9_2_out(.a(u_csamul_cska32_and9_2[0]), .b(u_csamul_cska32_ha10_1_xor0[0]), .cin(u_csamul_cska32_ha9_1_and0[0]), .fa_xor1(u_csamul_cska32_fa9_2_xor1), .fa_or0(u_csamul_cska32_fa9_2_or0));
  and_gate and_gate_u_csamul_cska32_and10_2(.a(a[10]), .b(b[2]), .out(u_csamul_cska32_and10_2));
  fa fa_u_csamul_cska32_fa10_2_out(.a(u_csamul_cska32_and10_2[0]), .b(u_csamul_cska32_ha11_1_xor0[0]), .cin(u_csamul_cska32_ha10_1_and0[0]), .fa_xor1(u_csamul_cska32_fa10_2_xor1), .fa_or0(u_csamul_cska32_fa10_2_or0));
  and_gate and_gate_u_csamul_cska32_and11_2(.a(a[11]), .b(b[2]), .out(u_csamul_cska32_and11_2));
  fa fa_u_csamul_cska32_fa11_2_out(.a(u_csamul_cska32_and11_2[0]), .b(u_csamul_cska32_ha12_1_xor0[0]), .cin(u_csamul_cska32_ha11_1_and0[0]), .fa_xor1(u_csamul_cska32_fa11_2_xor1), .fa_or0(u_csamul_cska32_fa11_2_or0));
  and_gate and_gate_u_csamul_cska32_and12_2(.a(a[12]), .b(b[2]), .out(u_csamul_cska32_and12_2));
  fa fa_u_csamul_cska32_fa12_2_out(.a(u_csamul_cska32_and12_2[0]), .b(u_csamul_cska32_ha13_1_xor0[0]), .cin(u_csamul_cska32_ha12_1_and0[0]), .fa_xor1(u_csamul_cska32_fa12_2_xor1), .fa_or0(u_csamul_cska32_fa12_2_or0));
  and_gate and_gate_u_csamul_cska32_and13_2(.a(a[13]), .b(b[2]), .out(u_csamul_cska32_and13_2));
  fa fa_u_csamul_cska32_fa13_2_out(.a(u_csamul_cska32_and13_2[0]), .b(u_csamul_cska32_ha14_1_xor0[0]), .cin(u_csamul_cska32_ha13_1_and0[0]), .fa_xor1(u_csamul_cska32_fa13_2_xor1), .fa_or0(u_csamul_cska32_fa13_2_or0));
  and_gate and_gate_u_csamul_cska32_and14_2(.a(a[14]), .b(b[2]), .out(u_csamul_cska32_and14_2));
  fa fa_u_csamul_cska32_fa14_2_out(.a(u_csamul_cska32_and14_2[0]), .b(u_csamul_cska32_ha15_1_xor0[0]), .cin(u_csamul_cska32_ha14_1_and0[0]), .fa_xor1(u_csamul_cska32_fa14_2_xor1), .fa_or0(u_csamul_cska32_fa14_2_or0));
  and_gate and_gate_u_csamul_cska32_and15_2(.a(a[15]), .b(b[2]), .out(u_csamul_cska32_and15_2));
  fa fa_u_csamul_cska32_fa15_2_out(.a(u_csamul_cska32_and15_2[0]), .b(u_csamul_cska32_ha16_1_xor0[0]), .cin(u_csamul_cska32_ha15_1_and0[0]), .fa_xor1(u_csamul_cska32_fa15_2_xor1), .fa_or0(u_csamul_cska32_fa15_2_or0));
  and_gate and_gate_u_csamul_cska32_and16_2(.a(a[16]), .b(b[2]), .out(u_csamul_cska32_and16_2));
  fa fa_u_csamul_cska32_fa16_2_out(.a(u_csamul_cska32_and16_2[0]), .b(u_csamul_cska32_ha17_1_xor0[0]), .cin(u_csamul_cska32_ha16_1_and0[0]), .fa_xor1(u_csamul_cska32_fa16_2_xor1), .fa_or0(u_csamul_cska32_fa16_2_or0));
  and_gate and_gate_u_csamul_cska32_and17_2(.a(a[17]), .b(b[2]), .out(u_csamul_cska32_and17_2));
  fa fa_u_csamul_cska32_fa17_2_out(.a(u_csamul_cska32_and17_2[0]), .b(u_csamul_cska32_ha18_1_xor0[0]), .cin(u_csamul_cska32_ha17_1_and0[0]), .fa_xor1(u_csamul_cska32_fa17_2_xor1), .fa_or0(u_csamul_cska32_fa17_2_or0));
  and_gate and_gate_u_csamul_cska32_and18_2(.a(a[18]), .b(b[2]), .out(u_csamul_cska32_and18_2));
  fa fa_u_csamul_cska32_fa18_2_out(.a(u_csamul_cska32_and18_2[0]), .b(u_csamul_cska32_ha19_1_xor0[0]), .cin(u_csamul_cska32_ha18_1_and0[0]), .fa_xor1(u_csamul_cska32_fa18_2_xor1), .fa_or0(u_csamul_cska32_fa18_2_or0));
  and_gate and_gate_u_csamul_cska32_and19_2(.a(a[19]), .b(b[2]), .out(u_csamul_cska32_and19_2));
  fa fa_u_csamul_cska32_fa19_2_out(.a(u_csamul_cska32_and19_2[0]), .b(u_csamul_cska32_ha20_1_xor0[0]), .cin(u_csamul_cska32_ha19_1_and0[0]), .fa_xor1(u_csamul_cska32_fa19_2_xor1), .fa_or0(u_csamul_cska32_fa19_2_or0));
  and_gate and_gate_u_csamul_cska32_and20_2(.a(a[20]), .b(b[2]), .out(u_csamul_cska32_and20_2));
  fa fa_u_csamul_cska32_fa20_2_out(.a(u_csamul_cska32_and20_2[0]), .b(u_csamul_cska32_ha21_1_xor0[0]), .cin(u_csamul_cska32_ha20_1_and0[0]), .fa_xor1(u_csamul_cska32_fa20_2_xor1), .fa_or0(u_csamul_cska32_fa20_2_or0));
  and_gate and_gate_u_csamul_cska32_and21_2(.a(a[21]), .b(b[2]), .out(u_csamul_cska32_and21_2));
  fa fa_u_csamul_cska32_fa21_2_out(.a(u_csamul_cska32_and21_2[0]), .b(u_csamul_cska32_ha22_1_xor0[0]), .cin(u_csamul_cska32_ha21_1_and0[0]), .fa_xor1(u_csamul_cska32_fa21_2_xor1), .fa_or0(u_csamul_cska32_fa21_2_or0));
  and_gate and_gate_u_csamul_cska32_and22_2(.a(a[22]), .b(b[2]), .out(u_csamul_cska32_and22_2));
  fa fa_u_csamul_cska32_fa22_2_out(.a(u_csamul_cska32_and22_2[0]), .b(u_csamul_cska32_ha23_1_xor0[0]), .cin(u_csamul_cska32_ha22_1_and0[0]), .fa_xor1(u_csamul_cska32_fa22_2_xor1), .fa_or0(u_csamul_cska32_fa22_2_or0));
  and_gate and_gate_u_csamul_cska32_and23_2(.a(a[23]), .b(b[2]), .out(u_csamul_cska32_and23_2));
  fa fa_u_csamul_cska32_fa23_2_out(.a(u_csamul_cska32_and23_2[0]), .b(u_csamul_cska32_ha24_1_xor0[0]), .cin(u_csamul_cska32_ha23_1_and0[0]), .fa_xor1(u_csamul_cska32_fa23_2_xor1), .fa_or0(u_csamul_cska32_fa23_2_or0));
  and_gate and_gate_u_csamul_cska32_and24_2(.a(a[24]), .b(b[2]), .out(u_csamul_cska32_and24_2));
  fa fa_u_csamul_cska32_fa24_2_out(.a(u_csamul_cska32_and24_2[0]), .b(u_csamul_cska32_ha25_1_xor0[0]), .cin(u_csamul_cska32_ha24_1_and0[0]), .fa_xor1(u_csamul_cska32_fa24_2_xor1), .fa_or0(u_csamul_cska32_fa24_2_or0));
  and_gate and_gate_u_csamul_cska32_and25_2(.a(a[25]), .b(b[2]), .out(u_csamul_cska32_and25_2));
  fa fa_u_csamul_cska32_fa25_2_out(.a(u_csamul_cska32_and25_2[0]), .b(u_csamul_cska32_ha26_1_xor0[0]), .cin(u_csamul_cska32_ha25_1_and0[0]), .fa_xor1(u_csamul_cska32_fa25_2_xor1), .fa_or0(u_csamul_cska32_fa25_2_or0));
  and_gate and_gate_u_csamul_cska32_and26_2(.a(a[26]), .b(b[2]), .out(u_csamul_cska32_and26_2));
  fa fa_u_csamul_cska32_fa26_2_out(.a(u_csamul_cska32_and26_2[0]), .b(u_csamul_cska32_ha27_1_xor0[0]), .cin(u_csamul_cska32_ha26_1_and0[0]), .fa_xor1(u_csamul_cska32_fa26_2_xor1), .fa_or0(u_csamul_cska32_fa26_2_or0));
  and_gate and_gate_u_csamul_cska32_and27_2(.a(a[27]), .b(b[2]), .out(u_csamul_cska32_and27_2));
  fa fa_u_csamul_cska32_fa27_2_out(.a(u_csamul_cska32_and27_2[0]), .b(u_csamul_cska32_ha28_1_xor0[0]), .cin(u_csamul_cska32_ha27_1_and0[0]), .fa_xor1(u_csamul_cska32_fa27_2_xor1), .fa_or0(u_csamul_cska32_fa27_2_or0));
  and_gate and_gate_u_csamul_cska32_and28_2(.a(a[28]), .b(b[2]), .out(u_csamul_cska32_and28_2));
  fa fa_u_csamul_cska32_fa28_2_out(.a(u_csamul_cska32_and28_2[0]), .b(u_csamul_cska32_ha29_1_xor0[0]), .cin(u_csamul_cska32_ha28_1_and0[0]), .fa_xor1(u_csamul_cska32_fa28_2_xor1), .fa_or0(u_csamul_cska32_fa28_2_or0));
  and_gate and_gate_u_csamul_cska32_and29_2(.a(a[29]), .b(b[2]), .out(u_csamul_cska32_and29_2));
  fa fa_u_csamul_cska32_fa29_2_out(.a(u_csamul_cska32_and29_2[0]), .b(u_csamul_cska32_ha30_1_xor0[0]), .cin(u_csamul_cska32_ha29_1_and0[0]), .fa_xor1(u_csamul_cska32_fa29_2_xor1), .fa_or0(u_csamul_cska32_fa29_2_or0));
  and_gate and_gate_u_csamul_cska32_and30_2(.a(a[30]), .b(b[2]), .out(u_csamul_cska32_and30_2));
  fa fa_u_csamul_cska32_fa30_2_out(.a(u_csamul_cska32_and30_2[0]), .b(u_csamul_cska32_and31_1[0]), .cin(u_csamul_cska32_ha30_1_and0[0]), .fa_xor1(u_csamul_cska32_fa30_2_xor1), .fa_or0(u_csamul_cska32_fa30_2_or0));
  and_gate and_gate_u_csamul_cska32_and31_2(.a(a[31]), .b(b[2]), .out(u_csamul_cska32_and31_2));
  and_gate and_gate_u_csamul_cska32_and0_3(.a(a[0]), .b(b[3]), .out(u_csamul_cska32_and0_3));
  fa fa_u_csamul_cska32_fa0_3_out(.a(u_csamul_cska32_and0_3[0]), .b(u_csamul_cska32_fa1_2_xor1[0]), .cin(u_csamul_cska32_fa0_2_or0[0]), .fa_xor1(u_csamul_cska32_fa0_3_xor1), .fa_or0(u_csamul_cska32_fa0_3_or0));
  and_gate and_gate_u_csamul_cska32_and1_3(.a(a[1]), .b(b[3]), .out(u_csamul_cska32_and1_3));
  fa fa_u_csamul_cska32_fa1_3_out(.a(u_csamul_cska32_and1_3[0]), .b(u_csamul_cska32_fa2_2_xor1[0]), .cin(u_csamul_cska32_fa1_2_or0[0]), .fa_xor1(u_csamul_cska32_fa1_3_xor1), .fa_or0(u_csamul_cska32_fa1_3_or0));
  and_gate and_gate_u_csamul_cska32_and2_3(.a(a[2]), .b(b[3]), .out(u_csamul_cska32_and2_3));
  fa fa_u_csamul_cska32_fa2_3_out(.a(u_csamul_cska32_and2_3[0]), .b(u_csamul_cska32_fa3_2_xor1[0]), .cin(u_csamul_cska32_fa2_2_or0[0]), .fa_xor1(u_csamul_cska32_fa2_3_xor1), .fa_or0(u_csamul_cska32_fa2_3_or0));
  and_gate and_gate_u_csamul_cska32_and3_3(.a(a[3]), .b(b[3]), .out(u_csamul_cska32_and3_3));
  fa fa_u_csamul_cska32_fa3_3_out(.a(u_csamul_cska32_and3_3[0]), .b(u_csamul_cska32_fa4_2_xor1[0]), .cin(u_csamul_cska32_fa3_2_or0[0]), .fa_xor1(u_csamul_cska32_fa3_3_xor1), .fa_or0(u_csamul_cska32_fa3_3_or0));
  and_gate and_gate_u_csamul_cska32_and4_3(.a(a[4]), .b(b[3]), .out(u_csamul_cska32_and4_3));
  fa fa_u_csamul_cska32_fa4_3_out(.a(u_csamul_cska32_and4_3[0]), .b(u_csamul_cska32_fa5_2_xor1[0]), .cin(u_csamul_cska32_fa4_2_or0[0]), .fa_xor1(u_csamul_cska32_fa4_3_xor1), .fa_or0(u_csamul_cska32_fa4_3_or0));
  and_gate and_gate_u_csamul_cska32_and5_3(.a(a[5]), .b(b[3]), .out(u_csamul_cska32_and5_3));
  fa fa_u_csamul_cska32_fa5_3_out(.a(u_csamul_cska32_and5_3[0]), .b(u_csamul_cska32_fa6_2_xor1[0]), .cin(u_csamul_cska32_fa5_2_or0[0]), .fa_xor1(u_csamul_cska32_fa5_3_xor1), .fa_or0(u_csamul_cska32_fa5_3_or0));
  and_gate and_gate_u_csamul_cska32_and6_3(.a(a[6]), .b(b[3]), .out(u_csamul_cska32_and6_3));
  fa fa_u_csamul_cska32_fa6_3_out(.a(u_csamul_cska32_and6_3[0]), .b(u_csamul_cska32_fa7_2_xor1[0]), .cin(u_csamul_cska32_fa6_2_or0[0]), .fa_xor1(u_csamul_cska32_fa6_3_xor1), .fa_or0(u_csamul_cska32_fa6_3_or0));
  and_gate and_gate_u_csamul_cska32_and7_3(.a(a[7]), .b(b[3]), .out(u_csamul_cska32_and7_3));
  fa fa_u_csamul_cska32_fa7_3_out(.a(u_csamul_cska32_and7_3[0]), .b(u_csamul_cska32_fa8_2_xor1[0]), .cin(u_csamul_cska32_fa7_2_or0[0]), .fa_xor1(u_csamul_cska32_fa7_3_xor1), .fa_or0(u_csamul_cska32_fa7_3_or0));
  and_gate and_gate_u_csamul_cska32_and8_3(.a(a[8]), .b(b[3]), .out(u_csamul_cska32_and8_3));
  fa fa_u_csamul_cska32_fa8_3_out(.a(u_csamul_cska32_and8_3[0]), .b(u_csamul_cska32_fa9_2_xor1[0]), .cin(u_csamul_cska32_fa8_2_or0[0]), .fa_xor1(u_csamul_cska32_fa8_3_xor1), .fa_or0(u_csamul_cska32_fa8_3_or0));
  and_gate and_gate_u_csamul_cska32_and9_3(.a(a[9]), .b(b[3]), .out(u_csamul_cska32_and9_3));
  fa fa_u_csamul_cska32_fa9_3_out(.a(u_csamul_cska32_and9_3[0]), .b(u_csamul_cska32_fa10_2_xor1[0]), .cin(u_csamul_cska32_fa9_2_or0[0]), .fa_xor1(u_csamul_cska32_fa9_3_xor1), .fa_or0(u_csamul_cska32_fa9_3_or0));
  and_gate and_gate_u_csamul_cska32_and10_3(.a(a[10]), .b(b[3]), .out(u_csamul_cska32_and10_3));
  fa fa_u_csamul_cska32_fa10_3_out(.a(u_csamul_cska32_and10_3[0]), .b(u_csamul_cska32_fa11_2_xor1[0]), .cin(u_csamul_cska32_fa10_2_or0[0]), .fa_xor1(u_csamul_cska32_fa10_3_xor1), .fa_or0(u_csamul_cska32_fa10_3_or0));
  and_gate and_gate_u_csamul_cska32_and11_3(.a(a[11]), .b(b[3]), .out(u_csamul_cska32_and11_3));
  fa fa_u_csamul_cska32_fa11_3_out(.a(u_csamul_cska32_and11_3[0]), .b(u_csamul_cska32_fa12_2_xor1[0]), .cin(u_csamul_cska32_fa11_2_or0[0]), .fa_xor1(u_csamul_cska32_fa11_3_xor1), .fa_or0(u_csamul_cska32_fa11_3_or0));
  and_gate and_gate_u_csamul_cska32_and12_3(.a(a[12]), .b(b[3]), .out(u_csamul_cska32_and12_3));
  fa fa_u_csamul_cska32_fa12_3_out(.a(u_csamul_cska32_and12_3[0]), .b(u_csamul_cska32_fa13_2_xor1[0]), .cin(u_csamul_cska32_fa12_2_or0[0]), .fa_xor1(u_csamul_cska32_fa12_3_xor1), .fa_or0(u_csamul_cska32_fa12_3_or0));
  and_gate and_gate_u_csamul_cska32_and13_3(.a(a[13]), .b(b[3]), .out(u_csamul_cska32_and13_3));
  fa fa_u_csamul_cska32_fa13_3_out(.a(u_csamul_cska32_and13_3[0]), .b(u_csamul_cska32_fa14_2_xor1[0]), .cin(u_csamul_cska32_fa13_2_or0[0]), .fa_xor1(u_csamul_cska32_fa13_3_xor1), .fa_or0(u_csamul_cska32_fa13_3_or0));
  and_gate and_gate_u_csamul_cska32_and14_3(.a(a[14]), .b(b[3]), .out(u_csamul_cska32_and14_3));
  fa fa_u_csamul_cska32_fa14_3_out(.a(u_csamul_cska32_and14_3[0]), .b(u_csamul_cska32_fa15_2_xor1[0]), .cin(u_csamul_cska32_fa14_2_or0[0]), .fa_xor1(u_csamul_cska32_fa14_3_xor1), .fa_or0(u_csamul_cska32_fa14_3_or0));
  and_gate and_gate_u_csamul_cska32_and15_3(.a(a[15]), .b(b[3]), .out(u_csamul_cska32_and15_3));
  fa fa_u_csamul_cska32_fa15_3_out(.a(u_csamul_cska32_and15_3[0]), .b(u_csamul_cska32_fa16_2_xor1[0]), .cin(u_csamul_cska32_fa15_2_or0[0]), .fa_xor1(u_csamul_cska32_fa15_3_xor1), .fa_or0(u_csamul_cska32_fa15_3_or0));
  and_gate and_gate_u_csamul_cska32_and16_3(.a(a[16]), .b(b[3]), .out(u_csamul_cska32_and16_3));
  fa fa_u_csamul_cska32_fa16_3_out(.a(u_csamul_cska32_and16_3[0]), .b(u_csamul_cska32_fa17_2_xor1[0]), .cin(u_csamul_cska32_fa16_2_or0[0]), .fa_xor1(u_csamul_cska32_fa16_3_xor1), .fa_or0(u_csamul_cska32_fa16_3_or0));
  and_gate and_gate_u_csamul_cska32_and17_3(.a(a[17]), .b(b[3]), .out(u_csamul_cska32_and17_3));
  fa fa_u_csamul_cska32_fa17_3_out(.a(u_csamul_cska32_and17_3[0]), .b(u_csamul_cska32_fa18_2_xor1[0]), .cin(u_csamul_cska32_fa17_2_or0[0]), .fa_xor1(u_csamul_cska32_fa17_3_xor1), .fa_or0(u_csamul_cska32_fa17_3_or0));
  and_gate and_gate_u_csamul_cska32_and18_3(.a(a[18]), .b(b[3]), .out(u_csamul_cska32_and18_3));
  fa fa_u_csamul_cska32_fa18_3_out(.a(u_csamul_cska32_and18_3[0]), .b(u_csamul_cska32_fa19_2_xor1[0]), .cin(u_csamul_cska32_fa18_2_or0[0]), .fa_xor1(u_csamul_cska32_fa18_3_xor1), .fa_or0(u_csamul_cska32_fa18_3_or0));
  and_gate and_gate_u_csamul_cska32_and19_3(.a(a[19]), .b(b[3]), .out(u_csamul_cska32_and19_3));
  fa fa_u_csamul_cska32_fa19_3_out(.a(u_csamul_cska32_and19_3[0]), .b(u_csamul_cska32_fa20_2_xor1[0]), .cin(u_csamul_cska32_fa19_2_or0[0]), .fa_xor1(u_csamul_cska32_fa19_3_xor1), .fa_or0(u_csamul_cska32_fa19_3_or0));
  and_gate and_gate_u_csamul_cska32_and20_3(.a(a[20]), .b(b[3]), .out(u_csamul_cska32_and20_3));
  fa fa_u_csamul_cska32_fa20_3_out(.a(u_csamul_cska32_and20_3[0]), .b(u_csamul_cska32_fa21_2_xor1[0]), .cin(u_csamul_cska32_fa20_2_or0[0]), .fa_xor1(u_csamul_cska32_fa20_3_xor1), .fa_or0(u_csamul_cska32_fa20_3_or0));
  and_gate and_gate_u_csamul_cska32_and21_3(.a(a[21]), .b(b[3]), .out(u_csamul_cska32_and21_3));
  fa fa_u_csamul_cska32_fa21_3_out(.a(u_csamul_cska32_and21_3[0]), .b(u_csamul_cska32_fa22_2_xor1[0]), .cin(u_csamul_cska32_fa21_2_or0[0]), .fa_xor1(u_csamul_cska32_fa21_3_xor1), .fa_or0(u_csamul_cska32_fa21_3_or0));
  and_gate and_gate_u_csamul_cska32_and22_3(.a(a[22]), .b(b[3]), .out(u_csamul_cska32_and22_3));
  fa fa_u_csamul_cska32_fa22_3_out(.a(u_csamul_cska32_and22_3[0]), .b(u_csamul_cska32_fa23_2_xor1[0]), .cin(u_csamul_cska32_fa22_2_or0[0]), .fa_xor1(u_csamul_cska32_fa22_3_xor1), .fa_or0(u_csamul_cska32_fa22_3_or0));
  and_gate and_gate_u_csamul_cska32_and23_3(.a(a[23]), .b(b[3]), .out(u_csamul_cska32_and23_3));
  fa fa_u_csamul_cska32_fa23_3_out(.a(u_csamul_cska32_and23_3[0]), .b(u_csamul_cska32_fa24_2_xor1[0]), .cin(u_csamul_cska32_fa23_2_or0[0]), .fa_xor1(u_csamul_cska32_fa23_3_xor1), .fa_or0(u_csamul_cska32_fa23_3_or0));
  and_gate and_gate_u_csamul_cska32_and24_3(.a(a[24]), .b(b[3]), .out(u_csamul_cska32_and24_3));
  fa fa_u_csamul_cska32_fa24_3_out(.a(u_csamul_cska32_and24_3[0]), .b(u_csamul_cska32_fa25_2_xor1[0]), .cin(u_csamul_cska32_fa24_2_or0[0]), .fa_xor1(u_csamul_cska32_fa24_3_xor1), .fa_or0(u_csamul_cska32_fa24_3_or0));
  and_gate and_gate_u_csamul_cska32_and25_3(.a(a[25]), .b(b[3]), .out(u_csamul_cska32_and25_3));
  fa fa_u_csamul_cska32_fa25_3_out(.a(u_csamul_cska32_and25_3[0]), .b(u_csamul_cska32_fa26_2_xor1[0]), .cin(u_csamul_cska32_fa25_2_or0[0]), .fa_xor1(u_csamul_cska32_fa25_3_xor1), .fa_or0(u_csamul_cska32_fa25_3_or0));
  and_gate and_gate_u_csamul_cska32_and26_3(.a(a[26]), .b(b[3]), .out(u_csamul_cska32_and26_3));
  fa fa_u_csamul_cska32_fa26_3_out(.a(u_csamul_cska32_and26_3[0]), .b(u_csamul_cska32_fa27_2_xor1[0]), .cin(u_csamul_cska32_fa26_2_or0[0]), .fa_xor1(u_csamul_cska32_fa26_3_xor1), .fa_or0(u_csamul_cska32_fa26_3_or0));
  and_gate and_gate_u_csamul_cska32_and27_3(.a(a[27]), .b(b[3]), .out(u_csamul_cska32_and27_3));
  fa fa_u_csamul_cska32_fa27_3_out(.a(u_csamul_cska32_and27_3[0]), .b(u_csamul_cska32_fa28_2_xor1[0]), .cin(u_csamul_cska32_fa27_2_or0[0]), .fa_xor1(u_csamul_cska32_fa27_3_xor1), .fa_or0(u_csamul_cska32_fa27_3_or0));
  and_gate and_gate_u_csamul_cska32_and28_3(.a(a[28]), .b(b[3]), .out(u_csamul_cska32_and28_3));
  fa fa_u_csamul_cska32_fa28_3_out(.a(u_csamul_cska32_and28_3[0]), .b(u_csamul_cska32_fa29_2_xor1[0]), .cin(u_csamul_cska32_fa28_2_or0[0]), .fa_xor1(u_csamul_cska32_fa28_3_xor1), .fa_or0(u_csamul_cska32_fa28_3_or0));
  and_gate and_gate_u_csamul_cska32_and29_3(.a(a[29]), .b(b[3]), .out(u_csamul_cska32_and29_3));
  fa fa_u_csamul_cska32_fa29_3_out(.a(u_csamul_cska32_and29_3[0]), .b(u_csamul_cska32_fa30_2_xor1[0]), .cin(u_csamul_cska32_fa29_2_or0[0]), .fa_xor1(u_csamul_cska32_fa29_3_xor1), .fa_or0(u_csamul_cska32_fa29_3_or0));
  and_gate and_gate_u_csamul_cska32_and30_3(.a(a[30]), .b(b[3]), .out(u_csamul_cska32_and30_3));
  fa fa_u_csamul_cska32_fa30_3_out(.a(u_csamul_cska32_and30_3[0]), .b(u_csamul_cska32_and31_2[0]), .cin(u_csamul_cska32_fa30_2_or0[0]), .fa_xor1(u_csamul_cska32_fa30_3_xor1), .fa_or0(u_csamul_cska32_fa30_3_or0));
  and_gate and_gate_u_csamul_cska32_and31_3(.a(a[31]), .b(b[3]), .out(u_csamul_cska32_and31_3));
  and_gate and_gate_u_csamul_cska32_and0_4(.a(a[0]), .b(b[4]), .out(u_csamul_cska32_and0_4));
  fa fa_u_csamul_cska32_fa0_4_out(.a(u_csamul_cska32_and0_4[0]), .b(u_csamul_cska32_fa1_3_xor1[0]), .cin(u_csamul_cska32_fa0_3_or0[0]), .fa_xor1(u_csamul_cska32_fa0_4_xor1), .fa_or0(u_csamul_cska32_fa0_4_or0));
  and_gate and_gate_u_csamul_cska32_and1_4(.a(a[1]), .b(b[4]), .out(u_csamul_cska32_and1_4));
  fa fa_u_csamul_cska32_fa1_4_out(.a(u_csamul_cska32_and1_4[0]), .b(u_csamul_cska32_fa2_3_xor1[0]), .cin(u_csamul_cska32_fa1_3_or0[0]), .fa_xor1(u_csamul_cska32_fa1_4_xor1), .fa_or0(u_csamul_cska32_fa1_4_or0));
  and_gate and_gate_u_csamul_cska32_and2_4(.a(a[2]), .b(b[4]), .out(u_csamul_cska32_and2_4));
  fa fa_u_csamul_cska32_fa2_4_out(.a(u_csamul_cska32_and2_4[0]), .b(u_csamul_cska32_fa3_3_xor1[0]), .cin(u_csamul_cska32_fa2_3_or0[0]), .fa_xor1(u_csamul_cska32_fa2_4_xor1), .fa_or0(u_csamul_cska32_fa2_4_or0));
  and_gate and_gate_u_csamul_cska32_and3_4(.a(a[3]), .b(b[4]), .out(u_csamul_cska32_and3_4));
  fa fa_u_csamul_cska32_fa3_4_out(.a(u_csamul_cska32_and3_4[0]), .b(u_csamul_cska32_fa4_3_xor1[0]), .cin(u_csamul_cska32_fa3_3_or0[0]), .fa_xor1(u_csamul_cska32_fa3_4_xor1), .fa_or0(u_csamul_cska32_fa3_4_or0));
  and_gate and_gate_u_csamul_cska32_and4_4(.a(a[4]), .b(b[4]), .out(u_csamul_cska32_and4_4));
  fa fa_u_csamul_cska32_fa4_4_out(.a(u_csamul_cska32_and4_4[0]), .b(u_csamul_cska32_fa5_3_xor1[0]), .cin(u_csamul_cska32_fa4_3_or0[0]), .fa_xor1(u_csamul_cska32_fa4_4_xor1), .fa_or0(u_csamul_cska32_fa4_4_or0));
  and_gate and_gate_u_csamul_cska32_and5_4(.a(a[5]), .b(b[4]), .out(u_csamul_cska32_and5_4));
  fa fa_u_csamul_cska32_fa5_4_out(.a(u_csamul_cska32_and5_4[0]), .b(u_csamul_cska32_fa6_3_xor1[0]), .cin(u_csamul_cska32_fa5_3_or0[0]), .fa_xor1(u_csamul_cska32_fa5_4_xor1), .fa_or0(u_csamul_cska32_fa5_4_or0));
  and_gate and_gate_u_csamul_cska32_and6_4(.a(a[6]), .b(b[4]), .out(u_csamul_cska32_and6_4));
  fa fa_u_csamul_cska32_fa6_4_out(.a(u_csamul_cska32_and6_4[0]), .b(u_csamul_cska32_fa7_3_xor1[0]), .cin(u_csamul_cska32_fa6_3_or0[0]), .fa_xor1(u_csamul_cska32_fa6_4_xor1), .fa_or0(u_csamul_cska32_fa6_4_or0));
  and_gate and_gate_u_csamul_cska32_and7_4(.a(a[7]), .b(b[4]), .out(u_csamul_cska32_and7_4));
  fa fa_u_csamul_cska32_fa7_4_out(.a(u_csamul_cska32_and7_4[0]), .b(u_csamul_cska32_fa8_3_xor1[0]), .cin(u_csamul_cska32_fa7_3_or0[0]), .fa_xor1(u_csamul_cska32_fa7_4_xor1), .fa_or0(u_csamul_cska32_fa7_4_or0));
  and_gate and_gate_u_csamul_cska32_and8_4(.a(a[8]), .b(b[4]), .out(u_csamul_cska32_and8_4));
  fa fa_u_csamul_cska32_fa8_4_out(.a(u_csamul_cska32_and8_4[0]), .b(u_csamul_cska32_fa9_3_xor1[0]), .cin(u_csamul_cska32_fa8_3_or0[0]), .fa_xor1(u_csamul_cska32_fa8_4_xor1), .fa_or0(u_csamul_cska32_fa8_4_or0));
  and_gate and_gate_u_csamul_cska32_and9_4(.a(a[9]), .b(b[4]), .out(u_csamul_cska32_and9_4));
  fa fa_u_csamul_cska32_fa9_4_out(.a(u_csamul_cska32_and9_4[0]), .b(u_csamul_cska32_fa10_3_xor1[0]), .cin(u_csamul_cska32_fa9_3_or0[0]), .fa_xor1(u_csamul_cska32_fa9_4_xor1), .fa_or0(u_csamul_cska32_fa9_4_or0));
  and_gate and_gate_u_csamul_cska32_and10_4(.a(a[10]), .b(b[4]), .out(u_csamul_cska32_and10_4));
  fa fa_u_csamul_cska32_fa10_4_out(.a(u_csamul_cska32_and10_4[0]), .b(u_csamul_cska32_fa11_3_xor1[0]), .cin(u_csamul_cska32_fa10_3_or0[0]), .fa_xor1(u_csamul_cska32_fa10_4_xor1), .fa_or0(u_csamul_cska32_fa10_4_or0));
  and_gate and_gate_u_csamul_cska32_and11_4(.a(a[11]), .b(b[4]), .out(u_csamul_cska32_and11_4));
  fa fa_u_csamul_cska32_fa11_4_out(.a(u_csamul_cska32_and11_4[0]), .b(u_csamul_cska32_fa12_3_xor1[0]), .cin(u_csamul_cska32_fa11_3_or0[0]), .fa_xor1(u_csamul_cska32_fa11_4_xor1), .fa_or0(u_csamul_cska32_fa11_4_or0));
  and_gate and_gate_u_csamul_cska32_and12_4(.a(a[12]), .b(b[4]), .out(u_csamul_cska32_and12_4));
  fa fa_u_csamul_cska32_fa12_4_out(.a(u_csamul_cska32_and12_4[0]), .b(u_csamul_cska32_fa13_3_xor1[0]), .cin(u_csamul_cska32_fa12_3_or0[0]), .fa_xor1(u_csamul_cska32_fa12_4_xor1), .fa_or0(u_csamul_cska32_fa12_4_or0));
  and_gate and_gate_u_csamul_cska32_and13_4(.a(a[13]), .b(b[4]), .out(u_csamul_cska32_and13_4));
  fa fa_u_csamul_cska32_fa13_4_out(.a(u_csamul_cska32_and13_4[0]), .b(u_csamul_cska32_fa14_3_xor1[0]), .cin(u_csamul_cska32_fa13_3_or0[0]), .fa_xor1(u_csamul_cska32_fa13_4_xor1), .fa_or0(u_csamul_cska32_fa13_4_or0));
  and_gate and_gate_u_csamul_cska32_and14_4(.a(a[14]), .b(b[4]), .out(u_csamul_cska32_and14_4));
  fa fa_u_csamul_cska32_fa14_4_out(.a(u_csamul_cska32_and14_4[0]), .b(u_csamul_cska32_fa15_3_xor1[0]), .cin(u_csamul_cska32_fa14_3_or0[0]), .fa_xor1(u_csamul_cska32_fa14_4_xor1), .fa_or0(u_csamul_cska32_fa14_4_or0));
  and_gate and_gate_u_csamul_cska32_and15_4(.a(a[15]), .b(b[4]), .out(u_csamul_cska32_and15_4));
  fa fa_u_csamul_cska32_fa15_4_out(.a(u_csamul_cska32_and15_4[0]), .b(u_csamul_cska32_fa16_3_xor1[0]), .cin(u_csamul_cska32_fa15_3_or0[0]), .fa_xor1(u_csamul_cska32_fa15_4_xor1), .fa_or0(u_csamul_cska32_fa15_4_or0));
  and_gate and_gate_u_csamul_cska32_and16_4(.a(a[16]), .b(b[4]), .out(u_csamul_cska32_and16_4));
  fa fa_u_csamul_cska32_fa16_4_out(.a(u_csamul_cska32_and16_4[0]), .b(u_csamul_cska32_fa17_3_xor1[0]), .cin(u_csamul_cska32_fa16_3_or0[0]), .fa_xor1(u_csamul_cska32_fa16_4_xor1), .fa_or0(u_csamul_cska32_fa16_4_or0));
  and_gate and_gate_u_csamul_cska32_and17_4(.a(a[17]), .b(b[4]), .out(u_csamul_cska32_and17_4));
  fa fa_u_csamul_cska32_fa17_4_out(.a(u_csamul_cska32_and17_4[0]), .b(u_csamul_cska32_fa18_3_xor1[0]), .cin(u_csamul_cska32_fa17_3_or0[0]), .fa_xor1(u_csamul_cska32_fa17_4_xor1), .fa_or0(u_csamul_cska32_fa17_4_or0));
  and_gate and_gate_u_csamul_cska32_and18_4(.a(a[18]), .b(b[4]), .out(u_csamul_cska32_and18_4));
  fa fa_u_csamul_cska32_fa18_4_out(.a(u_csamul_cska32_and18_4[0]), .b(u_csamul_cska32_fa19_3_xor1[0]), .cin(u_csamul_cska32_fa18_3_or0[0]), .fa_xor1(u_csamul_cska32_fa18_4_xor1), .fa_or0(u_csamul_cska32_fa18_4_or0));
  and_gate and_gate_u_csamul_cska32_and19_4(.a(a[19]), .b(b[4]), .out(u_csamul_cska32_and19_4));
  fa fa_u_csamul_cska32_fa19_4_out(.a(u_csamul_cska32_and19_4[0]), .b(u_csamul_cska32_fa20_3_xor1[0]), .cin(u_csamul_cska32_fa19_3_or0[0]), .fa_xor1(u_csamul_cska32_fa19_4_xor1), .fa_or0(u_csamul_cska32_fa19_4_or0));
  and_gate and_gate_u_csamul_cska32_and20_4(.a(a[20]), .b(b[4]), .out(u_csamul_cska32_and20_4));
  fa fa_u_csamul_cska32_fa20_4_out(.a(u_csamul_cska32_and20_4[0]), .b(u_csamul_cska32_fa21_3_xor1[0]), .cin(u_csamul_cska32_fa20_3_or0[0]), .fa_xor1(u_csamul_cska32_fa20_4_xor1), .fa_or0(u_csamul_cska32_fa20_4_or0));
  and_gate and_gate_u_csamul_cska32_and21_4(.a(a[21]), .b(b[4]), .out(u_csamul_cska32_and21_4));
  fa fa_u_csamul_cska32_fa21_4_out(.a(u_csamul_cska32_and21_4[0]), .b(u_csamul_cska32_fa22_3_xor1[0]), .cin(u_csamul_cska32_fa21_3_or0[0]), .fa_xor1(u_csamul_cska32_fa21_4_xor1), .fa_or0(u_csamul_cska32_fa21_4_or0));
  and_gate and_gate_u_csamul_cska32_and22_4(.a(a[22]), .b(b[4]), .out(u_csamul_cska32_and22_4));
  fa fa_u_csamul_cska32_fa22_4_out(.a(u_csamul_cska32_and22_4[0]), .b(u_csamul_cska32_fa23_3_xor1[0]), .cin(u_csamul_cska32_fa22_3_or0[0]), .fa_xor1(u_csamul_cska32_fa22_4_xor1), .fa_or0(u_csamul_cska32_fa22_4_or0));
  and_gate and_gate_u_csamul_cska32_and23_4(.a(a[23]), .b(b[4]), .out(u_csamul_cska32_and23_4));
  fa fa_u_csamul_cska32_fa23_4_out(.a(u_csamul_cska32_and23_4[0]), .b(u_csamul_cska32_fa24_3_xor1[0]), .cin(u_csamul_cska32_fa23_3_or0[0]), .fa_xor1(u_csamul_cska32_fa23_4_xor1), .fa_or0(u_csamul_cska32_fa23_4_or0));
  and_gate and_gate_u_csamul_cska32_and24_4(.a(a[24]), .b(b[4]), .out(u_csamul_cska32_and24_4));
  fa fa_u_csamul_cska32_fa24_4_out(.a(u_csamul_cska32_and24_4[0]), .b(u_csamul_cska32_fa25_3_xor1[0]), .cin(u_csamul_cska32_fa24_3_or0[0]), .fa_xor1(u_csamul_cska32_fa24_4_xor1), .fa_or0(u_csamul_cska32_fa24_4_or0));
  and_gate and_gate_u_csamul_cska32_and25_4(.a(a[25]), .b(b[4]), .out(u_csamul_cska32_and25_4));
  fa fa_u_csamul_cska32_fa25_4_out(.a(u_csamul_cska32_and25_4[0]), .b(u_csamul_cska32_fa26_3_xor1[0]), .cin(u_csamul_cska32_fa25_3_or0[0]), .fa_xor1(u_csamul_cska32_fa25_4_xor1), .fa_or0(u_csamul_cska32_fa25_4_or0));
  and_gate and_gate_u_csamul_cska32_and26_4(.a(a[26]), .b(b[4]), .out(u_csamul_cska32_and26_4));
  fa fa_u_csamul_cska32_fa26_4_out(.a(u_csamul_cska32_and26_4[0]), .b(u_csamul_cska32_fa27_3_xor1[0]), .cin(u_csamul_cska32_fa26_3_or0[0]), .fa_xor1(u_csamul_cska32_fa26_4_xor1), .fa_or0(u_csamul_cska32_fa26_4_or0));
  and_gate and_gate_u_csamul_cska32_and27_4(.a(a[27]), .b(b[4]), .out(u_csamul_cska32_and27_4));
  fa fa_u_csamul_cska32_fa27_4_out(.a(u_csamul_cska32_and27_4[0]), .b(u_csamul_cska32_fa28_3_xor1[0]), .cin(u_csamul_cska32_fa27_3_or0[0]), .fa_xor1(u_csamul_cska32_fa27_4_xor1), .fa_or0(u_csamul_cska32_fa27_4_or0));
  and_gate and_gate_u_csamul_cska32_and28_4(.a(a[28]), .b(b[4]), .out(u_csamul_cska32_and28_4));
  fa fa_u_csamul_cska32_fa28_4_out(.a(u_csamul_cska32_and28_4[0]), .b(u_csamul_cska32_fa29_3_xor1[0]), .cin(u_csamul_cska32_fa28_3_or0[0]), .fa_xor1(u_csamul_cska32_fa28_4_xor1), .fa_or0(u_csamul_cska32_fa28_4_or0));
  and_gate and_gate_u_csamul_cska32_and29_4(.a(a[29]), .b(b[4]), .out(u_csamul_cska32_and29_4));
  fa fa_u_csamul_cska32_fa29_4_out(.a(u_csamul_cska32_and29_4[0]), .b(u_csamul_cska32_fa30_3_xor1[0]), .cin(u_csamul_cska32_fa29_3_or0[0]), .fa_xor1(u_csamul_cska32_fa29_4_xor1), .fa_or0(u_csamul_cska32_fa29_4_or0));
  and_gate and_gate_u_csamul_cska32_and30_4(.a(a[30]), .b(b[4]), .out(u_csamul_cska32_and30_4));
  fa fa_u_csamul_cska32_fa30_4_out(.a(u_csamul_cska32_and30_4[0]), .b(u_csamul_cska32_and31_3[0]), .cin(u_csamul_cska32_fa30_3_or0[0]), .fa_xor1(u_csamul_cska32_fa30_4_xor1), .fa_or0(u_csamul_cska32_fa30_4_or0));
  and_gate and_gate_u_csamul_cska32_and31_4(.a(a[31]), .b(b[4]), .out(u_csamul_cska32_and31_4));
  and_gate and_gate_u_csamul_cska32_and0_5(.a(a[0]), .b(b[5]), .out(u_csamul_cska32_and0_5));
  fa fa_u_csamul_cska32_fa0_5_out(.a(u_csamul_cska32_and0_5[0]), .b(u_csamul_cska32_fa1_4_xor1[0]), .cin(u_csamul_cska32_fa0_4_or0[0]), .fa_xor1(u_csamul_cska32_fa0_5_xor1), .fa_or0(u_csamul_cska32_fa0_5_or0));
  and_gate and_gate_u_csamul_cska32_and1_5(.a(a[1]), .b(b[5]), .out(u_csamul_cska32_and1_5));
  fa fa_u_csamul_cska32_fa1_5_out(.a(u_csamul_cska32_and1_5[0]), .b(u_csamul_cska32_fa2_4_xor1[0]), .cin(u_csamul_cska32_fa1_4_or0[0]), .fa_xor1(u_csamul_cska32_fa1_5_xor1), .fa_or0(u_csamul_cska32_fa1_5_or0));
  and_gate and_gate_u_csamul_cska32_and2_5(.a(a[2]), .b(b[5]), .out(u_csamul_cska32_and2_5));
  fa fa_u_csamul_cska32_fa2_5_out(.a(u_csamul_cska32_and2_5[0]), .b(u_csamul_cska32_fa3_4_xor1[0]), .cin(u_csamul_cska32_fa2_4_or0[0]), .fa_xor1(u_csamul_cska32_fa2_5_xor1), .fa_or0(u_csamul_cska32_fa2_5_or0));
  and_gate and_gate_u_csamul_cska32_and3_5(.a(a[3]), .b(b[5]), .out(u_csamul_cska32_and3_5));
  fa fa_u_csamul_cska32_fa3_5_out(.a(u_csamul_cska32_and3_5[0]), .b(u_csamul_cska32_fa4_4_xor1[0]), .cin(u_csamul_cska32_fa3_4_or0[0]), .fa_xor1(u_csamul_cska32_fa3_5_xor1), .fa_or0(u_csamul_cska32_fa3_5_or0));
  and_gate and_gate_u_csamul_cska32_and4_5(.a(a[4]), .b(b[5]), .out(u_csamul_cska32_and4_5));
  fa fa_u_csamul_cska32_fa4_5_out(.a(u_csamul_cska32_and4_5[0]), .b(u_csamul_cska32_fa5_4_xor1[0]), .cin(u_csamul_cska32_fa4_4_or0[0]), .fa_xor1(u_csamul_cska32_fa4_5_xor1), .fa_or0(u_csamul_cska32_fa4_5_or0));
  and_gate and_gate_u_csamul_cska32_and5_5(.a(a[5]), .b(b[5]), .out(u_csamul_cska32_and5_5));
  fa fa_u_csamul_cska32_fa5_5_out(.a(u_csamul_cska32_and5_5[0]), .b(u_csamul_cska32_fa6_4_xor1[0]), .cin(u_csamul_cska32_fa5_4_or0[0]), .fa_xor1(u_csamul_cska32_fa5_5_xor1), .fa_or0(u_csamul_cska32_fa5_5_or0));
  and_gate and_gate_u_csamul_cska32_and6_5(.a(a[6]), .b(b[5]), .out(u_csamul_cska32_and6_5));
  fa fa_u_csamul_cska32_fa6_5_out(.a(u_csamul_cska32_and6_5[0]), .b(u_csamul_cska32_fa7_4_xor1[0]), .cin(u_csamul_cska32_fa6_4_or0[0]), .fa_xor1(u_csamul_cska32_fa6_5_xor1), .fa_or0(u_csamul_cska32_fa6_5_or0));
  and_gate and_gate_u_csamul_cska32_and7_5(.a(a[7]), .b(b[5]), .out(u_csamul_cska32_and7_5));
  fa fa_u_csamul_cska32_fa7_5_out(.a(u_csamul_cska32_and7_5[0]), .b(u_csamul_cska32_fa8_4_xor1[0]), .cin(u_csamul_cska32_fa7_4_or0[0]), .fa_xor1(u_csamul_cska32_fa7_5_xor1), .fa_or0(u_csamul_cska32_fa7_5_or0));
  and_gate and_gate_u_csamul_cska32_and8_5(.a(a[8]), .b(b[5]), .out(u_csamul_cska32_and8_5));
  fa fa_u_csamul_cska32_fa8_5_out(.a(u_csamul_cska32_and8_5[0]), .b(u_csamul_cska32_fa9_4_xor1[0]), .cin(u_csamul_cska32_fa8_4_or0[0]), .fa_xor1(u_csamul_cska32_fa8_5_xor1), .fa_or0(u_csamul_cska32_fa8_5_or0));
  and_gate and_gate_u_csamul_cska32_and9_5(.a(a[9]), .b(b[5]), .out(u_csamul_cska32_and9_5));
  fa fa_u_csamul_cska32_fa9_5_out(.a(u_csamul_cska32_and9_5[0]), .b(u_csamul_cska32_fa10_4_xor1[0]), .cin(u_csamul_cska32_fa9_4_or0[0]), .fa_xor1(u_csamul_cska32_fa9_5_xor1), .fa_or0(u_csamul_cska32_fa9_5_or0));
  and_gate and_gate_u_csamul_cska32_and10_5(.a(a[10]), .b(b[5]), .out(u_csamul_cska32_and10_5));
  fa fa_u_csamul_cska32_fa10_5_out(.a(u_csamul_cska32_and10_5[0]), .b(u_csamul_cska32_fa11_4_xor1[0]), .cin(u_csamul_cska32_fa10_4_or0[0]), .fa_xor1(u_csamul_cska32_fa10_5_xor1), .fa_or0(u_csamul_cska32_fa10_5_or0));
  and_gate and_gate_u_csamul_cska32_and11_5(.a(a[11]), .b(b[5]), .out(u_csamul_cska32_and11_5));
  fa fa_u_csamul_cska32_fa11_5_out(.a(u_csamul_cska32_and11_5[0]), .b(u_csamul_cska32_fa12_4_xor1[0]), .cin(u_csamul_cska32_fa11_4_or0[0]), .fa_xor1(u_csamul_cska32_fa11_5_xor1), .fa_or0(u_csamul_cska32_fa11_5_or0));
  and_gate and_gate_u_csamul_cska32_and12_5(.a(a[12]), .b(b[5]), .out(u_csamul_cska32_and12_5));
  fa fa_u_csamul_cska32_fa12_5_out(.a(u_csamul_cska32_and12_5[0]), .b(u_csamul_cska32_fa13_4_xor1[0]), .cin(u_csamul_cska32_fa12_4_or0[0]), .fa_xor1(u_csamul_cska32_fa12_5_xor1), .fa_or0(u_csamul_cska32_fa12_5_or0));
  and_gate and_gate_u_csamul_cska32_and13_5(.a(a[13]), .b(b[5]), .out(u_csamul_cska32_and13_5));
  fa fa_u_csamul_cska32_fa13_5_out(.a(u_csamul_cska32_and13_5[0]), .b(u_csamul_cska32_fa14_4_xor1[0]), .cin(u_csamul_cska32_fa13_4_or0[0]), .fa_xor1(u_csamul_cska32_fa13_5_xor1), .fa_or0(u_csamul_cska32_fa13_5_or0));
  and_gate and_gate_u_csamul_cska32_and14_5(.a(a[14]), .b(b[5]), .out(u_csamul_cska32_and14_5));
  fa fa_u_csamul_cska32_fa14_5_out(.a(u_csamul_cska32_and14_5[0]), .b(u_csamul_cska32_fa15_4_xor1[0]), .cin(u_csamul_cska32_fa14_4_or0[0]), .fa_xor1(u_csamul_cska32_fa14_5_xor1), .fa_or0(u_csamul_cska32_fa14_5_or0));
  and_gate and_gate_u_csamul_cska32_and15_5(.a(a[15]), .b(b[5]), .out(u_csamul_cska32_and15_5));
  fa fa_u_csamul_cska32_fa15_5_out(.a(u_csamul_cska32_and15_5[0]), .b(u_csamul_cska32_fa16_4_xor1[0]), .cin(u_csamul_cska32_fa15_4_or0[0]), .fa_xor1(u_csamul_cska32_fa15_5_xor1), .fa_or0(u_csamul_cska32_fa15_5_or0));
  and_gate and_gate_u_csamul_cska32_and16_5(.a(a[16]), .b(b[5]), .out(u_csamul_cska32_and16_5));
  fa fa_u_csamul_cska32_fa16_5_out(.a(u_csamul_cska32_and16_5[0]), .b(u_csamul_cska32_fa17_4_xor1[0]), .cin(u_csamul_cska32_fa16_4_or0[0]), .fa_xor1(u_csamul_cska32_fa16_5_xor1), .fa_or0(u_csamul_cska32_fa16_5_or0));
  and_gate and_gate_u_csamul_cska32_and17_5(.a(a[17]), .b(b[5]), .out(u_csamul_cska32_and17_5));
  fa fa_u_csamul_cska32_fa17_5_out(.a(u_csamul_cska32_and17_5[0]), .b(u_csamul_cska32_fa18_4_xor1[0]), .cin(u_csamul_cska32_fa17_4_or0[0]), .fa_xor1(u_csamul_cska32_fa17_5_xor1), .fa_or0(u_csamul_cska32_fa17_5_or0));
  and_gate and_gate_u_csamul_cska32_and18_5(.a(a[18]), .b(b[5]), .out(u_csamul_cska32_and18_5));
  fa fa_u_csamul_cska32_fa18_5_out(.a(u_csamul_cska32_and18_5[0]), .b(u_csamul_cska32_fa19_4_xor1[0]), .cin(u_csamul_cska32_fa18_4_or0[0]), .fa_xor1(u_csamul_cska32_fa18_5_xor1), .fa_or0(u_csamul_cska32_fa18_5_or0));
  and_gate and_gate_u_csamul_cska32_and19_5(.a(a[19]), .b(b[5]), .out(u_csamul_cska32_and19_5));
  fa fa_u_csamul_cska32_fa19_5_out(.a(u_csamul_cska32_and19_5[0]), .b(u_csamul_cska32_fa20_4_xor1[0]), .cin(u_csamul_cska32_fa19_4_or0[0]), .fa_xor1(u_csamul_cska32_fa19_5_xor1), .fa_or0(u_csamul_cska32_fa19_5_or0));
  and_gate and_gate_u_csamul_cska32_and20_5(.a(a[20]), .b(b[5]), .out(u_csamul_cska32_and20_5));
  fa fa_u_csamul_cska32_fa20_5_out(.a(u_csamul_cska32_and20_5[0]), .b(u_csamul_cska32_fa21_4_xor1[0]), .cin(u_csamul_cska32_fa20_4_or0[0]), .fa_xor1(u_csamul_cska32_fa20_5_xor1), .fa_or0(u_csamul_cska32_fa20_5_or0));
  and_gate and_gate_u_csamul_cska32_and21_5(.a(a[21]), .b(b[5]), .out(u_csamul_cska32_and21_5));
  fa fa_u_csamul_cska32_fa21_5_out(.a(u_csamul_cska32_and21_5[0]), .b(u_csamul_cska32_fa22_4_xor1[0]), .cin(u_csamul_cska32_fa21_4_or0[0]), .fa_xor1(u_csamul_cska32_fa21_5_xor1), .fa_or0(u_csamul_cska32_fa21_5_or0));
  and_gate and_gate_u_csamul_cska32_and22_5(.a(a[22]), .b(b[5]), .out(u_csamul_cska32_and22_5));
  fa fa_u_csamul_cska32_fa22_5_out(.a(u_csamul_cska32_and22_5[0]), .b(u_csamul_cska32_fa23_4_xor1[0]), .cin(u_csamul_cska32_fa22_4_or0[0]), .fa_xor1(u_csamul_cska32_fa22_5_xor1), .fa_or0(u_csamul_cska32_fa22_5_or0));
  and_gate and_gate_u_csamul_cska32_and23_5(.a(a[23]), .b(b[5]), .out(u_csamul_cska32_and23_5));
  fa fa_u_csamul_cska32_fa23_5_out(.a(u_csamul_cska32_and23_5[0]), .b(u_csamul_cska32_fa24_4_xor1[0]), .cin(u_csamul_cska32_fa23_4_or0[0]), .fa_xor1(u_csamul_cska32_fa23_5_xor1), .fa_or0(u_csamul_cska32_fa23_5_or0));
  and_gate and_gate_u_csamul_cska32_and24_5(.a(a[24]), .b(b[5]), .out(u_csamul_cska32_and24_5));
  fa fa_u_csamul_cska32_fa24_5_out(.a(u_csamul_cska32_and24_5[0]), .b(u_csamul_cska32_fa25_4_xor1[0]), .cin(u_csamul_cska32_fa24_4_or0[0]), .fa_xor1(u_csamul_cska32_fa24_5_xor1), .fa_or0(u_csamul_cska32_fa24_5_or0));
  and_gate and_gate_u_csamul_cska32_and25_5(.a(a[25]), .b(b[5]), .out(u_csamul_cska32_and25_5));
  fa fa_u_csamul_cska32_fa25_5_out(.a(u_csamul_cska32_and25_5[0]), .b(u_csamul_cska32_fa26_4_xor1[0]), .cin(u_csamul_cska32_fa25_4_or0[0]), .fa_xor1(u_csamul_cska32_fa25_5_xor1), .fa_or0(u_csamul_cska32_fa25_5_or0));
  and_gate and_gate_u_csamul_cska32_and26_5(.a(a[26]), .b(b[5]), .out(u_csamul_cska32_and26_5));
  fa fa_u_csamul_cska32_fa26_5_out(.a(u_csamul_cska32_and26_5[0]), .b(u_csamul_cska32_fa27_4_xor1[0]), .cin(u_csamul_cska32_fa26_4_or0[0]), .fa_xor1(u_csamul_cska32_fa26_5_xor1), .fa_or0(u_csamul_cska32_fa26_5_or0));
  and_gate and_gate_u_csamul_cska32_and27_5(.a(a[27]), .b(b[5]), .out(u_csamul_cska32_and27_5));
  fa fa_u_csamul_cska32_fa27_5_out(.a(u_csamul_cska32_and27_5[0]), .b(u_csamul_cska32_fa28_4_xor1[0]), .cin(u_csamul_cska32_fa27_4_or0[0]), .fa_xor1(u_csamul_cska32_fa27_5_xor1), .fa_or0(u_csamul_cska32_fa27_5_or0));
  and_gate and_gate_u_csamul_cska32_and28_5(.a(a[28]), .b(b[5]), .out(u_csamul_cska32_and28_5));
  fa fa_u_csamul_cska32_fa28_5_out(.a(u_csamul_cska32_and28_5[0]), .b(u_csamul_cska32_fa29_4_xor1[0]), .cin(u_csamul_cska32_fa28_4_or0[0]), .fa_xor1(u_csamul_cska32_fa28_5_xor1), .fa_or0(u_csamul_cska32_fa28_5_or0));
  and_gate and_gate_u_csamul_cska32_and29_5(.a(a[29]), .b(b[5]), .out(u_csamul_cska32_and29_5));
  fa fa_u_csamul_cska32_fa29_5_out(.a(u_csamul_cska32_and29_5[0]), .b(u_csamul_cska32_fa30_4_xor1[0]), .cin(u_csamul_cska32_fa29_4_or0[0]), .fa_xor1(u_csamul_cska32_fa29_5_xor1), .fa_or0(u_csamul_cska32_fa29_5_or0));
  and_gate and_gate_u_csamul_cska32_and30_5(.a(a[30]), .b(b[5]), .out(u_csamul_cska32_and30_5));
  fa fa_u_csamul_cska32_fa30_5_out(.a(u_csamul_cska32_and30_5[0]), .b(u_csamul_cska32_and31_4[0]), .cin(u_csamul_cska32_fa30_4_or0[0]), .fa_xor1(u_csamul_cska32_fa30_5_xor1), .fa_or0(u_csamul_cska32_fa30_5_or0));
  and_gate and_gate_u_csamul_cska32_and31_5(.a(a[31]), .b(b[5]), .out(u_csamul_cska32_and31_5));
  and_gate and_gate_u_csamul_cska32_and0_6(.a(a[0]), .b(b[6]), .out(u_csamul_cska32_and0_6));
  fa fa_u_csamul_cska32_fa0_6_out(.a(u_csamul_cska32_and0_6[0]), .b(u_csamul_cska32_fa1_5_xor1[0]), .cin(u_csamul_cska32_fa0_5_or0[0]), .fa_xor1(u_csamul_cska32_fa0_6_xor1), .fa_or0(u_csamul_cska32_fa0_6_or0));
  and_gate and_gate_u_csamul_cska32_and1_6(.a(a[1]), .b(b[6]), .out(u_csamul_cska32_and1_6));
  fa fa_u_csamul_cska32_fa1_6_out(.a(u_csamul_cska32_and1_6[0]), .b(u_csamul_cska32_fa2_5_xor1[0]), .cin(u_csamul_cska32_fa1_5_or0[0]), .fa_xor1(u_csamul_cska32_fa1_6_xor1), .fa_or0(u_csamul_cska32_fa1_6_or0));
  and_gate and_gate_u_csamul_cska32_and2_6(.a(a[2]), .b(b[6]), .out(u_csamul_cska32_and2_6));
  fa fa_u_csamul_cska32_fa2_6_out(.a(u_csamul_cska32_and2_6[0]), .b(u_csamul_cska32_fa3_5_xor1[0]), .cin(u_csamul_cska32_fa2_5_or0[0]), .fa_xor1(u_csamul_cska32_fa2_6_xor1), .fa_or0(u_csamul_cska32_fa2_6_or0));
  and_gate and_gate_u_csamul_cska32_and3_6(.a(a[3]), .b(b[6]), .out(u_csamul_cska32_and3_6));
  fa fa_u_csamul_cska32_fa3_6_out(.a(u_csamul_cska32_and3_6[0]), .b(u_csamul_cska32_fa4_5_xor1[0]), .cin(u_csamul_cska32_fa3_5_or0[0]), .fa_xor1(u_csamul_cska32_fa3_6_xor1), .fa_or0(u_csamul_cska32_fa3_6_or0));
  and_gate and_gate_u_csamul_cska32_and4_6(.a(a[4]), .b(b[6]), .out(u_csamul_cska32_and4_6));
  fa fa_u_csamul_cska32_fa4_6_out(.a(u_csamul_cska32_and4_6[0]), .b(u_csamul_cska32_fa5_5_xor1[0]), .cin(u_csamul_cska32_fa4_5_or0[0]), .fa_xor1(u_csamul_cska32_fa4_6_xor1), .fa_or0(u_csamul_cska32_fa4_6_or0));
  and_gate and_gate_u_csamul_cska32_and5_6(.a(a[5]), .b(b[6]), .out(u_csamul_cska32_and5_6));
  fa fa_u_csamul_cska32_fa5_6_out(.a(u_csamul_cska32_and5_6[0]), .b(u_csamul_cska32_fa6_5_xor1[0]), .cin(u_csamul_cska32_fa5_5_or0[0]), .fa_xor1(u_csamul_cska32_fa5_6_xor1), .fa_or0(u_csamul_cska32_fa5_6_or0));
  and_gate and_gate_u_csamul_cska32_and6_6(.a(a[6]), .b(b[6]), .out(u_csamul_cska32_and6_6));
  fa fa_u_csamul_cska32_fa6_6_out(.a(u_csamul_cska32_and6_6[0]), .b(u_csamul_cska32_fa7_5_xor1[0]), .cin(u_csamul_cska32_fa6_5_or0[0]), .fa_xor1(u_csamul_cska32_fa6_6_xor1), .fa_or0(u_csamul_cska32_fa6_6_or0));
  and_gate and_gate_u_csamul_cska32_and7_6(.a(a[7]), .b(b[6]), .out(u_csamul_cska32_and7_6));
  fa fa_u_csamul_cska32_fa7_6_out(.a(u_csamul_cska32_and7_6[0]), .b(u_csamul_cska32_fa8_5_xor1[0]), .cin(u_csamul_cska32_fa7_5_or0[0]), .fa_xor1(u_csamul_cska32_fa7_6_xor1), .fa_or0(u_csamul_cska32_fa7_6_or0));
  and_gate and_gate_u_csamul_cska32_and8_6(.a(a[8]), .b(b[6]), .out(u_csamul_cska32_and8_6));
  fa fa_u_csamul_cska32_fa8_6_out(.a(u_csamul_cska32_and8_6[0]), .b(u_csamul_cska32_fa9_5_xor1[0]), .cin(u_csamul_cska32_fa8_5_or0[0]), .fa_xor1(u_csamul_cska32_fa8_6_xor1), .fa_or0(u_csamul_cska32_fa8_6_or0));
  and_gate and_gate_u_csamul_cska32_and9_6(.a(a[9]), .b(b[6]), .out(u_csamul_cska32_and9_6));
  fa fa_u_csamul_cska32_fa9_6_out(.a(u_csamul_cska32_and9_6[0]), .b(u_csamul_cska32_fa10_5_xor1[0]), .cin(u_csamul_cska32_fa9_5_or0[0]), .fa_xor1(u_csamul_cska32_fa9_6_xor1), .fa_or0(u_csamul_cska32_fa9_6_or0));
  and_gate and_gate_u_csamul_cska32_and10_6(.a(a[10]), .b(b[6]), .out(u_csamul_cska32_and10_6));
  fa fa_u_csamul_cska32_fa10_6_out(.a(u_csamul_cska32_and10_6[0]), .b(u_csamul_cska32_fa11_5_xor1[0]), .cin(u_csamul_cska32_fa10_5_or0[0]), .fa_xor1(u_csamul_cska32_fa10_6_xor1), .fa_or0(u_csamul_cska32_fa10_6_or0));
  and_gate and_gate_u_csamul_cska32_and11_6(.a(a[11]), .b(b[6]), .out(u_csamul_cska32_and11_6));
  fa fa_u_csamul_cska32_fa11_6_out(.a(u_csamul_cska32_and11_6[0]), .b(u_csamul_cska32_fa12_5_xor1[0]), .cin(u_csamul_cska32_fa11_5_or0[0]), .fa_xor1(u_csamul_cska32_fa11_6_xor1), .fa_or0(u_csamul_cska32_fa11_6_or0));
  and_gate and_gate_u_csamul_cska32_and12_6(.a(a[12]), .b(b[6]), .out(u_csamul_cska32_and12_6));
  fa fa_u_csamul_cska32_fa12_6_out(.a(u_csamul_cska32_and12_6[0]), .b(u_csamul_cska32_fa13_5_xor1[0]), .cin(u_csamul_cska32_fa12_5_or0[0]), .fa_xor1(u_csamul_cska32_fa12_6_xor1), .fa_or0(u_csamul_cska32_fa12_6_or0));
  and_gate and_gate_u_csamul_cska32_and13_6(.a(a[13]), .b(b[6]), .out(u_csamul_cska32_and13_6));
  fa fa_u_csamul_cska32_fa13_6_out(.a(u_csamul_cska32_and13_6[0]), .b(u_csamul_cska32_fa14_5_xor1[0]), .cin(u_csamul_cska32_fa13_5_or0[0]), .fa_xor1(u_csamul_cska32_fa13_6_xor1), .fa_or0(u_csamul_cska32_fa13_6_or0));
  and_gate and_gate_u_csamul_cska32_and14_6(.a(a[14]), .b(b[6]), .out(u_csamul_cska32_and14_6));
  fa fa_u_csamul_cska32_fa14_6_out(.a(u_csamul_cska32_and14_6[0]), .b(u_csamul_cska32_fa15_5_xor1[0]), .cin(u_csamul_cska32_fa14_5_or0[0]), .fa_xor1(u_csamul_cska32_fa14_6_xor1), .fa_or0(u_csamul_cska32_fa14_6_or0));
  and_gate and_gate_u_csamul_cska32_and15_6(.a(a[15]), .b(b[6]), .out(u_csamul_cska32_and15_6));
  fa fa_u_csamul_cska32_fa15_6_out(.a(u_csamul_cska32_and15_6[0]), .b(u_csamul_cska32_fa16_5_xor1[0]), .cin(u_csamul_cska32_fa15_5_or0[0]), .fa_xor1(u_csamul_cska32_fa15_6_xor1), .fa_or0(u_csamul_cska32_fa15_6_or0));
  and_gate and_gate_u_csamul_cska32_and16_6(.a(a[16]), .b(b[6]), .out(u_csamul_cska32_and16_6));
  fa fa_u_csamul_cska32_fa16_6_out(.a(u_csamul_cska32_and16_6[0]), .b(u_csamul_cska32_fa17_5_xor1[0]), .cin(u_csamul_cska32_fa16_5_or0[0]), .fa_xor1(u_csamul_cska32_fa16_6_xor1), .fa_or0(u_csamul_cska32_fa16_6_or0));
  and_gate and_gate_u_csamul_cska32_and17_6(.a(a[17]), .b(b[6]), .out(u_csamul_cska32_and17_6));
  fa fa_u_csamul_cska32_fa17_6_out(.a(u_csamul_cska32_and17_6[0]), .b(u_csamul_cska32_fa18_5_xor1[0]), .cin(u_csamul_cska32_fa17_5_or0[0]), .fa_xor1(u_csamul_cska32_fa17_6_xor1), .fa_or0(u_csamul_cska32_fa17_6_or0));
  and_gate and_gate_u_csamul_cska32_and18_6(.a(a[18]), .b(b[6]), .out(u_csamul_cska32_and18_6));
  fa fa_u_csamul_cska32_fa18_6_out(.a(u_csamul_cska32_and18_6[0]), .b(u_csamul_cska32_fa19_5_xor1[0]), .cin(u_csamul_cska32_fa18_5_or0[0]), .fa_xor1(u_csamul_cska32_fa18_6_xor1), .fa_or0(u_csamul_cska32_fa18_6_or0));
  and_gate and_gate_u_csamul_cska32_and19_6(.a(a[19]), .b(b[6]), .out(u_csamul_cska32_and19_6));
  fa fa_u_csamul_cska32_fa19_6_out(.a(u_csamul_cska32_and19_6[0]), .b(u_csamul_cska32_fa20_5_xor1[0]), .cin(u_csamul_cska32_fa19_5_or0[0]), .fa_xor1(u_csamul_cska32_fa19_6_xor1), .fa_or0(u_csamul_cska32_fa19_6_or0));
  and_gate and_gate_u_csamul_cska32_and20_6(.a(a[20]), .b(b[6]), .out(u_csamul_cska32_and20_6));
  fa fa_u_csamul_cska32_fa20_6_out(.a(u_csamul_cska32_and20_6[0]), .b(u_csamul_cska32_fa21_5_xor1[0]), .cin(u_csamul_cska32_fa20_5_or0[0]), .fa_xor1(u_csamul_cska32_fa20_6_xor1), .fa_or0(u_csamul_cska32_fa20_6_or0));
  and_gate and_gate_u_csamul_cska32_and21_6(.a(a[21]), .b(b[6]), .out(u_csamul_cska32_and21_6));
  fa fa_u_csamul_cska32_fa21_6_out(.a(u_csamul_cska32_and21_6[0]), .b(u_csamul_cska32_fa22_5_xor1[0]), .cin(u_csamul_cska32_fa21_5_or0[0]), .fa_xor1(u_csamul_cska32_fa21_6_xor1), .fa_or0(u_csamul_cska32_fa21_6_or0));
  and_gate and_gate_u_csamul_cska32_and22_6(.a(a[22]), .b(b[6]), .out(u_csamul_cska32_and22_6));
  fa fa_u_csamul_cska32_fa22_6_out(.a(u_csamul_cska32_and22_6[0]), .b(u_csamul_cska32_fa23_5_xor1[0]), .cin(u_csamul_cska32_fa22_5_or0[0]), .fa_xor1(u_csamul_cska32_fa22_6_xor1), .fa_or0(u_csamul_cska32_fa22_6_or0));
  and_gate and_gate_u_csamul_cska32_and23_6(.a(a[23]), .b(b[6]), .out(u_csamul_cska32_and23_6));
  fa fa_u_csamul_cska32_fa23_6_out(.a(u_csamul_cska32_and23_6[0]), .b(u_csamul_cska32_fa24_5_xor1[0]), .cin(u_csamul_cska32_fa23_5_or0[0]), .fa_xor1(u_csamul_cska32_fa23_6_xor1), .fa_or0(u_csamul_cska32_fa23_6_or0));
  and_gate and_gate_u_csamul_cska32_and24_6(.a(a[24]), .b(b[6]), .out(u_csamul_cska32_and24_6));
  fa fa_u_csamul_cska32_fa24_6_out(.a(u_csamul_cska32_and24_6[0]), .b(u_csamul_cska32_fa25_5_xor1[0]), .cin(u_csamul_cska32_fa24_5_or0[0]), .fa_xor1(u_csamul_cska32_fa24_6_xor1), .fa_or0(u_csamul_cska32_fa24_6_or0));
  and_gate and_gate_u_csamul_cska32_and25_6(.a(a[25]), .b(b[6]), .out(u_csamul_cska32_and25_6));
  fa fa_u_csamul_cska32_fa25_6_out(.a(u_csamul_cska32_and25_6[0]), .b(u_csamul_cska32_fa26_5_xor1[0]), .cin(u_csamul_cska32_fa25_5_or0[0]), .fa_xor1(u_csamul_cska32_fa25_6_xor1), .fa_or0(u_csamul_cska32_fa25_6_or0));
  and_gate and_gate_u_csamul_cska32_and26_6(.a(a[26]), .b(b[6]), .out(u_csamul_cska32_and26_6));
  fa fa_u_csamul_cska32_fa26_6_out(.a(u_csamul_cska32_and26_6[0]), .b(u_csamul_cska32_fa27_5_xor1[0]), .cin(u_csamul_cska32_fa26_5_or0[0]), .fa_xor1(u_csamul_cska32_fa26_6_xor1), .fa_or0(u_csamul_cska32_fa26_6_or0));
  and_gate and_gate_u_csamul_cska32_and27_6(.a(a[27]), .b(b[6]), .out(u_csamul_cska32_and27_6));
  fa fa_u_csamul_cska32_fa27_6_out(.a(u_csamul_cska32_and27_6[0]), .b(u_csamul_cska32_fa28_5_xor1[0]), .cin(u_csamul_cska32_fa27_5_or0[0]), .fa_xor1(u_csamul_cska32_fa27_6_xor1), .fa_or0(u_csamul_cska32_fa27_6_or0));
  and_gate and_gate_u_csamul_cska32_and28_6(.a(a[28]), .b(b[6]), .out(u_csamul_cska32_and28_6));
  fa fa_u_csamul_cska32_fa28_6_out(.a(u_csamul_cska32_and28_6[0]), .b(u_csamul_cska32_fa29_5_xor1[0]), .cin(u_csamul_cska32_fa28_5_or0[0]), .fa_xor1(u_csamul_cska32_fa28_6_xor1), .fa_or0(u_csamul_cska32_fa28_6_or0));
  and_gate and_gate_u_csamul_cska32_and29_6(.a(a[29]), .b(b[6]), .out(u_csamul_cska32_and29_6));
  fa fa_u_csamul_cska32_fa29_6_out(.a(u_csamul_cska32_and29_6[0]), .b(u_csamul_cska32_fa30_5_xor1[0]), .cin(u_csamul_cska32_fa29_5_or0[0]), .fa_xor1(u_csamul_cska32_fa29_6_xor1), .fa_or0(u_csamul_cska32_fa29_6_or0));
  and_gate and_gate_u_csamul_cska32_and30_6(.a(a[30]), .b(b[6]), .out(u_csamul_cska32_and30_6));
  fa fa_u_csamul_cska32_fa30_6_out(.a(u_csamul_cska32_and30_6[0]), .b(u_csamul_cska32_and31_5[0]), .cin(u_csamul_cska32_fa30_5_or0[0]), .fa_xor1(u_csamul_cska32_fa30_6_xor1), .fa_or0(u_csamul_cska32_fa30_6_or0));
  and_gate and_gate_u_csamul_cska32_and31_6(.a(a[31]), .b(b[6]), .out(u_csamul_cska32_and31_6));
  and_gate and_gate_u_csamul_cska32_and0_7(.a(a[0]), .b(b[7]), .out(u_csamul_cska32_and0_7));
  fa fa_u_csamul_cska32_fa0_7_out(.a(u_csamul_cska32_and0_7[0]), .b(u_csamul_cska32_fa1_6_xor1[0]), .cin(u_csamul_cska32_fa0_6_or0[0]), .fa_xor1(u_csamul_cska32_fa0_7_xor1), .fa_or0(u_csamul_cska32_fa0_7_or0));
  and_gate and_gate_u_csamul_cska32_and1_7(.a(a[1]), .b(b[7]), .out(u_csamul_cska32_and1_7));
  fa fa_u_csamul_cska32_fa1_7_out(.a(u_csamul_cska32_and1_7[0]), .b(u_csamul_cska32_fa2_6_xor1[0]), .cin(u_csamul_cska32_fa1_6_or0[0]), .fa_xor1(u_csamul_cska32_fa1_7_xor1), .fa_or0(u_csamul_cska32_fa1_7_or0));
  and_gate and_gate_u_csamul_cska32_and2_7(.a(a[2]), .b(b[7]), .out(u_csamul_cska32_and2_7));
  fa fa_u_csamul_cska32_fa2_7_out(.a(u_csamul_cska32_and2_7[0]), .b(u_csamul_cska32_fa3_6_xor1[0]), .cin(u_csamul_cska32_fa2_6_or0[0]), .fa_xor1(u_csamul_cska32_fa2_7_xor1), .fa_or0(u_csamul_cska32_fa2_7_or0));
  and_gate and_gate_u_csamul_cska32_and3_7(.a(a[3]), .b(b[7]), .out(u_csamul_cska32_and3_7));
  fa fa_u_csamul_cska32_fa3_7_out(.a(u_csamul_cska32_and3_7[0]), .b(u_csamul_cska32_fa4_6_xor1[0]), .cin(u_csamul_cska32_fa3_6_or0[0]), .fa_xor1(u_csamul_cska32_fa3_7_xor1), .fa_or0(u_csamul_cska32_fa3_7_or0));
  and_gate and_gate_u_csamul_cska32_and4_7(.a(a[4]), .b(b[7]), .out(u_csamul_cska32_and4_7));
  fa fa_u_csamul_cska32_fa4_7_out(.a(u_csamul_cska32_and4_7[0]), .b(u_csamul_cska32_fa5_6_xor1[0]), .cin(u_csamul_cska32_fa4_6_or0[0]), .fa_xor1(u_csamul_cska32_fa4_7_xor1), .fa_or0(u_csamul_cska32_fa4_7_or0));
  and_gate and_gate_u_csamul_cska32_and5_7(.a(a[5]), .b(b[7]), .out(u_csamul_cska32_and5_7));
  fa fa_u_csamul_cska32_fa5_7_out(.a(u_csamul_cska32_and5_7[0]), .b(u_csamul_cska32_fa6_6_xor1[0]), .cin(u_csamul_cska32_fa5_6_or0[0]), .fa_xor1(u_csamul_cska32_fa5_7_xor1), .fa_or0(u_csamul_cska32_fa5_7_or0));
  and_gate and_gate_u_csamul_cska32_and6_7(.a(a[6]), .b(b[7]), .out(u_csamul_cska32_and6_7));
  fa fa_u_csamul_cska32_fa6_7_out(.a(u_csamul_cska32_and6_7[0]), .b(u_csamul_cska32_fa7_6_xor1[0]), .cin(u_csamul_cska32_fa6_6_or0[0]), .fa_xor1(u_csamul_cska32_fa6_7_xor1), .fa_or0(u_csamul_cska32_fa6_7_or0));
  and_gate and_gate_u_csamul_cska32_and7_7(.a(a[7]), .b(b[7]), .out(u_csamul_cska32_and7_7));
  fa fa_u_csamul_cska32_fa7_7_out(.a(u_csamul_cska32_and7_7[0]), .b(u_csamul_cska32_fa8_6_xor1[0]), .cin(u_csamul_cska32_fa7_6_or0[0]), .fa_xor1(u_csamul_cska32_fa7_7_xor1), .fa_or0(u_csamul_cska32_fa7_7_or0));
  and_gate and_gate_u_csamul_cska32_and8_7(.a(a[8]), .b(b[7]), .out(u_csamul_cska32_and8_7));
  fa fa_u_csamul_cska32_fa8_7_out(.a(u_csamul_cska32_and8_7[0]), .b(u_csamul_cska32_fa9_6_xor1[0]), .cin(u_csamul_cska32_fa8_6_or0[0]), .fa_xor1(u_csamul_cska32_fa8_7_xor1), .fa_or0(u_csamul_cska32_fa8_7_or0));
  and_gate and_gate_u_csamul_cska32_and9_7(.a(a[9]), .b(b[7]), .out(u_csamul_cska32_and9_7));
  fa fa_u_csamul_cska32_fa9_7_out(.a(u_csamul_cska32_and9_7[0]), .b(u_csamul_cska32_fa10_6_xor1[0]), .cin(u_csamul_cska32_fa9_6_or0[0]), .fa_xor1(u_csamul_cska32_fa9_7_xor1), .fa_or0(u_csamul_cska32_fa9_7_or0));
  and_gate and_gate_u_csamul_cska32_and10_7(.a(a[10]), .b(b[7]), .out(u_csamul_cska32_and10_7));
  fa fa_u_csamul_cska32_fa10_7_out(.a(u_csamul_cska32_and10_7[0]), .b(u_csamul_cska32_fa11_6_xor1[0]), .cin(u_csamul_cska32_fa10_6_or0[0]), .fa_xor1(u_csamul_cska32_fa10_7_xor1), .fa_or0(u_csamul_cska32_fa10_7_or0));
  and_gate and_gate_u_csamul_cska32_and11_7(.a(a[11]), .b(b[7]), .out(u_csamul_cska32_and11_7));
  fa fa_u_csamul_cska32_fa11_7_out(.a(u_csamul_cska32_and11_7[0]), .b(u_csamul_cska32_fa12_6_xor1[0]), .cin(u_csamul_cska32_fa11_6_or0[0]), .fa_xor1(u_csamul_cska32_fa11_7_xor1), .fa_or0(u_csamul_cska32_fa11_7_or0));
  and_gate and_gate_u_csamul_cska32_and12_7(.a(a[12]), .b(b[7]), .out(u_csamul_cska32_and12_7));
  fa fa_u_csamul_cska32_fa12_7_out(.a(u_csamul_cska32_and12_7[0]), .b(u_csamul_cska32_fa13_6_xor1[0]), .cin(u_csamul_cska32_fa12_6_or0[0]), .fa_xor1(u_csamul_cska32_fa12_7_xor1), .fa_or0(u_csamul_cska32_fa12_7_or0));
  and_gate and_gate_u_csamul_cska32_and13_7(.a(a[13]), .b(b[7]), .out(u_csamul_cska32_and13_7));
  fa fa_u_csamul_cska32_fa13_7_out(.a(u_csamul_cska32_and13_7[0]), .b(u_csamul_cska32_fa14_6_xor1[0]), .cin(u_csamul_cska32_fa13_6_or0[0]), .fa_xor1(u_csamul_cska32_fa13_7_xor1), .fa_or0(u_csamul_cska32_fa13_7_or0));
  and_gate and_gate_u_csamul_cska32_and14_7(.a(a[14]), .b(b[7]), .out(u_csamul_cska32_and14_7));
  fa fa_u_csamul_cska32_fa14_7_out(.a(u_csamul_cska32_and14_7[0]), .b(u_csamul_cska32_fa15_6_xor1[0]), .cin(u_csamul_cska32_fa14_6_or0[0]), .fa_xor1(u_csamul_cska32_fa14_7_xor1), .fa_or0(u_csamul_cska32_fa14_7_or0));
  and_gate and_gate_u_csamul_cska32_and15_7(.a(a[15]), .b(b[7]), .out(u_csamul_cska32_and15_7));
  fa fa_u_csamul_cska32_fa15_7_out(.a(u_csamul_cska32_and15_7[0]), .b(u_csamul_cska32_fa16_6_xor1[0]), .cin(u_csamul_cska32_fa15_6_or0[0]), .fa_xor1(u_csamul_cska32_fa15_7_xor1), .fa_or0(u_csamul_cska32_fa15_7_or0));
  and_gate and_gate_u_csamul_cska32_and16_7(.a(a[16]), .b(b[7]), .out(u_csamul_cska32_and16_7));
  fa fa_u_csamul_cska32_fa16_7_out(.a(u_csamul_cska32_and16_7[0]), .b(u_csamul_cska32_fa17_6_xor1[0]), .cin(u_csamul_cska32_fa16_6_or0[0]), .fa_xor1(u_csamul_cska32_fa16_7_xor1), .fa_or0(u_csamul_cska32_fa16_7_or0));
  and_gate and_gate_u_csamul_cska32_and17_7(.a(a[17]), .b(b[7]), .out(u_csamul_cska32_and17_7));
  fa fa_u_csamul_cska32_fa17_7_out(.a(u_csamul_cska32_and17_7[0]), .b(u_csamul_cska32_fa18_6_xor1[0]), .cin(u_csamul_cska32_fa17_6_or0[0]), .fa_xor1(u_csamul_cska32_fa17_7_xor1), .fa_or0(u_csamul_cska32_fa17_7_or0));
  and_gate and_gate_u_csamul_cska32_and18_7(.a(a[18]), .b(b[7]), .out(u_csamul_cska32_and18_7));
  fa fa_u_csamul_cska32_fa18_7_out(.a(u_csamul_cska32_and18_7[0]), .b(u_csamul_cska32_fa19_6_xor1[0]), .cin(u_csamul_cska32_fa18_6_or0[0]), .fa_xor1(u_csamul_cska32_fa18_7_xor1), .fa_or0(u_csamul_cska32_fa18_7_or0));
  and_gate and_gate_u_csamul_cska32_and19_7(.a(a[19]), .b(b[7]), .out(u_csamul_cska32_and19_7));
  fa fa_u_csamul_cska32_fa19_7_out(.a(u_csamul_cska32_and19_7[0]), .b(u_csamul_cska32_fa20_6_xor1[0]), .cin(u_csamul_cska32_fa19_6_or0[0]), .fa_xor1(u_csamul_cska32_fa19_7_xor1), .fa_or0(u_csamul_cska32_fa19_7_or0));
  and_gate and_gate_u_csamul_cska32_and20_7(.a(a[20]), .b(b[7]), .out(u_csamul_cska32_and20_7));
  fa fa_u_csamul_cska32_fa20_7_out(.a(u_csamul_cska32_and20_7[0]), .b(u_csamul_cska32_fa21_6_xor1[0]), .cin(u_csamul_cska32_fa20_6_or0[0]), .fa_xor1(u_csamul_cska32_fa20_7_xor1), .fa_or0(u_csamul_cska32_fa20_7_or0));
  and_gate and_gate_u_csamul_cska32_and21_7(.a(a[21]), .b(b[7]), .out(u_csamul_cska32_and21_7));
  fa fa_u_csamul_cska32_fa21_7_out(.a(u_csamul_cska32_and21_7[0]), .b(u_csamul_cska32_fa22_6_xor1[0]), .cin(u_csamul_cska32_fa21_6_or0[0]), .fa_xor1(u_csamul_cska32_fa21_7_xor1), .fa_or0(u_csamul_cska32_fa21_7_or0));
  and_gate and_gate_u_csamul_cska32_and22_7(.a(a[22]), .b(b[7]), .out(u_csamul_cska32_and22_7));
  fa fa_u_csamul_cska32_fa22_7_out(.a(u_csamul_cska32_and22_7[0]), .b(u_csamul_cska32_fa23_6_xor1[0]), .cin(u_csamul_cska32_fa22_6_or0[0]), .fa_xor1(u_csamul_cska32_fa22_7_xor1), .fa_or0(u_csamul_cska32_fa22_7_or0));
  and_gate and_gate_u_csamul_cska32_and23_7(.a(a[23]), .b(b[7]), .out(u_csamul_cska32_and23_7));
  fa fa_u_csamul_cska32_fa23_7_out(.a(u_csamul_cska32_and23_7[0]), .b(u_csamul_cska32_fa24_6_xor1[0]), .cin(u_csamul_cska32_fa23_6_or0[0]), .fa_xor1(u_csamul_cska32_fa23_7_xor1), .fa_or0(u_csamul_cska32_fa23_7_or0));
  and_gate and_gate_u_csamul_cska32_and24_7(.a(a[24]), .b(b[7]), .out(u_csamul_cska32_and24_7));
  fa fa_u_csamul_cska32_fa24_7_out(.a(u_csamul_cska32_and24_7[0]), .b(u_csamul_cska32_fa25_6_xor1[0]), .cin(u_csamul_cska32_fa24_6_or0[0]), .fa_xor1(u_csamul_cska32_fa24_7_xor1), .fa_or0(u_csamul_cska32_fa24_7_or0));
  and_gate and_gate_u_csamul_cska32_and25_7(.a(a[25]), .b(b[7]), .out(u_csamul_cska32_and25_7));
  fa fa_u_csamul_cska32_fa25_7_out(.a(u_csamul_cska32_and25_7[0]), .b(u_csamul_cska32_fa26_6_xor1[0]), .cin(u_csamul_cska32_fa25_6_or0[0]), .fa_xor1(u_csamul_cska32_fa25_7_xor1), .fa_or0(u_csamul_cska32_fa25_7_or0));
  and_gate and_gate_u_csamul_cska32_and26_7(.a(a[26]), .b(b[7]), .out(u_csamul_cska32_and26_7));
  fa fa_u_csamul_cska32_fa26_7_out(.a(u_csamul_cska32_and26_7[0]), .b(u_csamul_cska32_fa27_6_xor1[0]), .cin(u_csamul_cska32_fa26_6_or0[0]), .fa_xor1(u_csamul_cska32_fa26_7_xor1), .fa_or0(u_csamul_cska32_fa26_7_or0));
  and_gate and_gate_u_csamul_cska32_and27_7(.a(a[27]), .b(b[7]), .out(u_csamul_cska32_and27_7));
  fa fa_u_csamul_cska32_fa27_7_out(.a(u_csamul_cska32_and27_7[0]), .b(u_csamul_cska32_fa28_6_xor1[0]), .cin(u_csamul_cska32_fa27_6_or0[0]), .fa_xor1(u_csamul_cska32_fa27_7_xor1), .fa_or0(u_csamul_cska32_fa27_7_or0));
  and_gate and_gate_u_csamul_cska32_and28_7(.a(a[28]), .b(b[7]), .out(u_csamul_cska32_and28_7));
  fa fa_u_csamul_cska32_fa28_7_out(.a(u_csamul_cska32_and28_7[0]), .b(u_csamul_cska32_fa29_6_xor1[0]), .cin(u_csamul_cska32_fa28_6_or0[0]), .fa_xor1(u_csamul_cska32_fa28_7_xor1), .fa_or0(u_csamul_cska32_fa28_7_or0));
  and_gate and_gate_u_csamul_cska32_and29_7(.a(a[29]), .b(b[7]), .out(u_csamul_cska32_and29_7));
  fa fa_u_csamul_cska32_fa29_7_out(.a(u_csamul_cska32_and29_7[0]), .b(u_csamul_cska32_fa30_6_xor1[0]), .cin(u_csamul_cska32_fa29_6_or0[0]), .fa_xor1(u_csamul_cska32_fa29_7_xor1), .fa_or0(u_csamul_cska32_fa29_7_or0));
  and_gate and_gate_u_csamul_cska32_and30_7(.a(a[30]), .b(b[7]), .out(u_csamul_cska32_and30_7));
  fa fa_u_csamul_cska32_fa30_7_out(.a(u_csamul_cska32_and30_7[0]), .b(u_csamul_cska32_and31_6[0]), .cin(u_csamul_cska32_fa30_6_or0[0]), .fa_xor1(u_csamul_cska32_fa30_7_xor1), .fa_or0(u_csamul_cska32_fa30_7_or0));
  and_gate and_gate_u_csamul_cska32_and31_7(.a(a[31]), .b(b[7]), .out(u_csamul_cska32_and31_7));
  and_gate and_gate_u_csamul_cska32_and0_8(.a(a[0]), .b(b[8]), .out(u_csamul_cska32_and0_8));
  fa fa_u_csamul_cska32_fa0_8_out(.a(u_csamul_cska32_and0_8[0]), .b(u_csamul_cska32_fa1_7_xor1[0]), .cin(u_csamul_cska32_fa0_7_or0[0]), .fa_xor1(u_csamul_cska32_fa0_8_xor1), .fa_or0(u_csamul_cska32_fa0_8_or0));
  and_gate and_gate_u_csamul_cska32_and1_8(.a(a[1]), .b(b[8]), .out(u_csamul_cska32_and1_8));
  fa fa_u_csamul_cska32_fa1_8_out(.a(u_csamul_cska32_and1_8[0]), .b(u_csamul_cska32_fa2_7_xor1[0]), .cin(u_csamul_cska32_fa1_7_or0[0]), .fa_xor1(u_csamul_cska32_fa1_8_xor1), .fa_or0(u_csamul_cska32_fa1_8_or0));
  and_gate and_gate_u_csamul_cska32_and2_8(.a(a[2]), .b(b[8]), .out(u_csamul_cska32_and2_8));
  fa fa_u_csamul_cska32_fa2_8_out(.a(u_csamul_cska32_and2_8[0]), .b(u_csamul_cska32_fa3_7_xor1[0]), .cin(u_csamul_cska32_fa2_7_or0[0]), .fa_xor1(u_csamul_cska32_fa2_8_xor1), .fa_or0(u_csamul_cska32_fa2_8_or0));
  and_gate and_gate_u_csamul_cska32_and3_8(.a(a[3]), .b(b[8]), .out(u_csamul_cska32_and3_8));
  fa fa_u_csamul_cska32_fa3_8_out(.a(u_csamul_cska32_and3_8[0]), .b(u_csamul_cska32_fa4_7_xor1[0]), .cin(u_csamul_cska32_fa3_7_or0[0]), .fa_xor1(u_csamul_cska32_fa3_8_xor1), .fa_or0(u_csamul_cska32_fa3_8_or0));
  and_gate and_gate_u_csamul_cska32_and4_8(.a(a[4]), .b(b[8]), .out(u_csamul_cska32_and4_8));
  fa fa_u_csamul_cska32_fa4_8_out(.a(u_csamul_cska32_and4_8[0]), .b(u_csamul_cska32_fa5_7_xor1[0]), .cin(u_csamul_cska32_fa4_7_or0[0]), .fa_xor1(u_csamul_cska32_fa4_8_xor1), .fa_or0(u_csamul_cska32_fa4_8_or0));
  and_gate and_gate_u_csamul_cska32_and5_8(.a(a[5]), .b(b[8]), .out(u_csamul_cska32_and5_8));
  fa fa_u_csamul_cska32_fa5_8_out(.a(u_csamul_cska32_and5_8[0]), .b(u_csamul_cska32_fa6_7_xor1[0]), .cin(u_csamul_cska32_fa5_7_or0[0]), .fa_xor1(u_csamul_cska32_fa5_8_xor1), .fa_or0(u_csamul_cska32_fa5_8_or0));
  and_gate and_gate_u_csamul_cska32_and6_8(.a(a[6]), .b(b[8]), .out(u_csamul_cska32_and6_8));
  fa fa_u_csamul_cska32_fa6_8_out(.a(u_csamul_cska32_and6_8[0]), .b(u_csamul_cska32_fa7_7_xor1[0]), .cin(u_csamul_cska32_fa6_7_or0[0]), .fa_xor1(u_csamul_cska32_fa6_8_xor1), .fa_or0(u_csamul_cska32_fa6_8_or0));
  and_gate and_gate_u_csamul_cska32_and7_8(.a(a[7]), .b(b[8]), .out(u_csamul_cska32_and7_8));
  fa fa_u_csamul_cska32_fa7_8_out(.a(u_csamul_cska32_and7_8[0]), .b(u_csamul_cska32_fa8_7_xor1[0]), .cin(u_csamul_cska32_fa7_7_or0[0]), .fa_xor1(u_csamul_cska32_fa7_8_xor1), .fa_or0(u_csamul_cska32_fa7_8_or0));
  and_gate and_gate_u_csamul_cska32_and8_8(.a(a[8]), .b(b[8]), .out(u_csamul_cska32_and8_8));
  fa fa_u_csamul_cska32_fa8_8_out(.a(u_csamul_cska32_and8_8[0]), .b(u_csamul_cska32_fa9_7_xor1[0]), .cin(u_csamul_cska32_fa8_7_or0[0]), .fa_xor1(u_csamul_cska32_fa8_8_xor1), .fa_or0(u_csamul_cska32_fa8_8_or0));
  and_gate and_gate_u_csamul_cska32_and9_8(.a(a[9]), .b(b[8]), .out(u_csamul_cska32_and9_8));
  fa fa_u_csamul_cska32_fa9_8_out(.a(u_csamul_cska32_and9_8[0]), .b(u_csamul_cska32_fa10_7_xor1[0]), .cin(u_csamul_cska32_fa9_7_or0[0]), .fa_xor1(u_csamul_cska32_fa9_8_xor1), .fa_or0(u_csamul_cska32_fa9_8_or0));
  and_gate and_gate_u_csamul_cska32_and10_8(.a(a[10]), .b(b[8]), .out(u_csamul_cska32_and10_8));
  fa fa_u_csamul_cska32_fa10_8_out(.a(u_csamul_cska32_and10_8[0]), .b(u_csamul_cska32_fa11_7_xor1[0]), .cin(u_csamul_cska32_fa10_7_or0[0]), .fa_xor1(u_csamul_cska32_fa10_8_xor1), .fa_or0(u_csamul_cska32_fa10_8_or0));
  and_gate and_gate_u_csamul_cska32_and11_8(.a(a[11]), .b(b[8]), .out(u_csamul_cska32_and11_8));
  fa fa_u_csamul_cska32_fa11_8_out(.a(u_csamul_cska32_and11_8[0]), .b(u_csamul_cska32_fa12_7_xor1[0]), .cin(u_csamul_cska32_fa11_7_or0[0]), .fa_xor1(u_csamul_cska32_fa11_8_xor1), .fa_or0(u_csamul_cska32_fa11_8_or0));
  and_gate and_gate_u_csamul_cska32_and12_8(.a(a[12]), .b(b[8]), .out(u_csamul_cska32_and12_8));
  fa fa_u_csamul_cska32_fa12_8_out(.a(u_csamul_cska32_and12_8[0]), .b(u_csamul_cska32_fa13_7_xor1[0]), .cin(u_csamul_cska32_fa12_7_or0[0]), .fa_xor1(u_csamul_cska32_fa12_8_xor1), .fa_or0(u_csamul_cska32_fa12_8_or0));
  and_gate and_gate_u_csamul_cska32_and13_8(.a(a[13]), .b(b[8]), .out(u_csamul_cska32_and13_8));
  fa fa_u_csamul_cska32_fa13_8_out(.a(u_csamul_cska32_and13_8[0]), .b(u_csamul_cska32_fa14_7_xor1[0]), .cin(u_csamul_cska32_fa13_7_or0[0]), .fa_xor1(u_csamul_cska32_fa13_8_xor1), .fa_or0(u_csamul_cska32_fa13_8_or0));
  and_gate and_gate_u_csamul_cska32_and14_8(.a(a[14]), .b(b[8]), .out(u_csamul_cska32_and14_8));
  fa fa_u_csamul_cska32_fa14_8_out(.a(u_csamul_cska32_and14_8[0]), .b(u_csamul_cska32_fa15_7_xor1[0]), .cin(u_csamul_cska32_fa14_7_or0[0]), .fa_xor1(u_csamul_cska32_fa14_8_xor1), .fa_or0(u_csamul_cska32_fa14_8_or0));
  and_gate and_gate_u_csamul_cska32_and15_8(.a(a[15]), .b(b[8]), .out(u_csamul_cska32_and15_8));
  fa fa_u_csamul_cska32_fa15_8_out(.a(u_csamul_cska32_and15_8[0]), .b(u_csamul_cska32_fa16_7_xor1[0]), .cin(u_csamul_cska32_fa15_7_or0[0]), .fa_xor1(u_csamul_cska32_fa15_8_xor1), .fa_or0(u_csamul_cska32_fa15_8_or0));
  and_gate and_gate_u_csamul_cska32_and16_8(.a(a[16]), .b(b[8]), .out(u_csamul_cska32_and16_8));
  fa fa_u_csamul_cska32_fa16_8_out(.a(u_csamul_cska32_and16_8[0]), .b(u_csamul_cska32_fa17_7_xor1[0]), .cin(u_csamul_cska32_fa16_7_or0[0]), .fa_xor1(u_csamul_cska32_fa16_8_xor1), .fa_or0(u_csamul_cska32_fa16_8_or0));
  and_gate and_gate_u_csamul_cska32_and17_8(.a(a[17]), .b(b[8]), .out(u_csamul_cska32_and17_8));
  fa fa_u_csamul_cska32_fa17_8_out(.a(u_csamul_cska32_and17_8[0]), .b(u_csamul_cska32_fa18_7_xor1[0]), .cin(u_csamul_cska32_fa17_7_or0[0]), .fa_xor1(u_csamul_cska32_fa17_8_xor1), .fa_or0(u_csamul_cska32_fa17_8_or0));
  and_gate and_gate_u_csamul_cska32_and18_8(.a(a[18]), .b(b[8]), .out(u_csamul_cska32_and18_8));
  fa fa_u_csamul_cska32_fa18_8_out(.a(u_csamul_cska32_and18_8[0]), .b(u_csamul_cska32_fa19_7_xor1[0]), .cin(u_csamul_cska32_fa18_7_or0[0]), .fa_xor1(u_csamul_cska32_fa18_8_xor1), .fa_or0(u_csamul_cska32_fa18_8_or0));
  and_gate and_gate_u_csamul_cska32_and19_8(.a(a[19]), .b(b[8]), .out(u_csamul_cska32_and19_8));
  fa fa_u_csamul_cska32_fa19_8_out(.a(u_csamul_cska32_and19_8[0]), .b(u_csamul_cska32_fa20_7_xor1[0]), .cin(u_csamul_cska32_fa19_7_or0[0]), .fa_xor1(u_csamul_cska32_fa19_8_xor1), .fa_or0(u_csamul_cska32_fa19_8_or0));
  and_gate and_gate_u_csamul_cska32_and20_8(.a(a[20]), .b(b[8]), .out(u_csamul_cska32_and20_8));
  fa fa_u_csamul_cska32_fa20_8_out(.a(u_csamul_cska32_and20_8[0]), .b(u_csamul_cska32_fa21_7_xor1[0]), .cin(u_csamul_cska32_fa20_7_or0[0]), .fa_xor1(u_csamul_cska32_fa20_8_xor1), .fa_or0(u_csamul_cska32_fa20_8_or0));
  and_gate and_gate_u_csamul_cska32_and21_8(.a(a[21]), .b(b[8]), .out(u_csamul_cska32_and21_8));
  fa fa_u_csamul_cska32_fa21_8_out(.a(u_csamul_cska32_and21_8[0]), .b(u_csamul_cska32_fa22_7_xor1[0]), .cin(u_csamul_cska32_fa21_7_or0[0]), .fa_xor1(u_csamul_cska32_fa21_8_xor1), .fa_or0(u_csamul_cska32_fa21_8_or0));
  and_gate and_gate_u_csamul_cska32_and22_8(.a(a[22]), .b(b[8]), .out(u_csamul_cska32_and22_8));
  fa fa_u_csamul_cska32_fa22_8_out(.a(u_csamul_cska32_and22_8[0]), .b(u_csamul_cska32_fa23_7_xor1[0]), .cin(u_csamul_cska32_fa22_7_or0[0]), .fa_xor1(u_csamul_cska32_fa22_8_xor1), .fa_or0(u_csamul_cska32_fa22_8_or0));
  and_gate and_gate_u_csamul_cska32_and23_8(.a(a[23]), .b(b[8]), .out(u_csamul_cska32_and23_8));
  fa fa_u_csamul_cska32_fa23_8_out(.a(u_csamul_cska32_and23_8[0]), .b(u_csamul_cska32_fa24_7_xor1[0]), .cin(u_csamul_cska32_fa23_7_or0[0]), .fa_xor1(u_csamul_cska32_fa23_8_xor1), .fa_or0(u_csamul_cska32_fa23_8_or0));
  and_gate and_gate_u_csamul_cska32_and24_8(.a(a[24]), .b(b[8]), .out(u_csamul_cska32_and24_8));
  fa fa_u_csamul_cska32_fa24_8_out(.a(u_csamul_cska32_and24_8[0]), .b(u_csamul_cska32_fa25_7_xor1[0]), .cin(u_csamul_cska32_fa24_7_or0[0]), .fa_xor1(u_csamul_cska32_fa24_8_xor1), .fa_or0(u_csamul_cska32_fa24_8_or0));
  and_gate and_gate_u_csamul_cska32_and25_8(.a(a[25]), .b(b[8]), .out(u_csamul_cska32_and25_8));
  fa fa_u_csamul_cska32_fa25_8_out(.a(u_csamul_cska32_and25_8[0]), .b(u_csamul_cska32_fa26_7_xor1[0]), .cin(u_csamul_cska32_fa25_7_or0[0]), .fa_xor1(u_csamul_cska32_fa25_8_xor1), .fa_or0(u_csamul_cska32_fa25_8_or0));
  and_gate and_gate_u_csamul_cska32_and26_8(.a(a[26]), .b(b[8]), .out(u_csamul_cska32_and26_8));
  fa fa_u_csamul_cska32_fa26_8_out(.a(u_csamul_cska32_and26_8[0]), .b(u_csamul_cska32_fa27_7_xor1[0]), .cin(u_csamul_cska32_fa26_7_or0[0]), .fa_xor1(u_csamul_cska32_fa26_8_xor1), .fa_or0(u_csamul_cska32_fa26_8_or0));
  and_gate and_gate_u_csamul_cska32_and27_8(.a(a[27]), .b(b[8]), .out(u_csamul_cska32_and27_8));
  fa fa_u_csamul_cska32_fa27_8_out(.a(u_csamul_cska32_and27_8[0]), .b(u_csamul_cska32_fa28_7_xor1[0]), .cin(u_csamul_cska32_fa27_7_or0[0]), .fa_xor1(u_csamul_cska32_fa27_8_xor1), .fa_or0(u_csamul_cska32_fa27_8_or0));
  and_gate and_gate_u_csamul_cska32_and28_8(.a(a[28]), .b(b[8]), .out(u_csamul_cska32_and28_8));
  fa fa_u_csamul_cska32_fa28_8_out(.a(u_csamul_cska32_and28_8[0]), .b(u_csamul_cska32_fa29_7_xor1[0]), .cin(u_csamul_cska32_fa28_7_or0[0]), .fa_xor1(u_csamul_cska32_fa28_8_xor1), .fa_or0(u_csamul_cska32_fa28_8_or0));
  and_gate and_gate_u_csamul_cska32_and29_8(.a(a[29]), .b(b[8]), .out(u_csamul_cska32_and29_8));
  fa fa_u_csamul_cska32_fa29_8_out(.a(u_csamul_cska32_and29_8[0]), .b(u_csamul_cska32_fa30_7_xor1[0]), .cin(u_csamul_cska32_fa29_7_or0[0]), .fa_xor1(u_csamul_cska32_fa29_8_xor1), .fa_or0(u_csamul_cska32_fa29_8_or0));
  and_gate and_gate_u_csamul_cska32_and30_8(.a(a[30]), .b(b[8]), .out(u_csamul_cska32_and30_8));
  fa fa_u_csamul_cska32_fa30_8_out(.a(u_csamul_cska32_and30_8[0]), .b(u_csamul_cska32_and31_7[0]), .cin(u_csamul_cska32_fa30_7_or0[0]), .fa_xor1(u_csamul_cska32_fa30_8_xor1), .fa_or0(u_csamul_cska32_fa30_8_or0));
  and_gate and_gate_u_csamul_cska32_and31_8(.a(a[31]), .b(b[8]), .out(u_csamul_cska32_and31_8));
  and_gate and_gate_u_csamul_cska32_and0_9(.a(a[0]), .b(b[9]), .out(u_csamul_cska32_and0_9));
  fa fa_u_csamul_cska32_fa0_9_out(.a(u_csamul_cska32_and0_9[0]), .b(u_csamul_cska32_fa1_8_xor1[0]), .cin(u_csamul_cska32_fa0_8_or0[0]), .fa_xor1(u_csamul_cska32_fa0_9_xor1), .fa_or0(u_csamul_cska32_fa0_9_or0));
  and_gate and_gate_u_csamul_cska32_and1_9(.a(a[1]), .b(b[9]), .out(u_csamul_cska32_and1_9));
  fa fa_u_csamul_cska32_fa1_9_out(.a(u_csamul_cska32_and1_9[0]), .b(u_csamul_cska32_fa2_8_xor1[0]), .cin(u_csamul_cska32_fa1_8_or0[0]), .fa_xor1(u_csamul_cska32_fa1_9_xor1), .fa_or0(u_csamul_cska32_fa1_9_or0));
  and_gate and_gate_u_csamul_cska32_and2_9(.a(a[2]), .b(b[9]), .out(u_csamul_cska32_and2_9));
  fa fa_u_csamul_cska32_fa2_9_out(.a(u_csamul_cska32_and2_9[0]), .b(u_csamul_cska32_fa3_8_xor1[0]), .cin(u_csamul_cska32_fa2_8_or0[0]), .fa_xor1(u_csamul_cska32_fa2_9_xor1), .fa_or0(u_csamul_cska32_fa2_9_or0));
  and_gate and_gate_u_csamul_cska32_and3_9(.a(a[3]), .b(b[9]), .out(u_csamul_cska32_and3_9));
  fa fa_u_csamul_cska32_fa3_9_out(.a(u_csamul_cska32_and3_9[0]), .b(u_csamul_cska32_fa4_8_xor1[0]), .cin(u_csamul_cska32_fa3_8_or0[0]), .fa_xor1(u_csamul_cska32_fa3_9_xor1), .fa_or0(u_csamul_cska32_fa3_9_or0));
  and_gate and_gate_u_csamul_cska32_and4_9(.a(a[4]), .b(b[9]), .out(u_csamul_cska32_and4_9));
  fa fa_u_csamul_cska32_fa4_9_out(.a(u_csamul_cska32_and4_9[0]), .b(u_csamul_cska32_fa5_8_xor1[0]), .cin(u_csamul_cska32_fa4_8_or0[0]), .fa_xor1(u_csamul_cska32_fa4_9_xor1), .fa_or0(u_csamul_cska32_fa4_9_or0));
  and_gate and_gate_u_csamul_cska32_and5_9(.a(a[5]), .b(b[9]), .out(u_csamul_cska32_and5_9));
  fa fa_u_csamul_cska32_fa5_9_out(.a(u_csamul_cska32_and5_9[0]), .b(u_csamul_cska32_fa6_8_xor1[0]), .cin(u_csamul_cska32_fa5_8_or0[0]), .fa_xor1(u_csamul_cska32_fa5_9_xor1), .fa_or0(u_csamul_cska32_fa5_9_or0));
  and_gate and_gate_u_csamul_cska32_and6_9(.a(a[6]), .b(b[9]), .out(u_csamul_cska32_and6_9));
  fa fa_u_csamul_cska32_fa6_9_out(.a(u_csamul_cska32_and6_9[0]), .b(u_csamul_cska32_fa7_8_xor1[0]), .cin(u_csamul_cska32_fa6_8_or0[0]), .fa_xor1(u_csamul_cska32_fa6_9_xor1), .fa_or0(u_csamul_cska32_fa6_9_or0));
  and_gate and_gate_u_csamul_cska32_and7_9(.a(a[7]), .b(b[9]), .out(u_csamul_cska32_and7_9));
  fa fa_u_csamul_cska32_fa7_9_out(.a(u_csamul_cska32_and7_9[0]), .b(u_csamul_cska32_fa8_8_xor1[0]), .cin(u_csamul_cska32_fa7_8_or0[0]), .fa_xor1(u_csamul_cska32_fa7_9_xor1), .fa_or0(u_csamul_cska32_fa7_9_or0));
  and_gate and_gate_u_csamul_cska32_and8_9(.a(a[8]), .b(b[9]), .out(u_csamul_cska32_and8_9));
  fa fa_u_csamul_cska32_fa8_9_out(.a(u_csamul_cska32_and8_9[0]), .b(u_csamul_cska32_fa9_8_xor1[0]), .cin(u_csamul_cska32_fa8_8_or0[0]), .fa_xor1(u_csamul_cska32_fa8_9_xor1), .fa_or0(u_csamul_cska32_fa8_9_or0));
  and_gate and_gate_u_csamul_cska32_and9_9(.a(a[9]), .b(b[9]), .out(u_csamul_cska32_and9_9));
  fa fa_u_csamul_cska32_fa9_9_out(.a(u_csamul_cska32_and9_9[0]), .b(u_csamul_cska32_fa10_8_xor1[0]), .cin(u_csamul_cska32_fa9_8_or0[0]), .fa_xor1(u_csamul_cska32_fa9_9_xor1), .fa_or0(u_csamul_cska32_fa9_9_or0));
  and_gate and_gate_u_csamul_cska32_and10_9(.a(a[10]), .b(b[9]), .out(u_csamul_cska32_and10_9));
  fa fa_u_csamul_cska32_fa10_9_out(.a(u_csamul_cska32_and10_9[0]), .b(u_csamul_cska32_fa11_8_xor1[0]), .cin(u_csamul_cska32_fa10_8_or0[0]), .fa_xor1(u_csamul_cska32_fa10_9_xor1), .fa_or0(u_csamul_cska32_fa10_9_or0));
  and_gate and_gate_u_csamul_cska32_and11_9(.a(a[11]), .b(b[9]), .out(u_csamul_cska32_and11_9));
  fa fa_u_csamul_cska32_fa11_9_out(.a(u_csamul_cska32_and11_9[0]), .b(u_csamul_cska32_fa12_8_xor1[0]), .cin(u_csamul_cska32_fa11_8_or0[0]), .fa_xor1(u_csamul_cska32_fa11_9_xor1), .fa_or0(u_csamul_cska32_fa11_9_or0));
  and_gate and_gate_u_csamul_cska32_and12_9(.a(a[12]), .b(b[9]), .out(u_csamul_cska32_and12_9));
  fa fa_u_csamul_cska32_fa12_9_out(.a(u_csamul_cska32_and12_9[0]), .b(u_csamul_cska32_fa13_8_xor1[0]), .cin(u_csamul_cska32_fa12_8_or0[0]), .fa_xor1(u_csamul_cska32_fa12_9_xor1), .fa_or0(u_csamul_cska32_fa12_9_or0));
  and_gate and_gate_u_csamul_cska32_and13_9(.a(a[13]), .b(b[9]), .out(u_csamul_cska32_and13_9));
  fa fa_u_csamul_cska32_fa13_9_out(.a(u_csamul_cska32_and13_9[0]), .b(u_csamul_cska32_fa14_8_xor1[0]), .cin(u_csamul_cska32_fa13_8_or0[0]), .fa_xor1(u_csamul_cska32_fa13_9_xor1), .fa_or0(u_csamul_cska32_fa13_9_or0));
  and_gate and_gate_u_csamul_cska32_and14_9(.a(a[14]), .b(b[9]), .out(u_csamul_cska32_and14_9));
  fa fa_u_csamul_cska32_fa14_9_out(.a(u_csamul_cska32_and14_9[0]), .b(u_csamul_cska32_fa15_8_xor1[0]), .cin(u_csamul_cska32_fa14_8_or0[0]), .fa_xor1(u_csamul_cska32_fa14_9_xor1), .fa_or0(u_csamul_cska32_fa14_9_or0));
  and_gate and_gate_u_csamul_cska32_and15_9(.a(a[15]), .b(b[9]), .out(u_csamul_cska32_and15_9));
  fa fa_u_csamul_cska32_fa15_9_out(.a(u_csamul_cska32_and15_9[0]), .b(u_csamul_cska32_fa16_8_xor1[0]), .cin(u_csamul_cska32_fa15_8_or0[0]), .fa_xor1(u_csamul_cska32_fa15_9_xor1), .fa_or0(u_csamul_cska32_fa15_9_or0));
  and_gate and_gate_u_csamul_cska32_and16_9(.a(a[16]), .b(b[9]), .out(u_csamul_cska32_and16_9));
  fa fa_u_csamul_cska32_fa16_9_out(.a(u_csamul_cska32_and16_9[0]), .b(u_csamul_cska32_fa17_8_xor1[0]), .cin(u_csamul_cska32_fa16_8_or0[0]), .fa_xor1(u_csamul_cska32_fa16_9_xor1), .fa_or0(u_csamul_cska32_fa16_9_or0));
  and_gate and_gate_u_csamul_cska32_and17_9(.a(a[17]), .b(b[9]), .out(u_csamul_cska32_and17_9));
  fa fa_u_csamul_cska32_fa17_9_out(.a(u_csamul_cska32_and17_9[0]), .b(u_csamul_cska32_fa18_8_xor1[0]), .cin(u_csamul_cska32_fa17_8_or0[0]), .fa_xor1(u_csamul_cska32_fa17_9_xor1), .fa_or0(u_csamul_cska32_fa17_9_or0));
  and_gate and_gate_u_csamul_cska32_and18_9(.a(a[18]), .b(b[9]), .out(u_csamul_cska32_and18_9));
  fa fa_u_csamul_cska32_fa18_9_out(.a(u_csamul_cska32_and18_9[0]), .b(u_csamul_cska32_fa19_8_xor1[0]), .cin(u_csamul_cska32_fa18_8_or0[0]), .fa_xor1(u_csamul_cska32_fa18_9_xor1), .fa_or0(u_csamul_cska32_fa18_9_or0));
  and_gate and_gate_u_csamul_cska32_and19_9(.a(a[19]), .b(b[9]), .out(u_csamul_cska32_and19_9));
  fa fa_u_csamul_cska32_fa19_9_out(.a(u_csamul_cska32_and19_9[0]), .b(u_csamul_cska32_fa20_8_xor1[0]), .cin(u_csamul_cska32_fa19_8_or0[0]), .fa_xor1(u_csamul_cska32_fa19_9_xor1), .fa_or0(u_csamul_cska32_fa19_9_or0));
  and_gate and_gate_u_csamul_cska32_and20_9(.a(a[20]), .b(b[9]), .out(u_csamul_cska32_and20_9));
  fa fa_u_csamul_cska32_fa20_9_out(.a(u_csamul_cska32_and20_9[0]), .b(u_csamul_cska32_fa21_8_xor1[0]), .cin(u_csamul_cska32_fa20_8_or0[0]), .fa_xor1(u_csamul_cska32_fa20_9_xor1), .fa_or0(u_csamul_cska32_fa20_9_or0));
  and_gate and_gate_u_csamul_cska32_and21_9(.a(a[21]), .b(b[9]), .out(u_csamul_cska32_and21_9));
  fa fa_u_csamul_cska32_fa21_9_out(.a(u_csamul_cska32_and21_9[0]), .b(u_csamul_cska32_fa22_8_xor1[0]), .cin(u_csamul_cska32_fa21_8_or0[0]), .fa_xor1(u_csamul_cska32_fa21_9_xor1), .fa_or0(u_csamul_cska32_fa21_9_or0));
  and_gate and_gate_u_csamul_cska32_and22_9(.a(a[22]), .b(b[9]), .out(u_csamul_cska32_and22_9));
  fa fa_u_csamul_cska32_fa22_9_out(.a(u_csamul_cska32_and22_9[0]), .b(u_csamul_cska32_fa23_8_xor1[0]), .cin(u_csamul_cska32_fa22_8_or0[0]), .fa_xor1(u_csamul_cska32_fa22_9_xor1), .fa_or0(u_csamul_cska32_fa22_9_or0));
  and_gate and_gate_u_csamul_cska32_and23_9(.a(a[23]), .b(b[9]), .out(u_csamul_cska32_and23_9));
  fa fa_u_csamul_cska32_fa23_9_out(.a(u_csamul_cska32_and23_9[0]), .b(u_csamul_cska32_fa24_8_xor1[0]), .cin(u_csamul_cska32_fa23_8_or0[0]), .fa_xor1(u_csamul_cska32_fa23_9_xor1), .fa_or0(u_csamul_cska32_fa23_9_or0));
  and_gate and_gate_u_csamul_cska32_and24_9(.a(a[24]), .b(b[9]), .out(u_csamul_cska32_and24_9));
  fa fa_u_csamul_cska32_fa24_9_out(.a(u_csamul_cska32_and24_9[0]), .b(u_csamul_cska32_fa25_8_xor1[0]), .cin(u_csamul_cska32_fa24_8_or0[0]), .fa_xor1(u_csamul_cska32_fa24_9_xor1), .fa_or0(u_csamul_cska32_fa24_9_or0));
  and_gate and_gate_u_csamul_cska32_and25_9(.a(a[25]), .b(b[9]), .out(u_csamul_cska32_and25_9));
  fa fa_u_csamul_cska32_fa25_9_out(.a(u_csamul_cska32_and25_9[0]), .b(u_csamul_cska32_fa26_8_xor1[0]), .cin(u_csamul_cska32_fa25_8_or0[0]), .fa_xor1(u_csamul_cska32_fa25_9_xor1), .fa_or0(u_csamul_cska32_fa25_9_or0));
  and_gate and_gate_u_csamul_cska32_and26_9(.a(a[26]), .b(b[9]), .out(u_csamul_cska32_and26_9));
  fa fa_u_csamul_cska32_fa26_9_out(.a(u_csamul_cska32_and26_9[0]), .b(u_csamul_cska32_fa27_8_xor1[0]), .cin(u_csamul_cska32_fa26_8_or0[0]), .fa_xor1(u_csamul_cska32_fa26_9_xor1), .fa_or0(u_csamul_cska32_fa26_9_or0));
  and_gate and_gate_u_csamul_cska32_and27_9(.a(a[27]), .b(b[9]), .out(u_csamul_cska32_and27_9));
  fa fa_u_csamul_cska32_fa27_9_out(.a(u_csamul_cska32_and27_9[0]), .b(u_csamul_cska32_fa28_8_xor1[0]), .cin(u_csamul_cska32_fa27_8_or0[0]), .fa_xor1(u_csamul_cska32_fa27_9_xor1), .fa_or0(u_csamul_cska32_fa27_9_or0));
  and_gate and_gate_u_csamul_cska32_and28_9(.a(a[28]), .b(b[9]), .out(u_csamul_cska32_and28_9));
  fa fa_u_csamul_cska32_fa28_9_out(.a(u_csamul_cska32_and28_9[0]), .b(u_csamul_cska32_fa29_8_xor1[0]), .cin(u_csamul_cska32_fa28_8_or0[0]), .fa_xor1(u_csamul_cska32_fa28_9_xor1), .fa_or0(u_csamul_cska32_fa28_9_or0));
  and_gate and_gate_u_csamul_cska32_and29_9(.a(a[29]), .b(b[9]), .out(u_csamul_cska32_and29_9));
  fa fa_u_csamul_cska32_fa29_9_out(.a(u_csamul_cska32_and29_9[0]), .b(u_csamul_cska32_fa30_8_xor1[0]), .cin(u_csamul_cska32_fa29_8_or0[0]), .fa_xor1(u_csamul_cska32_fa29_9_xor1), .fa_or0(u_csamul_cska32_fa29_9_or0));
  and_gate and_gate_u_csamul_cska32_and30_9(.a(a[30]), .b(b[9]), .out(u_csamul_cska32_and30_9));
  fa fa_u_csamul_cska32_fa30_9_out(.a(u_csamul_cska32_and30_9[0]), .b(u_csamul_cska32_and31_8[0]), .cin(u_csamul_cska32_fa30_8_or0[0]), .fa_xor1(u_csamul_cska32_fa30_9_xor1), .fa_or0(u_csamul_cska32_fa30_9_or0));
  and_gate and_gate_u_csamul_cska32_and31_9(.a(a[31]), .b(b[9]), .out(u_csamul_cska32_and31_9));
  and_gate and_gate_u_csamul_cska32_and0_10(.a(a[0]), .b(b[10]), .out(u_csamul_cska32_and0_10));
  fa fa_u_csamul_cska32_fa0_10_out(.a(u_csamul_cska32_and0_10[0]), .b(u_csamul_cska32_fa1_9_xor1[0]), .cin(u_csamul_cska32_fa0_9_or0[0]), .fa_xor1(u_csamul_cska32_fa0_10_xor1), .fa_or0(u_csamul_cska32_fa0_10_or0));
  and_gate and_gate_u_csamul_cska32_and1_10(.a(a[1]), .b(b[10]), .out(u_csamul_cska32_and1_10));
  fa fa_u_csamul_cska32_fa1_10_out(.a(u_csamul_cska32_and1_10[0]), .b(u_csamul_cska32_fa2_9_xor1[0]), .cin(u_csamul_cska32_fa1_9_or0[0]), .fa_xor1(u_csamul_cska32_fa1_10_xor1), .fa_or0(u_csamul_cska32_fa1_10_or0));
  and_gate and_gate_u_csamul_cska32_and2_10(.a(a[2]), .b(b[10]), .out(u_csamul_cska32_and2_10));
  fa fa_u_csamul_cska32_fa2_10_out(.a(u_csamul_cska32_and2_10[0]), .b(u_csamul_cska32_fa3_9_xor1[0]), .cin(u_csamul_cska32_fa2_9_or0[0]), .fa_xor1(u_csamul_cska32_fa2_10_xor1), .fa_or0(u_csamul_cska32_fa2_10_or0));
  and_gate and_gate_u_csamul_cska32_and3_10(.a(a[3]), .b(b[10]), .out(u_csamul_cska32_and3_10));
  fa fa_u_csamul_cska32_fa3_10_out(.a(u_csamul_cska32_and3_10[0]), .b(u_csamul_cska32_fa4_9_xor1[0]), .cin(u_csamul_cska32_fa3_9_or0[0]), .fa_xor1(u_csamul_cska32_fa3_10_xor1), .fa_or0(u_csamul_cska32_fa3_10_or0));
  and_gate and_gate_u_csamul_cska32_and4_10(.a(a[4]), .b(b[10]), .out(u_csamul_cska32_and4_10));
  fa fa_u_csamul_cska32_fa4_10_out(.a(u_csamul_cska32_and4_10[0]), .b(u_csamul_cska32_fa5_9_xor1[0]), .cin(u_csamul_cska32_fa4_9_or0[0]), .fa_xor1(u_csamul_cska32_fa4_10_xor1), .fa_or0(u_csamul_cska32_fa4_10_or0));
  and_gate and_gate_u_csamul_cska32_and5_10(.a(a[5]), .b(b[10]), .out(u_csamul_cska32_and5_10));
  fa fa_u_csamul_cska32_fa5_10_out(.a(u_csamul_cska32_and5_10[0]), .b(u_csamul_cska32_fa6_9_xor1[0]), .cin(u_csamul_cska32_fa5_9_or0[0]), .fa_xor1(u_csamul_cska32_fa5_10_xor1), .fa_or0(u_csamul_cska32_fa5_10_or0));
  and_gate and_gate_u_csamul_cska32_and6_10(.a(a[6]), .b(b[10]), .out(u_csamul_cska32_and6_10));
  fa fa_u_csamul_cska32_fa6_10_out(.a(u_csamul_cska32_and6_10[0]), .b(u_csamul_cska32_fa7_9_xor1[0]), .cin(u_csamul_cska32_fa6_9_or0[0]), .fa_xor1(u_csamul_cska32_fa6_10_xor1), .fa_or0(u_csamul_cska32_fa6_10_or0));
  and_gate and_gate_u_csamul_cska32_and7_10(.a(a[7]), .b(b[10]), .out(u_csamul_cska32_and7_10));
  fa fa_u_csamul_cska32_fa7_10_out(.a(u_csamul_cska32_and7_10[0]), .b(u_csamul_cska32_fa8_9_xor1[0]), .cin(u_csamul_cska32_fa7_9_or0[0]), .fa_xor1(u_csamul_cska32_fa7_10_xor1), .fa_or0(u_csamul_cska32_fa7_10_or0));
  and_gate and_gate_u_csamul_cska32_and8_10(.a(a[8]), .b(b[10]), .out(u_csamul_cska32_and8_10));
  fa fa_u_csamul_cska32_fa8_10_out(.a(u_csamul_cska32_and8_10[0]), .b(u_csamul_cska32_fa9_9_xor1[0]), .cin(u_csamul_cska32_fa8_9_or0[0]), .fa_xor1(u_csamul_cska32_fa8_10_xor1), .fa_or0(u_csamul_cska32_fa8_10_or0));
  and_gate and_gate_u_csamul_cska32_and9_10(.a(a[9]), .b(b[10]), .out(u_csamul_cska32_and9_10));
  fa fa_u_csamul_cska32_fa9_10_out(.a(u_csamul_cska32_and9_10[0]), .b(u_csamul_cska32_fa10_9_xor1[0]), .cin(u_csamul_cska32_fa9_9_or0[0]), .fa_xor1(u_csamul_cska32_fa9_10_xor1), .fa_or0(u_csamul_cska32_fa9_10_or0));
  and_gate and_gate_u_csamul_cska32_and10_10(.a(a[10]), .b(b[10]), .out(u_csamul_cska32_and10_10));
  fa fa_u_csamul_cska32_fa10_10_out(.a(u_csamul_cska32_and10_10[0]), .b(u_csamul_cska32_fa11_9_xor1[0]), .cin(u_csamul_cska32_fa10_9_or0[0]), .fa_xor1(u_csamul_cska32_fa10_10_xor1), .fa_or0(u_csamul_cska32_fa10_10_or0));
  and_gate and_gate_u_csamul_cska32_and11_10(.a(a[11]), .b(b[10]), .out(u_csamul_cska32_and11_10));
  fa fa_u_csamul_cska32_fa11_10_out(.a(u_csamul_cska32_and11_10[0]), .b(u_csamul_cska32_fa12_9_xor1[0]), .cin(u_csamul_cska32_fa11_9_or0[0]), .fa_xor1(u_csamul_cska32_fa11_10_xor1), .fa_or0(u_csamul_cska32_fa11_10_or0));
  and_gate and_gate_u_csamul_cska32_and12_10(.a(a[12]), .b(b[10]), .out(u_csamul_cska32_and12_10));
  fa fa_u_csamul_cska32_fa12_10_out(.a(u_csamul_cska32_and12_10[0]), .b(u_csamul_cska32_fa13_9_xor1[0]), .cin(u_csamul_cska32_fa12_9_or0[0]), .fa_xor1(u_csamul_cska32_fa12_10_xor1), .fa_or0(u_csamul_cska32_fa12_10_or0));
  and_gate and_gate_u_csamul_cska32_and13_10(.a(a[13]), .b(b[10]), .out(u_csamul_cska32_and13_10));
  fa fa_u_csamul_cska32_fa13_10_out(.a(u_csamul_cska32_and13_10[0]), .b(u_csamul_cska32_fa14_9_xor1[0]), .cin(u_csamul_cska32_fa13_9_or0[0]), .fa_xor1(u_csamul_cska32_fa13_10_xor1), .fa_or0(u_csamul_cska32_fa13_10_or0));
  and_gate and_gate_u_csamul_cska32_and14_10(.a(a[14]), .b(b[10]), .out(u_csamul_cska32_and14_10));
  fa fa_u_csamul_cska32_fa14_10_out(.a(u_csamul_cska32_and14_10[0]), .b(u_csamul_cska32_fa15_9_xor1[0]), .cin(u_csamul_cska32_fa14_9_or0[0]), .fa_xor1(u_csamul_cska32_fa14_10_xor1), .fa_or0(u_csamul_cska32_fa14_10_or0));
  and_gate and_gate_u_csamul_cska32_and15_10(.a(a[15]), .b(b[10]), .out(u_csamul_cska32_and15_10));
  fa fa_u_csamul_cska32_fa15_10_out(.a(u_csamul_cska32_and15_10[0]), .b(u_csamul_cska32_fa16_9_xor1[0]), .cin(u_csamul_cska32_fa15_9_or0[0]), .fa_xor1(u_csamul_cska32_fa15_10_xor1), .fa_or0(u_csamul_cska32_fa15_10_or0));
  and_gate and_gate_u_csamul_cska32_and16_10(.a(a[16]), .b(b[10]), .out(u_csamul_cska32_and16_10));
  fa fa_u_csamul_cska32_fa16_10_out(.a(u_csamul_cska32_and16_10[0]), .b(u_csamul_cska32_fa17_9_xor1[0]), .cin(u_csamul_cska32_fa16_9_or0[0]), .fa_xor1(u_csamul_cska32_fa16_10_xor1), .fa_or0(u_csamul_cska32_fa16_10_or0));
  and_gate and_gate_u_csamul_cska32_and17_10(.a(a[17]), .b(b[10]), .out(u_csamul_cska32_and17_10));
  fa fa_u_csamul_cska32_fa17_10_out(.a(u_csamul_cska32_and17_10[0]), .b(u_csamul_cska32_fa18_9_xor1[0]), .cin(u_csamul_cska32_fa17_9_or0[0]), .fa_xor1(u_csamul_cska32_fa17_10_xor1), .fa_or0(u_csamul_cska32_fa17_10_or0));
  and_gate and_gate_u_csamul_cska32_and18_10(.a(a[18]), .b(b[10]), .out(u_csamul_cska32_and18_10));
  fa fa_u_csamul_cska32_fa18_10_out(.a(u_csamul_cska32_and18_10[0]), .b(u_csamul_cska32_fa19_9_xor1[0]), .cin(u_csamul_cska32_fa18_9_or0[0]), .fa_xor1(u_csamul_cska32_fa18_10_xor1), .fa_or0(u_csamul_cska32_fa18_10_or0));
  and_gate and_gate_u_csamul_cska32_and19_10(.a(a[19]), .b(b[10]), .out(u_csamul_cska32_and19_10));
  fa fa_u_csamul_cska32_fa19_10_out(.a(u_csamul_cska32_and19_10[0]), .b(u_csamul_cska32_fa20_9_xor1[0]), .cin(u_csamul_cska32_fa19_9_or0[0]), .fa_xor1(u_csamul_cska32_fa19_10_xor1), .fa_or0(u_csamul_cska32_fa19_10_or0));
  and_gate and_gate_u_csamul_cska32_and20_10(.a(a[20]), .b(b[10]), .out(u_csamul_cska32_and20_10));
  fa fa_u_csamul_cska32_fa20_10_out(.a(u_csamul_cska32_and20_10[0]), .b(u_csamul_cska32_fa21_9_xor1[0]), .cin(u_csamul_cska32_fa20_9_or0[0]), .fa_xor1(u_csamul_cska32_fa20_10_xor1), .fa_or0(u_csamul_cska32_fa20_10_or0));
  and_gate and_gate_u_csamul_cska32_and21_10(.a(a[21]), .b(b[10]), .out(u_csamul_cska32_and21_10));
  fa fa_u_csamul_cska32_fa21_10_out(.a(u_csamul_cska32_and21_10[0]), .b(u_csamul_cska32_fa22_9_xor1[0]), .cin(u_csamul_cska32_fa21_9_or0[0]), .fa_xor1(u_csamul_cska32_fa21_10_xor1), .fa_or0(u_csamul_cska32_fa21_10_or0));
  and_gate and_gate_u_csamul_cska32_and22_10(.a(a[22]), .b(b[10]), .out(u_csamul_cska32_and22_10));
  fa fa_u_csamul_cska32_fa22_10_out(.a(u_csamul_cska32_and22_10[0]), .b(u_csamul_cska32_fa23_9_xor1[0]), .cin(u_csamul_cska32_fa22_9_or0[0]), .fa_xor1(u_csamul_cska32_fa22_10_xor1), .fa_or0(u_csamul_cska32_fa22_10_or0));
  and_gate and_gate_u_csamul_cska32_and23_10(.a(a[23]), .b(b[10]), .out(u_csamul_cska32_and23_10));
  fa fa_u_csamul_cska32_fa23_10_out(.a(u_csamul_cska32_and23_10[0]), .b(u_csamul_cska32_fa24_9_xor1[0]), .cin(u_csamul_cska32_fa23_9_or0[0]), .fa_xor1(u_csamul_cska32_fa23_10_xor1), .fa_or0(u_csamul_cska32_fa23_10_or0));
  and_gate and_gate_u_csamul_cska32_and24_10(.a(a[24]), .b(b[10]), .out(u_csamul_cska32_and24_10));
  fa fa_u_csamul_cska32_fa24_10_out(.a(u_csamul_cska32_and24_10[0]), .b(u_csamul_cska32_fa25_9_xor1[0]), .cin(u_csamul_cska32_fa24_9_or0[0]), .fa_xor1(u_csamul_cska32_fa24_10_xor1), .fa_or0(u_csamul_cska32_fa24_10_or0));
  and_gate and_gate_u_csamul_cska32_and25_10(.a(a[25]), .b(b[10]), .out(u_csamul_cska32_and25_10));
  fa fa_u_csamul_cska32_fa25_10_out(.a(u_csamul_cska32_and25_10[0]), .b(u_csamul_cska32_fa26_9_xor1[0]), .cin(u_csamul_cska32_fa25_9_or0[0]), .fa_xor1(u_csamul_cska32_fa25_10_xor1), .fa_or0(u_csamul_cska32_fa25_10_or0));
  and_gate and_gate_u_csamul_cska32_and26_10(.a(a[26]), .b(b[10]), .out(u_csamul_cska32_and26_10));
  fa fa_u_csamul_cska32_fa26_10_out(.a(u_csamul_cska32_and26_10[0]), .b(u_csamul_cska32_fa27_9_xor1[0]), .cin(u_csamul_cska32_fa26_9_or0[0]), .fa_xor1(u_csamul_cska32_fa26_10_xor1), .fa_or0(u_csamul_cska32_fa26_10_or0));
  and_gate and_gate_u_csamul_cska32_and27_10(.a(a[27]), .b(b[10]), .out(u_csamul_cska32_and27_10));
  fa fa_u_csamul_cska32_fa27_10_out(.a(u_csamul_cska32_and27_10[0]), .b(u_csamul_cska32_fa28_9_xor1[0]), .cin(u_csamul_cska32_fa27_9_or0[0]), .fa_xor1(u_csamul_cska32_fa27_10_xor1), .fa_or0(u_csamul_cska32_fa27_10_or0));
  and_gate and_gate_u_csamul_cska32_and28_10(.a(a[28]), .b(b[10]), .out(u_csamul_cska32_and28_10));
  fa fa_u_csamul_cska32_fa28_10_out(.a(u_csamul_cska32_and28_10[0]), .b(u_csamul_cska32_fa29_9_xor1[0]), .cin(u_csamul_cska32_fa28_9_or0[0]), .fa_xor1(u_csamul_cska32_fa28_10_xor1), .fa_or0(u_csamul_cska32_fa28_10_or0));
  and_gate and_gate_u_csamul_cska32_and29_10(.a(a[29]), .b(b[10]), .out(u_csamul_cska32_and29_10));
  fa fa_u_csamul_cska32_fa29_10_out(.a(u_csamul_cska32_and29_10[0]), .b(u_csamul_cska32_fa30_9_xor1[0]), .cin(u_csamul_cska32_fa29_9_or0[0]), .fa_xor1(u_csamul_cska32_fa29_10_xor1), .fa_or0(u_csamul_cska32_fa29_10_or0));
  and_gate and_gate_u_csamul_cska32_and30_10(.a(a[30]), .b(b[10]), .out(u_csamul_cska32_and30_10));
  fa fa_u_csamul_cska32_fa30_10_out(.a(u_csamul_cska32_and30_10[0]), .b(u_csamul_cska32_and31_9[0]), .cin(u_csamul_cska32_fa30_9_or0[0]), .fa_xor1(u_csamul_cska32_fa30_10_xor1), .fa_or0(u_csamul_cska32_fa30_10_or0));
  and_gate and_gate_u_csamul_cska32_and31_10(.a(a[31]), .b(b[10]), .out(u_csamul_cska32_and31_10));
  and_gate and_gate_u_csamul_cska32_and0_11(.a(a[0]), .b(b[11]), .out(u_csamul_cska32_and0_11));
  fa fa_u_csamul_cska32_fa0_11_out(.a(u_csamul_cska32_and0_11[0]), .b(u_csamul_cska32_fa1_10_xor1[0]), .cin(u_csamul_cska32_fa0_10_or0[0]), .fa_xor1(u_csamul_cska32_fa0_11_xor1), .fa_or0(u_csamul_cska32_fa0_11_or0));
  and_gate and_gate_u_csamul_cska32_and1_11(.a(a[1]), .b(b[11]), .out(u_csamul_cska32_and1_11));
  fa fa_u_csamul_cska32_fa1_11_out(.a(u_csamul_cska32_and1_11[0]), .b(u_csamul_cska32_fa2_10_xor1[0]), .cin(u_csamul_cska32_fa1_10_or0[0]), .fa_xor1(u_csamul_cska32_fa1_11_xor1), .fa_or0(u_csamul_cska32_fa1_11_or0));
  and_gate and_gate_u_csamul_cska32_and2_11(.a(a[2]), .b(b[11]), .out(u_csamul_cska32_and2_11));
  fa fa_u_csamul_cska32_fa2_11_out(.a(u_csamul_cska32_and2_11[0]), .b(u_csamul_cska32_fa3_10_xor1[0]), .cin(u_csamul_cska32_fa2_10_or0[0]), .fa_xor1(u_csamul_cska32_fa2_11_xor1), .fa_or0(u_csamul_cska32_fa2_11_or0));
  and_gate and_gate_u_csamul_cska32_and3_11(.a(a[3]), .b(b[11]), .out(u_csamul_cska32_and3_11));
  fa fa_u_csamul_cska32_fa3_11_out(.a(u_csamul_cska32_and3_11[0]), .b(u_csamul_cska32_fa4_10_xor1[0]), .cin(u_csamul_cska32_fa3_10_or0[0]), .fa_xor1(u_csamul_cska32_fa3_11_xor1), .fa_or0(u_csamul_cska32_fa3_11_or0));
  and_gate and_gate_u_csamul_cska32_and4_11(.a(a[4]), .b(b[11]), .out(u_csamul_cska32_and4_11));
  fa fa_u_csamul_cska32_fa4_11_out(.a(u_csamul_cska32_and4_11[0]), .b(u_csamul_cska32_fa5_10_xor1[0]), .cin(u_csamul_cska32_fa4_10_or0[0]), .fa_xor1(u_csamul_cska32_fa4_11_xor1), .fa_or0(u_csamul_cska32_fa4_11_or0));
  and_gate and_gate_u_csamul_cska32_and5_11(.a(a[5]), .b(b[11]), .out(u_csamul_cska32_and5_11));
  fa fa_u_csamul_cska32_fa5_11_out(.a(u_csamul_cska32_and5_11[0]), .b(u_csamul_cska32_fa6_10_xor1[0]), .cin(u_csamul_cska32_fa5_10_or0[0]), .fa_xor1(u_csamul_cska32_fa5_11_xor1), .fa_or0(u_csamul_cska32_fa5_11_or0));
  and_gate and_gate_u_csamul_cska32_and6_11(.a(a[6]), .b(b[11]), .out(u_csamul_cska32_and6_11));
  fa fa_u_csamul_cska32_fa6_11_out(.a(u_csamul_cska32_and6_11[0]), .b(u_csamul_cska32_fa7_10_xor1[0]), .cin(u_csamul_cska32_fa6_10_or0[0]), .fa_xor1(u_csamul_cska32_fa6_11_xor1), .fa_or0(u_csamul_cska32_fa6_11_or0));
  and_gate and_gate_u_csamul_cska32_and7_11(.a(a[7]), .b(b[11]), .out(u_csamul_cska32_and7_11));
  fa fa_u_csamul_cska32_fa7_11_out(.a(u_csamul_cska32_and7_11[0]), .b(u_csamul_cska32_fa8_10_xor1[0]), .cin(u_csamul_cska32_fa7_10_or0[0]), .fa_xor1(u_csamul_cska32_fa7_11_xor1), .fa_or0(u_csamul_cska32_fa7_11_or0));
  and_gate and_gate_u_csamul_cska32_and8_11(.a(a[8]), .b(b[11]), .out(u_csamul_cska32_and8_11));
  fa fa_u_csamul_cska32_fa8_11_out(.a(u_csamul_cska32_and8_11[0]), .b(u_csamul_cska32_fa9_10_xor1[0]), .cin(u_csamul_cska32_fa8_10_or0[0]), .fa_xor1(u_csamul_cska32_fa8_11_xor1), .fa_or0(u_csamul_cska32_fa8_11_or0));
  and_gate and_gate_u_csamul_cska32_and9_11(.a(a[9]), .b(b[11]), .out(u_csamul_cska32_and9_11));
  fa fa_u_csamul_cska32_fa9_11_out(.a(u_csamul_cska32_and9_11[0]), .b(u_csamul_cska32_fa10_10_xor1[0]), .cin(u_csamul_cska32_fa9_10_or0[0]), .fa_xor1(u_csamul_cska32_fa9_11_xor1), .fa_or0(u_csamul_cska32_fa9_11_or0));
  and_gate and_gate_u_csamul_cska32_and10_11(.a(a[10]), .b(b[11]), .out(u_csamul_cska32_and10_11));
  fa fa_u_csamul_cska32_fa10_11_out(.a(u_csamul_cska32_and10_11[0]), .b(u_csamul_cska32_fa11_10_xor1[0]), .cin(u_csamul_cska32_fa10_10_or0[0]), .fa_xor1(u_csamul_cska32_fa10_11_xor1), .fa_or0(u_csamul_cska32_fa10_11_or0));
  and_gate and_gate_u_csamul_cska32_and11_11(.a(a[11]), .b(b[11]), .out(u_csamul_cska32_and11_11));
  fa fa_u_csamul_cska32_fa11_11_out(.a(u_csamul_cska32_and11_11[0]), .b(u_csamul_cska32_fa12_10_xor1[0]), .cin(u_csamul_cska32_fa11_10_or0[0]), .fa_xor1(u_csamul_cska32_fa11_11_xor1), .fa_or0(u_csamul_cska32_fa11_11_or0));
  and_gate and_gate_u_csamul_cska32_and12_11(.a(a[12]), .b(b[11]), .out(u_csamul_cska32_and12_11));
  fa fa_u_csamul_cska32_fa12_11_out(.a(u_csamul_cska32_and12_11[0]), .b(u_csamul_cska32_fa13_10_xor1[0]), .cin(u_csamul_cska32_fa12_10_or0[0]), .fa_xor1(u_csamul_cska32_fa12_11_xor1), .fa_or0(u_csamul_cska32_fa12_11_or0));
  and_gate and_gate_u_csamul_cska32_and13_11(.a(a[13]), .b(b[11]), .out(u_csamul_cska32_and13_11));
  fa fa_u_csamul_cska32_fa13_11_out(.a(u_csamul_cska32_and13_11[0]), .b(u_csamul_cska32_fa14_10_xor1[0]), .cin(u_csamul_cska32_fa13_10_or0[0]), .fa_xor1(u_csamul_cska32_fa13_11_xor1), .fa_or0(u_csamul_cska32_fa13_11_or0));
  and_gate and_gate_u_csamul_cska32_and14_11(.a(a[14]), .b(b[11]), .out(u_csamul_cska32_and14_11));
  fa fa_u_csamul_cska32_fa14_11_out(.a(u_csamul_cska32_and14_11[0]), .b(u_csamul_cska32_fa15_10_xor1[0]), .cin(u_csamul_cska32_fa14_10_or0[0]), .fa_xor1(u_csamul_cska32_fa14_11_xor1), .fa_or0(u_csamul_cska32_fa14_11_or0));
  and_gate and_gate_u_csamul_cska32_and15_11(.a(a[15]), .b(b[11]), .out(u_csamul_cska32_and15_11));
  fa fa_u_csamul_cska32_fa15_11_out(.a(u_csamul_cska32_and15_11[0]), .b(u_csamul_cska32_fa16_10_xor1[0]), .cin(u_csamul_cska32_fa15_10_or0[0]), .fa_xor1(u_csamul_cska32_fa15_11_xor1), .fa_or0(u_csamul_cska32_fa15_11_or0));
  and_gate and_gate_u_csamul_cska32_and16_11(.a(a[16]), .b(b[11]), .out(u_csamul_cska32_and16_11));
  fa fa_u_csamul_cska32_fa16_11_out(.a(u_csamul_cska32_and16_11[0]), .b(u_csamul_cska32_fa17_10_xor1[0]), .cin(u_csamul_cska32_fa16_10_or0[0]), .fa_xor1(u_csamul_cska32_fa16_11_xor1), .fa_or0(u_csamul_cska32_fa16_11_or0));
  and_gate and_gate_u_csamul_cska32_and17_11(.a(a[17]), .b(b[11]), .out(u_csamul_cska32_and17_11));
  fa fa_u_csamul_cska32_fa17_11_out(.a(u_csamul_cska32_and17_11[0]), .b(u_csamul_cska32_fa18_10_xor1[0]), .cin(u_csamul_cska32_fa17_10_or0[0]), .fa_xor1(u_csamul_cska32_fa17_11_xor1), .fa_or0(u_csamul_cska32_fa17_11_or0));
  and_gate and_gate_u_csamul_cska32_and18_11(.a(a[18]), .b(b[11]), .out(u_csamul_cska32_and18_11));
  fa fa_u_csamul_cska32_fa18_11_out(.a(u_csamul_cska32_and18_11[0]), .b(u_csamul_cska32_fa19_10_xor1[0]), .cin(u_csamul_cska32_fa18_10_or0[0]), .fa_xor1(u_csamul_cska32_fa18_11_xor1), .fa_or0(u_csamul_cska32_fa18_11_or0));
  and_gate and_gate_u_csamul_cska32_and19_11(.a(a[19]), .b(b[11]), .out(u_csamul_cska32_and19_11));
  fa fa_u_csamul_cska32_fa19_11_out(.a(u_csamul_cska32_and19_11[0]), .b(u_csamul_cska32_fa20_10_xor1[0]), .cin(u_csamul_cska32_fa19_10_or0[0]), .fa_xor1(u_csamul_cska32_fa19_11_xor1), .fa_or0(u_csamul_cska32_fa19_11_or0));
  and_gate and_gate_u_csamul_cska32_and20_11(.a(a[20]), .b(b[11]), .out(u_csamul_cska32_and20_11));
  fa fa_u_csamul_cska32_fa20_11_out(.a(u_csamul_cska32_and20_11[0]), .b(u_csamul_cska32_fa21_10_xor1[0]), .cin(u_csamul_cska32_fa20_10_or0[0]), .fa_xor1(u_csamul_cska32_fa20_11_xor1), .fa_or0(u_csamul_cska32_fa20_11_or0));
  and_gate and_gate_u_csamul_cska32_and21_11(.a(a[21]), .b(b[11]), .out(u_csamul_cska32_and21_11));
  fa fa_u_csamul_cska32_fa21_11_out(.a(u_csamul_cska32_and21_11[0]), .b(u_csamul_cska32_fa22_10_xor1[0]), .cin(u_csamul_cska32_fa21_10_or0[0]), .fa_xor1(u_csamul_cska32_fa21_11_xor1), .fa_or0(u_csamul_cska32_fa21_11_or0));
  and_gate and_gate_u_csamul_cska32_and22_11(.a(a[22]), .b(b[11]), .out(u_csamul_cska32_and22_11));
  fa fa_u_csamul_cska32_fa22_11_out(.a(u_csamul_cska32_and22_11[0]), .b(u_csamul_cska32_fa23_10_xor1[0]), .cin(u_csamul_cska32_fa22_10_or0[0]), .fa_xor1(u_csamul_cska32_fa22_11_xor1), .fa_or0(u_csamul_cska32_fa22_11_or0));
  and_gate and_gate_u_csamul_cska32_and23_11(.a(a[23]), .b(b[11]), .out(u_csamul_cska32_and23_11));
  fa fa_u_csamul_cska32_fa23_11_out(.a(u_csamul_cska32_and23_11[0]), .b(u_csamul_cska32_fa24_10_xor1[0]), .cin(u_csamul_cska32_fa23_10_or0[0]), .fa_xor1(u_csamul_cska32_fa23_11_xor1), .fa_or0(u_csamul_cska32_fa23_11_or0));
  and_gate and_gate_u_csamul_cska32_and24_11(.a(a[24]), .b(b[11]), .out(u_csamul_cska32_and24_11));
  fa fa_u_csamul_cska32_fa24_11_out(.a(u_csamul_cska32_and24_11[0]), .b(u_csamul_cska32_fa25_10_xor1[0]), .cin(u_csamul_cska32_fa24_10_or0[0]), .fa_xor1(u_csamul_cska32_fa24_11_xor1), .fa_or0(u_csamul_cska32_fa24_11_or0));
  and_gate and_gate_u_csamul_cska32_and25_11(.a(a[25]), .b(b[11]), .out(u_csamul_cska32_and25_11));
  fa fa_u_csamul_cska32_fa25_11_out(.a(u_csamul_cska32_and25_11[0]), .b(u_csamul_cska32_fa26_10_xor1[0]), .cin(u_csamul_cska32_fa25_10_or0[0]), .fa_xor1(u_csamul_cska32_fa25_11_xor1), .fa_or0(u_csamul_cska32_fa25_11_or0));
  and_gate and_gate_u_csamul_cska32_and26_11(.a(a[26]), .b(b[11]), .out(u_csamul_cska32_and26_11));
  fa fa_u_csamul_cska32_fa26_11_out(.a(u_csamul_cska32_and26_11[0]), .b(u_csamul_cska32_fa27_10_xor1[0]), .cin(u_csamul_cska32_fa26_10_or0[0]), .fa_xor1(u_csamul_cska32_fa26_11_xor1), .fa_or0(u_csamul_cska32_fa26_11_or0));
  and_gate and_gate_u_csamul_cska32_and27_11(.a(a[27]), .b(b[11]), .out(u_csamul_cska32_and27_11));
  fa fa_u_csamul_cska32_fa27_11_out(.a(u_csamul_cska32_and27_11[0]), .b(u_csamul_cska32_fa28_10_xor1[0]), .cin(u_csamul_cska32_fa27_10_or0[0]), .fa_xor1(u_csamul_cska32_fa27_11_xor1), .fa_or0(u_csamul_cska32_fa27_11_or0));
  and_gate and_gate_u_csamul_cska32_and28_11(.a(a[28]), .b(b[11]), .out(u_csamul_cska32_and28_11));
  fa fa_u_csamul_cska32_fa28_11_out(.a(u_csamul_cska32_and28_11[0]), .b(u_csamul_cska32_fa29_10_xor1[0]), .cin(u_csamul_cska32_fa28_10_or0[0]), .fa_xor1(u_csamul_cska32_fa28_11_xor1), .fa_or0(u_csamul_cska32_fa28_11_or0));
  and_gate and_gate_u_csamul_cska32_and29_11(.a(a[29]), .b(b[11]), .out(u_csamul_cska32_and29_11));
  fa fa_u_csamul_cska32_fa29_11_out(.a(u_csamul_cska32_and29_11[0]), .b(u_csamul_cska32_fa30_10_xor1[0]), .cin(u_csamul_cska32_fa29_10_or0[0]), .fa_xor1(u_csamul_cska32_fa29_11_xor1), .fa_or0(u_csamul_cska32_fa29_11_or0));
  and_gate and_gate_u_csamul_cska32_and30_11(.a(a[30]), .b(b[11]), .out(u_csamul_cska32_and30_11));
  fa fa_u_csamul_cska32_fa30_11_out(.a(u_csamul_cska32_and30_11[0]), .b(u_csamul_cska32_and31_10[0]), .cin(u_csamul_cska32_fa30_10_or0[0]), .fa_xor1(u_csamul_cska32_fa30_11_xor1), .fa_or0(u_csamul_cska32_fa30_11_or0));
  and_gate and_gate_u_csamul_cska32_and31_11(.a(a[31]), .b(b[11]), .out(u_csamul_cska32_and31_11));
  and_gate and_gate_u_csamul_cska32_and0_12(.a(a[0]), .b(b[12]), .out(u_csamul_cska32_and0_12));
  fa fa_u_csamul_cska32_fa0_12_out(.a(u_csamul_cska32_and0_12[0]), .b(u_csamul_cska32_fa1_11_xor1[0]), .cin(u_csamul_cska32_fa0_11_or0[0]), .fa_xor1(u_csamul_cska32_fa0_12_xor1), .fa_or0(u_csamul_cska32_fa0_12_or0));
  and_gate and_gate_u_csamul_cska32_and1_12(.a(a[1]), .b(b[12]), .out(u_csamul_cska32_and1_12));
  fa fa_u_csamul_cska32_fa1_12_out(.a(u_csamul_cska32_and1_12[0]), .b(u_csamul_cska32_fa2_11_xor1[0]), .cin(u_csamul_cska32_fa1_11_or0[0]), .fa_xor1(u_csamul_cska32_fa1_12_xor1), .fa_or0(u_csamul_cska32_fa1_12_or0));
  and_gate and_gate_u_csamul_cska32_and2_12(.a(a[2]), .b(b[12]), .out(u_csamul_cska32_and2_12));
  fa fa_u_csamul_cska32_fa2_12_out(.a(u_csamul_cska32_and2_12[0]), .b(u_csamul_cska32_fa3_11_xor1[0]), .cin(u_csamul_cska32_fa2_11_or0[0]), .fa_xor1(u_csamul_cska32_fa2_12_xor1), .fa_or0(u_csamul_cska32_fa2_12_or0));
  and_gate and_gate_u_csamul_cska32_and3_12(.a(a[3]), .b(b[12]), .out(u_csamul_cska32_and3_12));
  fa fa_u_csamul_cska32_fa3_12_out(.a(u_csamul_cska32_and3_12[0]), .b(u_csamul_cska32_fa4_11_xor1[0]), .cin(u_csamul_cska32_fa3_11_or0[0]), .fa_xor1(u_csamul_cska32_fa3_12_xor1), .fa_or0(u_csamul_cska32_fa3_12_or0));
  and_gate and_gate_u_csamul_cska32_and4_12(.a(a[4]), .b(b[12]), .out(u_csamul_cska32_and4_12));
  fa fa_u_csamul_cska32_fa4_12_out(.a(u_csamul_cska32_and4_12[0]), .b(u_csamul_cska32_fa5_11_xor1[0]), .cin(u_csamul_cska32_fa4_11_or0[0]), .fa_xor1(u_csamul_cska32_fa4_12_xor1), .fa_or0(u_csamul_cska32_fa4_12_or0));
  and_gate and_gate_u_csamul_cska32_and5_12(.a(a[5]), .b(b[12]), .out(u_csamul_cska32_and5_12));
  fa fa_u_csamul_cska32_fa5_12_out(.a(u_csamul_cska32_and5_12[0]), .b(u_csamul_cska32_fa6_11_xor1[0]), .cin(u_csamul_cska32_fa5_11_or0[0]), .fa_xor1(u_csamul_cska32_fa5_12_xor1), .fa_or0(u_csamul_cska32_fa5_12_or0));
  and_gate and_gate_u_csamul_cska32_and6_12(.a(a[6]), .b(b[12]), .out(u_csamul_cska32_and6_12));
  fa fa_u_csamul_cska32_fa6_12_out(.a(u_csamul_cska32_and6_12[0]), .b(u_csamul_cska32_fa7_11_xor1[0]), .cin(u_csamul_cska32_fa6_11_or0[0]), .fa_xor1(u_csamul_cska32_fa6_12_xor1), .fa_or0(u_csamul_cska32_fa6_12_or0));
  and_gate and_gate_u_csamul_cska32_and7_12(.a(a[7]), .b(b[12]), .out(u_csamul_cska32_and7_12));
  fa fa_u_csamul_cska32_fa7_12_out(.a(u_csamul_cska32_and7_12[0]), .b(u_csamul_cska32_fa8_11_xor1[0]), .cin(u_csamul_cska32_fa7_11_or0[0]), .fa_xor1(u_csamul_cska32_fa7_12_xor1), .fa_or0(u_csamul_cska32_fa7_12_or0));
  and_gate and_gate_u_csamul_cska32_and8_12(.a(a[8]), .b(b[12]), .out(u_csamul_cska32_and8_12));
  fa fa_u_csamul_cska32_fa8_12_out(.a(u_csamul_cska32_and8_12[0]), .b(u_csamul_cska32_fa9_11_xor1[0]), .cin(u_csamul_cska32_fa8_11_or0[0]), .fa_xor1(u_csamul_cska32_fa8_12_xor1), .fa_or0(u_csamul_cska32_fa8_12_or0));
  and_gate and_gate_u_csamul_cska32_and9_12(.a(a[9]), .b(b[12]), .out(u_csamul_cska32_and9_12));
  fa fa_u_csamul_cska32_fa9_12_out(.a(u_csamul_cska32_and9_12[0]), .b(u_csamul_cska32_fa10_11_xor1[0]), .cin(u_csamul_cska32_fa9_11_or0[0]), .fa_xor1(u_csamul_cska32_fa9_12_xor1), .fa_or0(u_csamul_cska32_fa9_12_or0));
  and_gate and_gate_u_csamul_cska32_and10_12(.a(a[10]), .b(b[12]), .out(u_csamul_cska32_and10_12));
  fa fa_u_csamul_cska32_fa10_12_out(.a(u_csamul_cska32_and10_12[0]), .b(u_csamul_cska32_fa11_11_xor1[0]), .cin(u_csamul_cska32_fa10_11_or0[0]), .fa_xor1(u_csamul_cska32_fa10_12_xor1), .fa_or0(u_csamul_cska32_fa10_12_or0));
  and_gate and_gate_u_csamul_cska32_and11_12(.a(a[11]), .b(b[12]), .out(u_csamul_cska32_and11_12));
  fa fa_u_csamul_cska32_fa11_12_out(.a(u_csamul_cska32_and11_12[0]), .b(u_csamul_cska32_fa12_11_xor1[0]), .cin(u_csamul_cska32_fa11_11_or0[0]), .fa_xor1(u_csamul_cska32_fa11_12_xor1), .fa_or0(u_csamul_cska32_fa11_12_or0));
  and_gate and_gate_u_csamul_cska32_and12_12(.a(a[12]), .b(b[12]), .out(u_csamul_cska32_and12_12));
  fa fa_u_csamul_cska32_fa12_12_out(.a(u_csamul_cska32_and12_12[0]), .b(u_csamul_cska32_fa13_11_xor1[0]), .cin(u_csamul_cska32_fa12_11_or0[0]), .fa_xor1(u_csamul_cska32_fa12_12_xor1), .fa_or0(u_csamul_cska32_fa12_12_or0));
  and_gate and_gate_u_csamul_cska32_and13_12(.a(a[13]), .b(b[12]), .out(u_csamul_cska32_and13_12));
  fa fa_u_csamul_cska32_fa13_12_out(.a(u_csamul_cska32_and13_12[0]), .b(u_csamul_cska32_fa14_11_xor1[0]), .cin(u_csamul_cska32_fa13_11_or0[0]), .fa_xor1(u_csamul_cska32_fa13_12_xor1), .fa_or0(u_csamul_cska32_fa13_12_or0));
  and_gate and_gate_u_csamul_cska32_and14_12(.a(a[14]), .b(b[12]), .out(u_csamul_cska32_and14_12));
  fa fa_u_csamul_cska32_fa14_12_out(.a(u_csamul_cska32_and14_12[0]), .b(u_csamul_cska32_fa15_11_xor1[0]), .cin(u_csamul_cska32_fa14_11_or0[0]), .fa_xor1(u_csamul_cska32_fa14_12_xor1), .fa_or0(u_csamul_cska32_fa14_12_or0));
  and_gate and_gate_u_csamul_cska32_and15_12(.a(a[15]), .b(b[12]), .out(u_csamul_cska32_and15_12));
  fa fa_u_csamul_cska32_fa15_12_out(.a(u_csamul_cska32_and15_12[0]), .b(u_csamul_cska32_fa16_11_xor1[0]), .cin(u_csamul_cska32_fa15_11_or0[0]), .fa_xor1(u_csamul_cska32_fa15_12_xor1), .fa_or0(u_csamul_cska32_fa15_12_or0));
  and_gate and_gate_u_csamul_cska32_and16_12(.a(a[16]), .b(b[12]), .out(u_csamul_cska32_and16_12));
  fa fa_u_csamul_cska32_fa16_12_out(.a(u_csamul_cska32_and16_12[0]), .b(u_csamul_cska32_fa17_11_xor1[0]), .cin(u_csamul_cska32_fa16_11_or0[0]), .fa_xor1(u_csamul_cska32_fa16_12_xor1), .fa_or0(u_csamul_cska32_fa16_12_or0));
  and_gate and_gate_u_csamul_cska32_and17_12(.a(a[17]), .b(b[12]), .out(u_csamul_cska32_and17_12));
  fa fa_u_csamul_cska32_fa17_12_out(.a(u_csamul_cska32_and17_12[0]), .b(u_csamul_cska32_fa18_11_xor1[0]), .cin(u_csamul_cska32_fa17_11_or0[0]), .fa_xor1(u_csamul_cska32_fa17_12_xor1), .fa_or0(u_csamul_cska32_fa17_12_or0));
  and_gate and_gate_u_csamul_cska32_and18_12(.a(a[18]), .b(b[12]), .out(u_csamul_cska32_and18_12));
  fa fa_u_csamul_cska32_fa18_12_out(.a(u_csamul_cska32_and18_12[0]), .b(u_csamul_cska32_fa19_11_xor1[0]), .cin(u_csamul_cska32_fa18_11_or0[0]), .fa_xor1(u_csamul_cska32_fa18_12_xor1), .fa_or0(u_csamul_cska32_fa18_12_or0));
  and_gate and_gate_u_csamul_cska32_and19_12(.a(a[19]), .b(b[12]), .out(u_csamul_cska32_and19_12));
  fa fa_u_csamul_cska32_fa19_12_out(.a(u_csamul_cska32_and19_12[0]), .b(u_csamul_cska32_fa20_11_xor1[0]), .cin(u_csamul_cska32_fa19_11_or0[0]), .fa_xor1(u_csamul_cska32_fa19_12_xor1), .fa_or0(u_csamul_cska32_fa19_12_or0));
  and_gate and_gate_u_csamul_cska32_and20_12(.a(a[20]), .b(b[12]), .out(u_csamul_cska32_and20_12));
  fa fa_u_csamul_cska32_fa20_12_out(.a(u_csamul_cska32_and20_12[0]), .b(u_csamul_cska32_fa21_11_xor1[0]), .cin(u_csamul_cska32_fa20_11_or0[0]), .fa_xor1(u_csamul_cska32_fa20_12_xor1), .fa_or0(u_csamul_cska32_fa20_12_or0));
  and_gate and_gate_u_csamul_cska32_and21_12(.a(a[21]), .b(b[12]), .out(u_csamul_cska32_and21_12));
  fa fa_u_csamul_cska32_fa21_12_out(.a(u_csamul_cska32_and21_12[0]), .b(u_csamul_cska32_fa22_11_xor1[0]), .cin(u_csamul_cska32_fa21_11_or0[0]), .fa_xor1(u_csamul_cska32_fa21_12_xor1), .fa_or0(u_csamul_cska32_fa21_12_or0));
  and_gate and_gate_u_csamul_cska32_and22_12(.a(a[22]), .b(b[12]), .out(u_csamul_cska32_and22_12));
  fa fa_u_csamul_cska32_fa22_12_out(.a(u_csamul_cska32_and22_12[0]), .b(u_csamul_cska32_fa23_11_xor1[0]), .cin(u_csamul_cska32_fa22_11_or0[0]), .fa_xor1(u_csamul_cska32_fa22_12_xor1), .fa_or0(u_csamul_cska32_fa22_12_or0));
  and_gate and_gate_u_csamul_cska32_and23_12(.a(a[23]), .b(b[12]), .out(u_csamul_cska32_and23_12));
  fa fa_u_csamul_cska32_fa23_12_out(.a(u_csamul_cska32_and23_12[0]), .b(u_csamul_cska32_fa24_11_xor1[0]), .cin(u_csamul_cska32_fa23_11_or0[0]), .fa_xor1(u_csamul_cska32_fa23_12_xor1), .fa_or0(u_csamul_cska32_fa23_12_or0));
  and_gate and_gate_u_csamul_cska32_and24_12(.a(a[24]), .b(b[12]), .out(u_csamul_cska32_and24_12));
  fa fa_u_csamul_cska32_fa24_12_out(.a(u_csamul_cska32_and24_12[0]), .b(u_csamul_cska32_fa25_11_xor1[0]), .cin(u_csamul_cska32_fa24_11_or0[0]), .fa_xor1(u_csamul_cska32_fa24_12_xor1), .fa_or0(u_csamul_cska32_fa24_12_or0));
  and_gate and_gate_u_csamul_cska32_and25_12(.a(a[25]), .b(b[12]), .out(u_csamul_cska32_and25_12));
  fa fa_u_csamul_cska32_fa25_12_out(.a(u_csamul_cska32_and25_12[0]), .b(u_csamul_cska32_fa26_11_xor1[0]), .cin(u_csamul_cska32_fa25_11_or0[0]), .fa_xor1(u_csamul_cska32_fa25_12_xor1), .fa_or0(u_csamul_cska32_fa25_12_or0));
  and_gate and_gate_u_csamul_cska32_and26_12(.a(a[26]), .b(b[12]), .out(u_csamul_cska32_and26_12));
  fa fa_u_csamul_cska32_fa26_12_out(.a(u_csamul_cska32_and26_12[0]), .b(u_csamul_cska32_fa27_11_xor1[0]), .cin(u_csamul_cska32_fa26_11_or0[0]), .fa_xor1(u_csamul_cska32_fa26_12_xor1), .fa_or0(u_csamul_cska32_fa26_12_or0));
  and_gate and_gate_u_csamul_cska32_and27_12(.a(a[27]), .b(b[12]), .out(u_csamul_cska32_and27_12));
  fa fa_u_csamul_cska32_fa27_12_out(.a(u_csamul_cska32_and27_12[0]), .b(u_csamul_cska32_fa28_11_xor1[0]), .cin(u_csamul_cska32_fa27_11_or0[0]), .fa_xor1(u_csamul_cska32_fa27_12_xor1), .fa_or0(u_csamul_cska32_fa27_12_or0));
  and_gate and_gate_u_csamul_cska32_and28_12(.a(a[28]), .b(b[12]), .out(u_csamul_cska32_and28_12));
  fa fa_u_csamul_cska32_fa28_12_out(.a(u_csamul_cska32_and28_12[0]), .b(u_csamul_cska32_fa29_11_xor1[0]), .cin(u_csamul_cska32_fa28_11_or0[0]), .fa_xor1(u_csamul_cska32_fa28_12_xor1), .fa_or0(u_csamul_cska32_fa28_12_or0));
  and_gate and_gate_u_csamul_cska32_and29_12(.a(a[29]), .b(b[12]), .out(u_csamul_cska32_and29_12));
  fa fa_u_csamul_cska32_fa29_12_out(.a(u_csamul_cska32_and29_12[0]), .b(u_csamul_cska32_fa30_11_xor1[0]), .cin(u_csamul_cska32_fa29_11_or0[0]), .fa_xor1(u_csamul_cska32_fa29_12_xor1), .fa_or0(u_csamul_cska32_fa29_12_or0));
  and_gate and_gate_u_csamul_cska32_and30_12(.a(a[30]), .b(b[12]), .out(u_csamul_cska32_and30_12));
  fa fa_u_csamul_cska32_fa30_12_out(.a(u_csamul_cska32_and30_12[0]), .b(u_csamul_cska32_and31_11[0]), .cin(u_csamul_cska32_fa30_11_or0[0]), .fa_xor1(u_csamul_cska32_fa30_12_xor1), .fa_or0(u_csamul_cska32_fa30_12_or0));
  and_gate and_gate_u_csamul_cska32_and31_12(.a(a[31]), .b(b[12]), .out(u_csamul_cska32_and31_12));
  and_gate and_gate_u_csamul_cska32_and0_13(.a(a[0]), .b(b[13]), .out(u_csamul_cska32_and0_13));
  fa fa_u_csamul_cska32_fa0_13_out(.a(u_csamul_cska32_and0_13[0]), .b(u_csamul_cska32_fa1_12_xor1[0]), .cin(u_csamul_cska32_fa0_12_or0[0]), .fa_xor1(u_csamul_cska32_fa0_13_xor1), .fa_or0(u_csamul_cska32_fa0_13_or0));
  and_gate and_gate_u_csamul_cska32_and1_13(.a(a[1]), .b(b[13]), .out(u_csamul_cska32_and1_13));
  fa fa_u_csamul_cska32_fa1_13_out(.a(u_csamul_cska32_and1_13[0]), .b(u_csamul_cska32_fa2_12_xor1[0]), .cin(u_csamul_cska32_fa1_12_or0[0]), .fa_xor1(u_csamul_cska32_fa1_13_xor1), .fa_or0(u_csamul_cska32_fa1_13_or0));
  and_gate and_gate_u_csamul_cska32_and2_13(.a(a[2]), .b(b[13]), .out(u_csamul_cska32_and2_13));
  fa fa_u_csamul_cska32_fa2_13_out(.a(u_csamul_cska32_and2_13[0]), .b(u_csamul_cska32_fa3_12_xor1[0]), .cin(u_csamul_cska32_fa2_12_or0[0]), .fa_xor1(u_csamul_cska32_fa2_13_xor1), .fa_or0(u_csamul_cska32_fa2_13_or0));
  and_gate and_gate_u_csamul_cska32_and3_13(.a(a[3]), .b(b[13]), .out(u_csamul_cska32_and3_13));
  fa fa_u_csamul_cska32_fa3_13_out(.a(u_csamul_cska32_and3_13[0]), .b(u_csamul_cska32_fa4_12_xor1[0]), .cin(u_csamul_cska32_fa3_12_or0[0]), .fa_xor1(u_csamul_cska32_fa3_13_xor1), .fa_or0(u_csamul_cska32_fa3_13_or0));
  and_gate and_gate_u_csamul_cska32_and4_13(.a(a[4]), .b(b[13]), .out(u_csamul_cska32_and4_13));
  fa fa_u_csamul_cska32_fa4_13_out(.a(u_csamul_cska32_and4_13[0]), .b(u_csamul_cska32_fa5_12_xor1[0]), .cin(u_csamul_cska32_fa4_12_or0[0]), .fa_xor1(u_csamul_cska32_fa4_13_xor1), .fa_or0(u_csamul_cska32_fa4_13_or0));
  and_gate and_gate_u_csamul_cska32_and5_13(.a(a[5]), .b(b[13]), .out(u_csamul_cska32_and5_13));
  fa fa_u_csamul_cska32_fa5_13_out(.a(u_csamul_cska32_and5_13[0]), .b(u_csamul_cska32_fa6_12_xor1[0]), .cin(u_csamul_cska32_fa5_12_or0[0]), .fa_xor1(u_csamul_cska32_fa5_13_xor1), .fa_or0(u_csamul_cska32_fa5_13_or0));
  and_gate and_gate_u_csamul_cska32_and6_13(.a(a[6]), .b(b[13]), .out(u_csamul_cska32_and6_13));
  fa fa_u_csamul_cska32_fa6_13_out(.a(u_csamul_cska32_and6_13[0]), .b(u_csamul_cska32_fa7_12_xor1[0]), .cin(u_csamul_cska32_fa6_12_or0[0]), .fa_xor1(u_csamul_cska32_fa6_13_xor1), .fa_or0(u_csamul_cska32_fa6_13_or0));
  and_gate and_gate_u_csamul_cska32_and7_13(.a(a[7]), .b(b[13]), .out(u_csamul_cska32_and7_13));
  fa fa_u_csamul_cska32_fa7_13_out(.a(u_csamul_cska32_and7_13[0]), .b(u_csamul_cska32_fa8_12_xor1[0]), .cin(u_csamul_cska32_fa7_12_or0[0]), .fa_xor1(u_csamul_cska32_fa7_13_xor1), .fa_or0(u_csamul_cska32_fa7_13_or0));
  and_gate and_gate_u_csamul_cska32_and8_13(.a(a[8]), .b(b[13]), .out(u_csamul_cska32_and8_13));
  fa fa_u_csamul_cska32_fa8_13_out(.a(u_csamul_cska32_and8_13[0]), .b(u_csamul_cska32_fa9_12_xor1[0]), .cin(u_csamul_cska32_fa8_12_or0[0]), .fa_xor1(u_csamul_cska32_fa8_13_xor1), .fa_or0(u_csamul_cska32_fa8_13_or0));
  and_gate and_gate_u_csamul_cska32_and9_13(.a(a[9]), .b(b[13]), .out(u_csamul_cska32_and9_13));
  fa fa_u_csamul_cska32_fa9_13_out(.a(u_csamul_cska32_and9_13[0]), .b(u_csamul_cska32_fa10_12_xor1[0]), .cin(u_csamul_cska32_fa9_12_or0[0]), .fa_xor1(u_csamul_cska32_fa9_13_xor1), .fa_or0(u_csamul_cska32_fa9_13_or0));
  and_gate and_gate_u_csamul_cska32_and10_13(.a(a[10]), .b(b[13]), .out(u_csamul_cska32_and10_13));
  fa fa_u_csamul_cska32_fa10_13_out(.a(u_csamul_cska32_and10_13[0]), .b(u_csamul_cska32_fa11_12_xor1[0]), .cin(u_csamul_cska32_fa10_12_or0[0]), .fa_xor1(u_csamul_cska32_fa10_13_xor1), .fa_or0(u_csamul_cska32_fa10_13_or0));
  and_gate and_gate_u_csamul_cska32_and11_13(.a(a[11]), .b(b[13]), .out(u_csamul_cska32_and11_13));
  fa fa_u_csamul_cska32_fa11_13_out(.a(u_csamul_cska32_and11_13[0]), .b(u_csamul_cska32_fa12_12_xor1[0]), .cin(u_csamul_cska32_fa11_12_or0[0]), .fa_xor1(u_csamul_cska32_fa11_13_xor1), .fa_or0(u_csamul_cska32_fa11_13_or0));
  and_gate and_gate_u_csamul_cska32_and12_13(.a(a[12]), .b(b[13]), .out(u_csamul_cska32_and12_13));
  fa fa_u_csamul_cska32_fa12_13_out(.a(u_csamul_cska32_and12_13[0]), .b(u_csamul_cska32_fa13_12_xor1[0]), .cin(u_csamul_cska32_fa12_12_or0[0]), .fa_xor1(u_csamul_cska32_fa12_13_xor1), .fa_or0(u_csamul_cska32_fa12_13_or0));
  and_gate and_gate_u_csamul_cska32_and13_13(.a(a[13]), .b(b[13]), .out(u_csamul_cska32_and13_13));
  fa fa_u_csamul_cska32_fa13_13_out(.a(u_csamul_cska32_and13_13[0]), .b(u_csamul_cska32_fa14_12_xor1[0]), .cin(u_csamul_cska32_fa13_12_or0[0]), .fa_xor1(u_csamul_cska32_fa13_13_xor1), .fa_or0(u_csamul_cska32_fa13_13_or0));
  and_gate and_gate_u_csamul_cska32_and14_13(.a(a[14]), .b(b[13]), .out(u_csamul_cska32_and14_13));
  fa fa_u_csamul_cska32_fa14_13_out(.a(u_csamul_cska32_and14_13[0]), .b(u_csamul_cska32_fa15_12_xor1[0]), .cin(u_csamul_cska32_fa14_12_or0[0]), .fa_xor1(u_csamul_cska32_fa14_13_xor1), .fa_or0(u_csamul_cska32_fa14_13_or0));
  and_gate and_gate_u_csamul_cska32_and15_13(.a(a[15]), .b(b[13]), .out(u_csamul_cska32_and15_13));
  fa fa_u_csamul_cska32_fa15_13_out(.a(u_csamul_cska32_and15_13[0]), .b(u_csamul_cska32_fa16_12_xor1[0]), .cin(u_csamul_cska32_fa15_12_or0[0]), .fa_xor1(u_csamul_cska32_fa15_13_xor1), .fa_or0(u_csamul_cska32_fa15_13_or0));
  and_gate and_gate_u_csamul_cska32_and16_13(.a(a[16]), .b(b[13]), .out(u_csamul_cska32_and16_13));
  fa fa_u_csamul_cska32_fa16_13_out(.a(u_csamul_cska32_and16_13[0]), .b(u_csamul_cska32_fa17_12_xor1[0]), .cin(u_csamul_cska32_fa16_12_or0[0]), .fa_xor1(u_csamul_cska32_fa16_13_xor1), .fa_or0(u_csamul_cska32_fa16_13_or0));
  and_gate and_gate_u_csamul_cska32_and17_13(.a(a[17]), .b(b[13]), .out(u_csamul_cska32_and17_13));
  fa fa_u_csamul_cska32_fa17_13_out(.a(u_csamul_cska32_and17_13[0]), .b(u_csamul_cska32_fa18_12_xor1[0]), .cin(u_csamul_cska32_fa17_12_or0[0]), .fa_xor1(u_csamul_cska32_fa17_13_xor1), .fa_or0(u_csamul_cska32_fa17_13_or0));
  and_gate and_gate_u_csamul_cska32_and18_13(.a(a[18]), .b(b[13]), .out(u_csamul_cska32_and18_13));
  fa fa_u_csamul_cska32_fa18_13_out(.a(u_csamul_cska32_and18_13[0]), .b(u_csamul_cska32_fa19_12_xor1[0]), .cin(u_csamul_cska32_fa18_12_or0[0]), .fa_xor1(u_csamul_cska32_fa18_13_xor1), .fa_or0(u_csamul_cska32_fa18_13_or0));
  and_gate and_gate_u_csamul_cska32_and19_13(.a(a[19]), .b(b[13]), .out(u_csamul_cska32_and19_13));
  fa fa_u_csamul_cska32_fa19_13_out(.a(u_csamul_cska32_and19_13[0]), .b(u_csamul_cska32_fa20_12_xor1[0]), .cin(u_csamul_cska32_fa19_12_or0[0]), .fa_xor1(u_csamul_cska32_fa19_13_xor1), .fa_or0(u_csamul_cska32_fa19_13_or0));
  and_gate and_gate_u_csamul_cska32_and20_13(.a(a[20]), .b(b[13]), .out(u_csamul_cska32_and20_13));
  fa fa_u_csamul_cska32_fa20_13_out(.a(u_csamul_cska32_and20_13[0]), .b(u_csamul_cska32_fa21_12_xor1[0]), .cin(u_csamul_cska32_fa20_12_or0[0]), .fa_xor1(u_csamul_cska32_fa20_13_xor1), .fa_or0(u_csamul_cska32_fa20_13_or0));
  and_gate and_gate_u_csamul_cska32_and21_13(.a(a[21]), .b(b[13]), .out(u_csamul_cska32_and21_13));
  fa fa_u_csamul_cska32_fa21_13_out(.a(u_csamul_cska32_and21_13[0]), .b(u_csamul_cska32_fa22_12_xor1[0]), .cin(u_csamul_cska32_fa21_12_or0[0]), .fa_xor1(u_csamul_cska32_fa21_13_xor1), .fa_or0(u_csamul_cska32_fa21_13_or0));
  and_gate and_gate_u_csamul_cska32_and22_13(.a(a[22]), .b(b[13]), .out(u_csamul_cska32_and22_13));
  fa fa_u_csamul_cska32_fa22_13_out(.a(u_csamul_cska32_and22_13[0]), .b(u_csamul_cska32_fa23_12_xor1[0]), .cin(u_csamul_cska32_fa22_12_or0[0]), .fa_xor1(u_csamul_cska32_fa22_13_xor1), .fa_or0(u_csamul_cska32_fa22_13_or0));
  and_gate and_gate_u_csamul_cska32_and23_13(.a(a[23]), .b(b[13]), .out(u_csamul_cska32_and23_13));
  fa fa_u_csamul_cska32_fa23_13_out(.a(u_csamul_cska32_and23_13[0]), .b(u_csamul_cska32_fa24_12_xor1[0]), .cin(u_csamul_cska32_fa23_12_or0[0]), .fa_xor1(u_csamul_cska32_fa23_13_xor1), .fa_or0(u_csamul_cska32_fa23_13_or0));
  and_gate and_gate_u_csamul_cska32_and24_13(.a(a[24]), .b(b[13]), .out(u_csamul_cska32_and24_13));
  fa fa_u_csamul_cska32_fa24_13_out(.a(u_csamul_cska32_and24_13[0]), .b(u_csamul_cska32_fa25_12_xor1[0]), .cin(u_csamul_cska32_fa24_12_or0[0]), .fa_xor1(u_csamul_cska32_fa24_13_xor1), .fa_or0(u_csamul_cska32_fa24_13_or0));
  and_gate and_gate_u_csamul_cska32_and25_13(.a(a[25]), .b(b[13]), .out(u_csamul_cska32_and25_13));
  fa fa_u_csamul_cska32_fa25_13_out(.a(u_csamul_cska32_and25_13[0]), .b(u_csamul_cska32_fa26_12_xor1[0]), .cin(u_csamul_cska32_fa25_12_or0[0]), .fa_xor1(u_csamul_cska32_fa25_13_xor1), .fa_or0(u_csamul_cska32_fa25_13_or0));
  and_gate and_gate_u_csamul_cska32_and26_13(.a(a[26]), .b(b[13]), .out(u_csamul_cska32_and26_13));
  fa fa_u_csamul_cska32_fa26_13_out(.a(u_csamul_cska32_and26_13[0]), .b(u_csamul_cska32_fa27_12_xor1[0]), .cin(u_csamul_cska32_fa26_12_or0[0]), .fa_xor1(u_csamul_cska32_fa26_13_xor1), .fa_or0(u_csamul_cska32_fa26_13_or0));
  and_gate and_gate_u_csamul_cska32_and27_13(.a(a[27]), .b(b[13]), .out(u_csamul_cska32_and27_13));
  fa fa_u_csamul_cska32_fa27_13_out(.a(u_csamul_cska32_and27_13[0]), .b(u_csamul_cska32_fa28_12_xor1[0]), .cin(u_csamul_cska32_fa27_12_or0[0]), .fa_xor1(u_csamul_cska32_fa27_13_xor1), .fa_or0(u_csamul_cska32_fa27_13_or0));
  and_gate and_gate_u_csamul_cska32_and28_13(.a(a[28]), .b(b[13]), .out(u_csamul_cska32_and28_13));
  fa fa_u_csamul_cska32_fa28_13_out(.a(u_csamul_cska32_and28_13[0]), .b(u_csamul_cska32_fa29_12_xor1[0]), .cin(u_csamul_cska32_fa28_12_or0[0]), .fa_xor1(u_csamul_cska32_fa28_13_xor1), .fa_or0(u_csamul_cska32_fa28_13_or0));
  and_gate and_gate_u_csamul_cska32_and29_13(.a(a[29]), .b(b[13]), .out(u_csamul_cska32_and29_13));
  fa fa_u_csamul_cska32_fa29_13_out(.a(u_csamul_cska32_and29_13[0]), .b(u_csamul_cska32_fa30_12_xor1[0]), .cin(u_csamul_cska32_fa29_12_or0[0]), .fa_xor1(u_csamul_cska32_fa29_13_xor1), .fa_or0(u_csamul_cska32_fa29_13_or0));
  and_gate and_gate_u_csamul_cska32_and30_13(.a(a[30]), .b(b[13]), .out(u_csamul_cska32_and30_13));
  fa fa_u_csamul_cska32_fa30_13_out(.a(u_csamul_cska32_and30_13[0]), .b(u_csamul_cska32_and31_12[0]), .cin(u_csamul_cska32_fa30_12_or0[0]), .fa_xor1(u_csamul_cska32_fa30_13_xor1), .fa_or0(u_csamul_cska32_fa30_13_or0));
  and_gate and_gate_u_csamul_cska32_and31_13(.a(a[31]), .b(b[13]), .out(u_csamul_cska32_and31_13));
  and_gate and_gate_u_csamul_cska32_and0_14(.a(a[0]), .b(b[14]), .out(u_csamul_cska32_and0_14));
  fa fa_u_csamul_cska32_fa0_14_out(.a(u_csamul_cska32_and0_14[0]), .b(u_csamul_cska32_fa1_13_xor1[0]), .cin(u_csamul_cska32_fa0_13_or0[0]), .fa_xor1(u_csamul_cska32_fa0_14_xor1), .fa_or0(u_csamul_cska32_fa0_14_or0));
  and_gate and_gate_u_csamul_cska32_and1_14(.a(a[1]), .b(b[14]), .out(u_csamul_cska32_and1_14));
  fa fa_u_csamul_cska32_fa1_14_out(.a(u_csamul_cska32_and1_14[0]), .b(u_csamul_cska32_fa2_13_xor1[0]), .cin(u_csamul_cska32_fa1_13_or0[0]), .fa_xor1(u_csamul_cska32_fa1_14_xor1), .fa_or0(u_csamul_cska32_fa1_14_or0));
  and_gate and_gate_u_csamul_cska32_and2_14(.a(a[2]), .b(b[14]), .out(u_csamul_cska32_and2_14));
  fa fa_u_csamul_cska32_fa2_14_out(.a(u_csamul_cska32_and2_14[0]), .b(u_csamul_cska32_fa3_13_xor1[0]), .cin(u_csamul_cska32_fa2_13_or0[0]), .fa_xor1(u_csamul_cska32_fa2_14_xor1), .fa_or0(u_csamul_cska32_fa2_14_or0));
  and_gate and_gate_u_csamul_cska32_and3_14(.a(a[3]), .b(b[14]), .out(u_csamul_cska32_and3_14));
  fa fa_u_csamul_cska32_fa3_14_out(.a(u_csamul_cska32_and3_14[0]), .b(u_csamul_cska32_fa4_13_xor1[0]), .cin(u_csamul_cska32_fa3_13_or0[0]), .fa_xor1(u_csamul_cska32_fa3_14_xor1), .fa_or0(u_csamul_cska32_fa3_14_or0));
  and_gate and_gate_u_csamul_cska32_and4_14(.a(a[4]), .b(b[14]), .out(u_csamul_cska32_and4_14));
  fa fa_u_csamul_cska32_fa4_14_out(.a(u_csamul_cska32_and4_14[0]), .b(u_csamul_cska32_fa5_13_xor1[0]), .cin(u_csamul_cska32_fa4_13_or0[0]), .fa_xor1(u_csamul_cska32_fa4_14_xor1), .fa_or0(u_csamul_cska32_fa4_14_or0));
  and_gate and_gate_u_csamul_cska32_and5_14(.a(a[5]), .b(b[14]), .out(u_csamul_cska32_and5_14));
  fa fa_u_csamul_cska32_fa5_14_out(.a(u_csamul_cska32_and5_14[0]), .b(u_csamul_cska32_fa6_13_xor1[0]), .cin(u_csamul_cska32_fa5_13_or0[0]), .fa_xor1(u_csamul_cska32_fa5_14_xor1), .fa_or0(u_csamul_cska32_fa5_14_or0));
  and_gate and_gate_u_csamul_cska32_and6_14(.a(a[6]), .b(b[14]), .out(u_csamul_cska32_and6_14));
  fa fa_u_csamul_cska32_fa6_14_out(.a(u_csamul_cska32_and6_14[0]), .b(u_csamul_cska32_fa7_13_xor1[0]), .cin(u_csamul_cska32_fa6_13_or0[0]), .fa_xor1(u_csamul_cska32_fa6_14_xor1), .fa_or0(u_csamul_cska32_fa6_14_or0));
  and_gate and_gate_u_csamul_cska32_and7_14(.a(a[7]), .b(b[14]), .out(u_csamul_cska32_and7_14));
  fa fa_u_csamul_cska32_fa7_14_out(.a(u_csamul_cska32_and7_14[0]), .b(u_csamul_cska32_fa8_13_xor1[0]), .cin(u_csamul_cska32_fa7_13_or0[0]), .fa_xor1(u_csamul_cska32_fa7_14_xor1), .fa_or0(u_csamul_cska32_fa7_14_or0));
  and_gate and_gate_u_csamul_cska32_and8_14(.a(a[8]), .b(b[14]), .out(u_csamul_cska32_and8_14));
  fa fa_u_csamul_cska32_fa8_14_out(.a(u_csamul_cska32_and8_14[0]), .b(u_csamul_cska32_fa9_13_xor1[0]), .cin(u_csamul_cska32_fa8_13_or0[0]), .fa_xor1(u_csamul_cska32_fa8_14_xor1), .fa_or0(u_csamul_cska32_fa8_14_or0));
  and_gate and_gate_u_csamul_cska32_and9_14(.a(a[9]), .b(b[14]), .out(u_csamul_cska32_and9_14));
  fa fa_u_csamul_cska32_fa9_14_out(.a(u_csamul_cska32_and9_14[0]), .b(u_csamul_cska32_fa10_13_xor1[0]), .cin(u_csamul_cska32_fa9_13_or0[0]), .fa_xor1(u_csamul_cska32_fa9_14_xor1), .fa_or0(u_csamul_cska32_fa9_14_or0));
  and_gate and_gate_u_csamul_cska32_and10_14(.a(a[10]), .b(b[14]), .out(u_csamul_cska32_and10_14));
  fa fa_u_csamul_cska32_fa10_14_out(.a(u_csamul_cska32_and10_14[0]), .b(u_csamul_cska32_fa11_13_xor1[0]), .cin(u_csamul_cska32_fa10_13_or0[0]), .fa_xor1(u_csamul_cska32_fa10_14_xor1), .fa_or0(u_csamul_cska32_fa10_14_or0));
  and_gate and_gate_u_csamul_cska32_and11_14(.a(a[11]), .b(b[14]), .out(u_csamul_cska32_and11_14));
  fa fa_u_csamul_cska32_fa11_14_out(.a(u_csamul_cska32_and11_14[0]), .b(u_csamul_cska32_fa12_13_xor1[0]), .cin(u_csamul_cska32_fa11_13_or0[0]), .fa_xor1(u_csamul_cska32_fa11_14_xor1), .fa_or0(u_csamul_cska32_fa11_14_or0));
  and_gate and_gate_u_csamul_cska32_and12_14(.a(a[12]), .b(b[14]), .out(u_csamul_cska32_and12_14));
  fa fa_u_csamul_cska32_fa12_14_out(.a(u_csamul_cska32_and12_14[0]), .b(u_csamul_cska32_fa13_13_xor1[0]), .cin(u_csamul_cska32_fa12_13_or0[0]), .fa_xor1(u_csamul_cska32_fa12_14_xor1), .fa_or0(u_csamul_cska32_fa12_14_or0));
  and_gate and_gate_u_csamul_cska32_and13_14(.a(a[13]), .b(b[14]), .out(u_csamul_cska32_and13_14));
  fa fa_u_csamul_cska32_fa13_14_out(.a(u_csamul_cska32_and13_14[0]), .b(u_csamul_cska32_fa14_13_xor1[0]), .cin(u_csamul_cska32_fa13_13_or0[0]), .fa_xor1(u_csamul_cska32_fa13_14_xor1), .fa_or0(u_csamul_cska32_fa13_14_or0));
  and_gate and_gate_u_csamul_cska32_and14_14(.a(a[14]), .b(b[14]), .out(u_csamul_cska32_and14_14));
  fa fa_u_csamul_cska32_fa14_14_out(.a(u_csamul_cska32_and14_14[0]), .b(u_csamul_cska32_fa15_13_xor1[0]), .cin(u_csamul_cska32_fa14_13_or0[0]), .fa_xor1(u_csamul_cska32_fa14_14_xor1), .fa_or0(u_csamul_cska32_fa14_14_or0));
  and_gate and_gate_u_csamul_cska32_and15_14(.a(a[15]), .b(b[14]), .out(u_csamul_cska32_and15_14));
  fa fa_u_csamul_cska32_fa15_14_out(.a(u_csamul_cska32_and15_14[0]), .b(u_csamul_cska32_fa16_13_xor1[0]), .cin(u_csamul_cska32_fa15_13_or0[0]), .fa_xor1(u_csamul_cska32_fa15_14_xor1), .fa_or0(u_csamul_cska32_fa15_14_or0));
  and_gate and_gate_u_csamul_cska32_and16_14(.a(a[16]), .b(b[14]), .out(u_csamul_cska32_and16_14));
  fa fa_u_csamul_cska32_fa16_14_out(.a(u_csamul_cska32_and16_14[0]), .b(u_csamul_cska32_fa17_13_xor1[0]), .cin(u_csamul_cska32_fa16_13_or0[0]), .fa_xor1(u_csamul_cska32_fa16_14_xor1), .fa_or0(u_csamul_cska32_fa16_14_or0));
  and_gate and_gate_u_csamul_cska32_and17_14(.a(a[17]), .b(b[14]), .out(u_csamul_cska32_and17_14));
  fa fa_u_csamul_cska32_fa17_14_out(.a(u_csamul_cska32_and17_14[0]), .b(u_csamul_cska32_fa18_13_xor1[0]), .cin(u_csamul_cska32_fa17_13_or0[0]), .fa_xor1(u_csamul_cska32_fa17_14_xor1), .fa_or0(u_csamul_cska32_fa17_14_or0));
  and_gate and_gate_u_csamul_cska32_and18_14(.a(a[18]), .b(b[14]), .out(u_csamul_cska32_and18_14));
  fa fa_u_csamul_cska32_fa18_14_out(.a(u_csamul_cska32_and18_14[0]), .b(u_csamul_cska32_fa19_13_xor1[0]), .cin(u_csamul_cska32_fa18_13_or0[0]), .fa_xor1(u_csamul_cska32_fa18_14_xor1), .fa_or0(u_csamul_cska32_fa18_14_or0));
  and_gate and_gate_u_csamul_cska32_and19_14(.a(a[19]), .b(b[14]), .out(u_csamul_cska32_and19_14));
  fa fa_u_csamul_cska32_fa19_14_out(.a(u_csamul_cska32_and19_14[0]), .b(u_csamul_cska32_fa20_13_xor1[0]), .cin(u_csamul_cska32_fa19_13_or0[0]), .fa_xor1(u_csamul_cska32_fa19_14_xor1), .fa_or0(u_csamul_cska32_fa19_14_or0));
  and_gate and_gate_u_csamul_cska32_and20_14(.a(a[20]), .b(b[14]), .out(u_csamul_cska32_and20_14));
  fa fa_u_csamul_cska32_fa20_14_out(.a(u_csamul_cska32_and20_14[0]), .b(u_csamul_cska32_fa21_13_xor1[0]), .cin(u_csamul_cska32_fa20_13_or0[0]), .fa_xor1(u_csamul_cska32_fa20_14_xor1), .fa_or0(u_csamul_cska32_fa20_14_or0));
  and_gate and_gate_u_csamul_cska32_and21_14(.a(a[21]), .b(b[14]), .out(u_csamul_cska32_and21_14));
  fa fa_u_csamul_cska32_fa21_14_out(.a(u_csamul_cska32_and21_14[0]), .b(u_csamul_cska32_fa22_13_xor1[0]), .cin(u_csamul_cska32_fa21_13_or0[0]), .fa_xor1(u_csamul_cska32_fa21_14_xor1), .fa_or0(u_csamul_cska32_fa21_14_or0));
  and_gate and_gate_u_csamul_cska32_and22_14(.a(a[22]), .b(b[14]), .out(u_csamul_cska32_and22_14));
  fa fa_u_csamul_cska32_fa22_14_out(.a(u_csamul_cska32_and22_14[0]), .b(u_csamul_cska32_fa23_13_xor1[0]), .cin(u_csamul_cska32_fa22_13_or0[0]), .fa_xor1(u_csamul_cska32_fa22_14_xor1), .fa_or0(u_csamul_cska32_fa22_14_or0));
  and_gate and_gate_u_csamul_cska32_and23_14(.a(a[23]), .b(b[14]), .out(u_csamul_cska32_and23_14));
  fa fa_u_csamul_cska32_fa23_14_out(.a(u_csamul_cska32_and23_14[0]), .b(u_csamul_cska32_fa24_13_xor1[0]), .cin(u_csamul_cska32_fa23_13_or0[0]), .fa_xor1(u_csamul_cska32_fa23_14_xor1), .fa_or0(u_csamul_cska32_fa23_14_or0));
  and_gate and_gate_u_csamul_cska32_and24_14(.a(a[24]), .b(b[14]), .out(u_csamul_cska32_and24_14));
  fa fa_u_csamul_cska32_fa24_14_out(.a(u_csamul_cska32_and24_14[0]), .b(u_csamul_cska32_fa25_13_xor1[0]), .cin(u_csamul_cska32_fa24_13_or0[0]), .fa_xor1(u_csamul_cska32_fa24_14_xor1), .fa_or0(u_csamul_cska32_fa24_14_or0));
  and_gate and_gate_u_csamul_cska32_and25_14(.a(a[25]), .b(b[14]), .out(u_csamul_cska32_and25_14));
  fa fa_u_csamul_cska32_fa25_14_out(.a(u_csamul_cska32_and25_14[0]), .b(u_csamul_cska32_fa26_13_xor1[0]), .cin(u_csamul_cska32_fa25_13_or0[0]), .fa_xor1(u_csamul_cska32_fa25_14_xor1), .fa_or0(u_csamul_cska32_fa25_14_or0));
  and_gate and_gate_u_csamul_cska32_and26_14(.a(a[26]), .b(b[14]), .out(u_csamul_cska32_and26_14));
  fa fa_u_csamul_cska32_fa26_14_out(.a(u_csamul_cska32_and26_14[0]), .b(u_csamul_cska32_fa27_13_xor1[0]), .cin(u_csamul_cska32_fa26_13_or0[0]), .fa_xor1(u_csamul_cska32_fa26_14_xor1), .fa_or0(u_csamul_cska32_fa26_14_or0));
  and_gate and_gate_u_csamul_cska32_and27_14(.a(a[27]), .b(b[14]), .out(u_csamul_cska32_and27_14));
  fa fa_u_csamul_cska32_fa27_14_out(.a(u_csamul_cska32_and27_14[0]), .b(u_csamul_cska32_fa28_13_xor1[0]), .cin(u_csamul_cska32_fa27_13_or0[0]), .fa_xor1(u_csamul_cska32_fa27_14_xor1), .fa_or0(u_csamul_cska32_fa27_14_or0));
  and_gate and_gate_u_csamul_cska32_and28_14(.a(a[28]), .b(b[14]), .out(u_csamul_cska32_and28_14));
  fa fa_u_csamul_cska32_fa28_14_out(.a(u_csamul_cska32_and28_14[0]), .b(u_csamul_cska32_fa29_13_xor1[0]), .cin(u_csamul_cska32_fa28_13_or0[0]), .fa_xor1(u_csamul_cska32_fa28_14_xor1), .fa_or0(u_csamul_cska32_fa28_14_or0));
  and_gate and_gate_u_csamul_cska32_and29_14(.a(a[29]), .b(b[14]), .out(u_csamul_cska32_and29_14));
  fa fa_u_csamul_cska32_fa29_14_out(.a(u_csamul_cska32_and29_14[0]), .b(u_csamul_cska32_fa30_13_xor1[0]), .cin(u_csamul_cska32_fa29_13_or0[0]), .fa_xor1(u_csamul_cska32_fa29_14_xor1), .fa_or0(u_csamul_cska32_fa29_14_or0));
  and_gate and_gate_u_csamul_cska32_and30_14(.a(a[30]), .b(b[14]), .out(u_csamul_cska32_and30_14));
  fa fa_u_csamul_cska32_fa30_14_out(.a(u_csamul_cska32_and30_14[0]), .b(u_csamul_cska32_and31_13[0]), .cin(u_csamul_cska32_fa30_13_or0[0]), .fa_xor1(u_csamul_cska32_fa30_14_xor1), .fa_or0(u_csamul_cska32_fa30_14_or0));
  and_gate and_gate_u_csamul_cska32_and31_14(.a(a[31]), .b(b[14]), .out(u_csamul_cska32_and31_14));
  and_gate and_gate_u_csamul_cska32_and0_15(.a(a[0]), .b(b[15]), .out(u_csamul_cska32_and0_15));
  fa fa_u_csamul_cska32_fa0_15_out(.a(u_csamul_cska32_and0_15[0]), .b(u_csamul_cska32_fa1_14_xor1[0]), .cin(u_csamul_cska32_fa0_14_or0[0]), .fa_xor1(u_csamul_cska32_fa0_15_xor1), .fa_or0(u_csamul_cska32_fa0_15_or0));
  and_gate and_gate_u_csamul_cska32_and1_15(.a(a[1]), .b(b[15]), .out(u_csamul_cska32_and1_15));
  fa fa_u_csamul_cska32_fa1_15_out(.a(u_csamul_cska32_and1_15[0]), .b(u_csamul_cska32_fa2_14_xor1[0]), .cin(u_csamul_cska32_fa1_14_or0[0]), .fa_xor1(u_csamul_cska32_fa1_15_xor1), .fa_or0(u_csamul_cska32_fa1_15_or0));
  and_gate and_gate_u_csamul_cska32_and2_15(.a(a[2]), .b(b[15]), .out(u_csamul_cska32_and2_15));
  fa fa_u_csamul_cska32_fa2_15_out(.a(u_csamul_cska32_and2_15[0]), .b(u_csamul_cska32_fa3_14_xor1[0]), .cin(u_csamul_cska32_fa2_14_or0[0]), .fa_xor1(u_csamul_cska32_fa2_15_xor1), .fa_or0(u_csamul_cska32_fa2_15_or0));
  and_gate and_gate_u_csamul_cska32_and3_15(.a(a[3]), .b(b[15]), .out(u_csamul_cska32_and3_15));
  fa fa_u_csamul_cska32_fa3_15_out(.a(u_csamul_cska32_and3_15[0]), .b(u_csamul_cska32_fa4_14_xor1[0]), .cin(u_csamul_cska32_fa3_14_or0[0]), .fa_xor1(u_csamul_cska32_fa3_15_xor1), .fa_or0(u_csamul_cska32_fa3_15_or0));
  and_gate and_gate_u_csamul_cska32_and4_15(.a(a[4]), .b(b[15]), .out(u_csamul_cska32_and4_15));
  fa fa_u_csamul_cska32_fa4_15_out(.a(u_csamul_cska32_and4_15[0]), .b(u_csamul_cska32_fa5_14_xor1[0]), .cin(u_csamul_cska32_fa4_14_or0[0]), .fa_xor1(u_csamul_cska32_fa4_15_xor1), .fa_or0(u_csamul_cska32_fa4_15_or0));
  and_gate and_gate_u_csamul_cska32_and5_15(.a(a[5]), .b(b[15]), .out(u_csamul_cska32_and5_15));
  fa fa_u_csamul_cska32_fa5_15_out(.a(u_csamul_cska32_and5_15[0]), .b(u_csamul_cska32_fa6_14_xor1[0]), .cin(u_csamul_cska32_fa5_14_or0[0]), .fa_xor1(u_csamul_cska32_fa5_15_xor1), .fa_or0(u_csamul_cska32_fa5_15_or0));
  and_gate and_gate_u_csamul_cska32_and6_15(.a(a[6]), .b(b[15]), .out(u_csamul_cska32_and6_15));
  fa fa_u_csamul_cska32_fa6_15_out(.a(u_csamul_cska32_and6_15[0]), .b(u_csamul_cska32_fa7_14_xor1[0]), .cin(u_csamul_cska32_fa6_14_or0[0]), .fa_xor1(u_csamul_cska32_fa6_15_xor1), .fa_or0(u_csamul_cska32_fa6_15_or0));
  and_gate and_gate_u_csamul_cska32_and7_15(.a(a[7]), .b(b[15]), .out(u_csamul_cska32_and7_15));
  fa fa_u_csamul_cska32_fa7_15_out(.a(u_csamul_cska32_and7_15[0]), .b(u_csamul_cska32_fa8_14_xor1[0]), .cin(u_csamul_cska32_fa7_14_or0[0]), .fa_xor1(u_csamul_cska32_fa7_15_xor1), .fa_or0(u_csamul_cska32_fa7_15_or0));
  and_gate and_gate_u_csamul_cska32_and8_15(.a(a[8]), .b(b[15]), .out(u_csamul_cska32_and8_15));
  fa fa_u_csamul_cska32_fa8_15_out(.a(u_csamul_cska32_and8_15[0]), .b(u_csamul_cska32_fa9_14_xor1[0]), .cin(u_csamul_cska32_fa8_14_or0[0]), .fa_xor1(u_csamul_cska32_fa8_15_xor1), .fa_or0(u_csamul_cska32_fa8_15_or0));
  and_gate and_gate_u_csamul_cska32_and9_15(.a(a[9]), .b(b[15]), .out(u_csamul_cska32_and9_15));
  fa fa_u_csamul_cska32_fa9_15_out(.a(u_csamul_cska32_and9_15[0]), .b(u_csamul_cska32_fa10_14_xor1[0]), .cin(u_csamul_cska32_fa9_14_or0[0]), .fa_xor1(u_csamul_cska32_fa9_15_xor1), .fa_or0(u_csamul_cska32_fa9_15_or0));
  and_gate and_gate_u_csamul_cska32_and10_15(.a(a[10]), .b(b[15]), .out(u_csamul_cska32_and10_15));
  fa fa_u_csamul_cska32_fa10_15_out(.a(u_csamul_cska32_and10_15[0]), .b(u_csamul_cska32_fa11_14_xor1[0]), .cin(u_csamul_cska32_fa10_14_or0[0]), .fa_xor1(u_csamul_cska32_fa10_15_xor1), .fa_or0(u_csamul_cska32_fa10_15_or0));
  and_gate and_gate_u_csamul_cska32_and11_15(.a(a[11]), .b(b[15]), .out(u_csamul_cska32_and11_15));
  fa fa_u_csamul_cska32_fa11_15_out(.a(u_csamul_cska32_and11_15[0]), .b(u_csamul_cska32_fa12_14_xor1[0]), .cin(u_csamul_cska32_fa11_14_or0[0]), .fa_xor1(u_csamul_cska32_fa11_15_xor1), .fa_or0(u_csamul_cska32_fa11_15_or0));
  and_gate and_gate_u_csamul_cska32_and12_15(.a(a[12]), .b(b[15]), .out(u_csamul_cska32_and12_15));
  fa fa_u_csamul_cska32_fa12_15_out(.a(u_csamul_cska32_and12_15[0]), .b(u_csamul_cska32_fa13_14_xor1[0]), .cin(u_csamul_cska32_fa12_14_or0[0]), .fa_xor1(u_csamul_cska32_fa12_15_xor1), .fa_or0(u_csamul_cska32_fa12_15_or0));
  and_gate and_gate_u_csamul_cska32_and13_15(.a(a[13]), .b(b[15]), .out(u_csamul_cska32_and13_15));
  fa fa_u_csamul_cska32_fa13_15_out(.a(u_csamul_cska32_and13_15[0]), .b(u_csamul_cska32_fa14_14_xor1[0]), .cin(u_csamul_cska32_fa13_14_or0[0]), .fa_xor1(u_csamul_cska32_fa13_15_xor1), .fa_or0(u_csamul_cska32_fa13_15_or0));
  and_gate and_gate_u_csamul_cska32_and14_15(.a(a[14]), .b(b[15]), .out(u_csamul_cska32_and14_15));
  fa fa_u_csamul_cska32_fa14_15_out(.a(u_csamul_cska32_and14_15[0]), .b(u_csamul_cska32_fa15_14_xor1[0]), .cin(u_csamul_cska32_fa14_14_or0[0]), .fa_xor1(u_csamul_cska32_fa14_15_xor1), .fa_or0(u_csamul_cska32_fa14_15_or0));
  and_gate and_gate_u_csamul_cska32_and15_15(.a(a[15]), .b(b[15]), .out(u_csamul_cska32_and15_15));
  fa fa_u_csamul_cska32_fa15_15_out(.a(u_csamul_cska32_and15_15[0]), .b(u_csamul_cska32_fa16_14_xor1[0]), .cin(u_csamul_cska32_fa15_14_or0[0]), .fa_xor1(u_csamul_cska32_fa15_15_xor1), .fa_or0(u_csamul_cska32_fa15_15_or0));
  and_gate and_gate_u_csamul_cska32_and16_15(.a(a[16]), .b(b[15]), .out(u_csamul_cska32_and16_15));
  fa fa_u_csamul_cska32_fa16_15_out(.a(u_csamul_cska32_and16_15[0]), .b(u_csamul_cska32_fa17_14_xor1[0]), .cin(u_csamul_cska32_fa16_14_or0[0]), .fa_xor1(u_csamul_cska32_fa16_15_xor1), .fa_or0(u_csamul_cska32_fa16_15_or0));
  and_gate and_gate_u_csamul_cska32_and17_15(.a(a[17]), .b(b[15]), .out(u_csamul_cska32_and17_15));
  fa fa_u_csamul_cska32_fa17_15_out(.a(u_csamul_cska32_and17_15[0]), .b(u_csamul_cska32_fa18_14_xor1[0]), .cin(u_csamul_cska32_fa17_14_or0[0]), .fa_xor1(u_csamul_cska32_fa17_15_xor1), .fa_or0(u_csamul_cska32_fa17_15_or0));
  and_gate and_gate_u_csamul_cska32_and18_15(.a(a[18]), .b(b[15]), .out(u_csamul_cska32_and18_15));
  fa fa_u_csamul_cska32_fa18_15_out(.a(u_csamul_cska32_and18_15[0]), .b(u_csamul_cska32_fa19_14_xor1[0]), .cin(u_csamul_cska32_fa18_14_or0[0]), .fa_xor1(u_csamul_cska32_fa18_15_xor1), .fa_or0(u_csamul_cska32_fa18_15_or0));
  and_gate and_gate_u_csamul_cska32_and19_15(.a(a[19]), .b(b[15]), .out(u_csamul_cska32_and19_15));
  fa fa_u_csamul_cska32_fa19_15_out(.a(u_csamul_cska32_and19_15[0]), .b(u_csamul_cska32_fa20_14_xor1[0]), .cin(u_csamul_cska32_fa19_14_or0[0]), .fa_xor1(u_csamul_cska32_fa19_15_xor1), .fa_or0(u_csamul_cska32_fa19_15_or0));
  and_gate and_gate_u_csamul_cska32_and20_15(.a(a[20]), .b(b[15]), .out(u_csamul_cska32_and20_15));
  fa fa_u_csamul_cska32_fa20_15_out(.a(u_csamul_cska32_and20_15[0]), .b(u_csamul_cska32_fa21_14_xor1[0]), .cin(u_csamul_cska32_fa20_14_or0[0]), .fa_xor1(u_csamul_cska32_fa20_15_xor1), .fa_or0(u_csamul_cska32_fa20_15_or0));
  and_gate and_gate_u_csamul_cska32_and21_15(.a(a[21]), .b(b[15]), .out(u_csamul_cska32_and21_15));
  fa fa_u_csamul_cska32_fa21_15_out(.a(u_csamul_cska32_and21_15[0]), .b(u_csamul_cska32_fa22_14_xor1[0]), .cin(u_csamul_cska32_fa21_14_or0[0]), .fa_xor1(u_csamul_cska32_fa21_15_xor1), .fa_or0(u_csamul_cska32_fa21_15_or0));
  and_gate and_gate_u_csamul_cska32_and22_15(.a(a[22]), .b(b[15]), .out(u_csamul_cska32_and22_15));
  fa fa_u_csamul_cska32_fa22_15_out(.a(u_csamul_cska32_and22_15[0]), .b(u_csamul_cska32_fa23_14_xor1[0]), .cin(u_csamul_cska32_fa22_14_or0[0]), .fa_xor1(u_csamul_cska32_fa22_15_xor1), .fa_or0(u_csamul_cska32_fa22_15_or0));
  and_gate and_gate_u_csamul_cska32_and23_15(.a(a[23]), .b(b[15]), .out(u_csamul_cska32_and23_15));
  fa fa_u_csamul_cska32_fa23_15_out(.a(u_csamul_cska32_and23_15[0]), .b(u_csamul_cska32_fa24_14_xor1[0]), .cin(u_csamul_cska32_fa23_14_or0[0]), .fa_xor1(u_csamul_cska32_fa23_15_xor1), .fa_or0(u_csamul_cska32_fa23_15_or0));
  and_gate and_gate_u_csamul_cska32_and24_15(.a(a[24]), .b(b[15]), .out(u_csamul_cska32_and24_15));
  fa fa_u_csamul_cska32_fa24_15_out(.a(u_csamul_cska32_and24_15[0]), .b(u_csamul_cska32_fa25_14_xor1[0]), .cin(u_csamul_cska32_fa24_14_or0[0]), .fa_xor1(u_csamul_cska32_fa24_15_xor1), .fa_or0(u_csamul_cska32_fa24_15_or0));
  and_gate and_gate_u_csamul_cska32_and25_15(.a(a[25]), .b(b[15]), .out(u_csamul_cska32_and25_15));
  fa fa_u_csamul_cska32_fa25_15_out(.a(u_csamul_cska32_and25_15[0]), .b(u_csamul_cska32_fa26_14_xor1[0]), .cin(u_csamul_cska32_fa25_14_or0[0]), .fa_xor1(u_csamul_cska32_fa25_15_xor1), .fa_or0(u_csamul_cska32_fa25_15_or0));
  and_gate and_gate_u_csamul_cska32_and26_15(.a(a[26]), .b(b[15]), .out(u_csamul_cska32_and26_15));
  fa fa_u_csamul_cska32_fa26_15_out(.a(u_csamul_cska32_and26_15[0]), .b(u_csamul_cska32_fa27_14_xor1[0]), .cin(u_csamul_cska32_fa26_14_or0[0]), .fa_xor1(u_csamul_cska32_fa26_15_xor1), .fa_or0(u_csamul_cska32_fa26_15_or0));
  and_gate and_gate_u_csamul_cska32_and27_15(.a(a[27]), .b(b[15]), .out(u_csamul_cska32_and27_15));
  fa fa_u_csamul_cska32_fa27_15_out(.a(u_csamul_cska32_and27_15[0]), .b(u_csamul_cska32_fa28_14_xor1[0]), .cin(u_csamul_cska32_fa27_14_or0[0]), .fa_xor1(u_csamul_cska32_fa27_15_xor1), .fa_or0(u_csamul_cska32_fa27_15_or0));
  and_gate and_gate_u_csamul_cska32_and28_15(.a(a[28]), .b(b[15]), .out(u_csamul_cska32_and28_15));
  fa fa_u_csamul_cska32_fa28_15_out(.a(u_csamul_cska32_and28_15[0]), .b(u_csamul_cska32_fa29_14_xor1[0]), .cin(u_csamul_cska32_fa28_14_or0[0]), .fa_xor1(u_csamul_cska32_fa28_15_xor1), .fa_or0(u_csamul_cska32_fa28_15_or0));
  and_gate and_gate_u_csamul_cska32_and29_15(.a(a[29]), .b(b[15]), .out(u_csamul_cska32_and29_15));
  fa fa_u_csamul_cska32_fa29_15_out(.a(u_csamul_cska32_and29_15[0]), .b(u_csamul_cska32_fa30_14_xor1[0]), .cin(u_csamul_cska32_fa29_14_or0[0]), .fa_xor1(u_csamul_cska32_fa29_15_xor1), .fa_or0(u_csamul_cska32_fa29_15_or0));
  and_gate and_gate_u_csamul_cska32_and30_15(.a(a[30]), .b(b[15]), .out(u_csamul_cska32_and30_15));
  fa fa_u_csamul_cska32_fa30_15_out(.a(u_csamul_cska32_and30_15[0]), .b(u_csamul_cska32_and31_14[0]), .cin(u_csamul_cska32_fa30_14_or0[0]), .fa_xor1(u_csamul_cska32_fa30_15_xor1), .fa_or0(u_csamul_cska32_fa30_15_or0));
  and_gate and_gate_u_csamul_cska32_and31_15(.a(a[31]), .b(b[15]), .out(u_csamul_cska32_and31_15));
  and_gate and_gate_u_csamul_cska32_and0_16(.a(a[0]), .b(b[16]), .out(u_csamul_cska32_and0_16));
  fa fa_u_csamul_cska32_fa0_16_out(.a(u_csamul_cska32_and0_16[0]), .b(u_csamul_cska32_fa1_15_xor1[0]), .cin(u_csamul_cska32_fa0_15_or0[0]), .fa_xor1(u_csamul_cska32_fa0_16_xor1), .fa_or0(u_csamul_cska32_fa0_16_or0));
  and_gate and_gate_u_csamul_cska32_and1_16(.a(a[1]), .b(b[16]), .out(u_csamul_cska32_and1_16));
  fa fa_u_csamul_cska32_fa1_16_out(.a(u_csamul_cska32_and1_16[0]), .b(u_csamul_cska32_fa2_15_xor1[0]), .cin(u_csamul_cska32_fa1_15_or0[0]), .fa_xor1(u_csamul_cska32_fa1_16_xor1), .fa_or0(u_csamul_cska32_fa1_16_or0));
  and_gate and_gate_u_csamul_cska32_and2_16(.a(a[2]), .b(b[16]), .out(u_csamul_cska32_and2_16));
  fa fa_u_csamul_cska32_fa2_16_out(.a(u_csamul_cska32_and2_16[0]), .b(u_csamul_cska32_fa3_15_xor1[0]), .cin(u_csamul_cska32_fa2_15_or0[0]), .fa_xor1(u_csamul_cska32_fa2_16_xor1), .fa_or0(u_csamul_cska32_fa2_16_or0));
  and_gate and_gate_u_csamul_cska32_and3_16(.a(a[3]), .b(b[16]), .out(u_csamul_cska32_and3_16));
  fa fa_u_csamul_cska32_fa3_16_out(.a(u_csamul_cska32_and3_16[0]), .b(u_csamul_cska32_fa4_15_xor1[0]), .cin(u_csamul_cska32_fa3_15_or0[0]), .fa_xor1(u_csamul_cska32_fa3_16_xor1), .fa_or0(u_csamul_cska32_fa3_16_or0));
  and_gate and_gate_u_csamul_cska32_and4_16(.a(a[4]), .b(b[16]), .out(u_csamul_cska32_and4_16));
  fa fa_u_csamul_cska32_fa4_16_out(.a(u_csamul_cska32_and4_16[0]), .b(u_csamul_cska32_fa5_15_xor1[0]), .cin(u_csamul_cska32_fa4_15_or0[0]), .fa_xor1(u_csamul_cska32_fa4_16_xor1), .fa_or0(u_csamul_cska32_fa4_16_or0));
  and_gate and_gate_u_csamul_cska32_and5_16(.a(a[5]), .b(b[16]), .out(u_csamul_cska32_and5_16));
  fa fa_u_csamul_cska32_fa5_16_out(.a(u_csamul_cska32_and5_16[0]), .b(u_csamul_cska32_fa6_15_xor1[0]), .cin(u_csamul_cska32_fa5_15_or0[0]), .fa_xor1(u_csamul_cska32_fa5_16_xor1), .fa_or0(u_csamul_cska32_fa5_16_or0));
  and_gate and_gate_u_csamul_cska32_and6_16(.a(a[6]), .b(b[16]), .out(u_csamul_cska32_and6_16));
  fa fa_u_csamul_cska32_fa6_16_out(.a(u_csamul_cska32_and6_16[0]), .b(u_csamul_cska32_fa7_15_xor1[0]), .cin(u_csamul_cska32_fa6_15_or0[0]), .fa_xor1(u_csamul_cska32_fa6_16_xor1), .fa_or0(u_csamul_cska32_fa6_16_or0));
  and_gate and_gate_u_csamul_cska32_and7_16(.a(a[7]), .b(b[16]), .out(u_csamul_cska32_and7_16));
  fa fa_u_csamul_cska32_fa7_16_out(.a(u_csamul_cska32_and7_16[0]), .b(u_csamul_cska32_fa8_15_xor1[0]), .cin(u_csamul_cska32_fa7_15_or0[0]), .fa_xor1(u_csamul_cska32_fa7_16_xor1), .fa_or0(u_csamul_cska32_fa7_16_or0));
  and_gate and_gate_u_csamul_cska32_and8_16(.a(a[8]), .b(b[16]), .out(u_csamul_cska32_and8_16));
  fa fa_u_csamul_cska32_fa8_16_out(.a(u_csamul_cska32_and8_16[0]), .b(u_csamul_cska32_fa9_15_xor1[0]), .cin(u_csamul_cska32_fa8_15_or0[0]), .fa_xor1(u_csamul_cska32_fa8_16_xor1), .fa_or0(u_csamul_cska32_fa8_16_or0));
  and_gate and_gate_u_csamul_cska32_and9_16(.a(a[9]), .b(b[16]), .out(u_csamul_cska32_and9_16));
  fa fa_u_csamul_cska32_fa9_16_out(.a(u_csamul_cska32_and9_16[0]), .b(u_csamul_cska32_fa10_15_xor1[0]), .cin(u_csamul_cska32_fa9_15_or0[0]), .fa_xor1(u_csamul_cska32_fa9_16_xor1), .fa_or0(u_csamul_cska32_fa9_16_or0));
  and_gate and_gate_u_csamul_cska32_and10_16(.a(a[10]), .b(b[16]), .out(u_csamul_cska32_and10_16));
  fa fa_u_csamul_cska32_fa10_16_out(.a(u_csamul_cska32_and10_16[0]), .b(u_csamul_cska32_fa11_15_xor1[0]), .cin(u_csamul_cska32_fa10_15_or0[0]), .fa_xor1(u_csamul_cska32_fa10_16_xor1), .fa_or0(u_csamul_cska32_fa10_16_or0));
  and_gate and_gate_u_csamul_cska32_and11_16(.a(a[11]), .b(b[16]), .out(u_csamul_cska32_and11_16));
  fa fa_u_csamul_cska32_fa11_16_out(.a(u_csamul_cska32_and11_16[0]), .b(u_csamul_cska32_fa12_15_xor1[0]), .cin(u_csamul_cska32_fa11_15_or0[0]), .fa_xor1(u_csamul_cska32_fa11_16_xor1), .fa_or0(u_csamul_cska32_fa11_16_or0));
  and_gate and_gate_u_csamul_cska32_and12_16(.a(a[12]), .b(b[16]), .out(u_csamul_cska32_and12_16));
  fa fa_u_csamul_cska32_fa12_16_out(.a(u_csamul_cska32_and12_16[0]), .b(u_csamul_cska32_fa13_15_xor1[0]), .cin(u_csamul_cska32_fa12_15_or0[0]), .fa_xor1(u_csamul_cska32_fa12_16_xor1), .fa_or0(u_csamul_cska32_fa12_16_or0));
  and_gate and_gate_u_csamul_cska32_and13_16(.a(a[13]), .b(b[16]), .out(u_csamul_cska32_and13_16));
  fa fa_u_csamul_cska32_fa13_16_out(.a(u_csamul_cska32_and13_16[0]), .b(u_csamul_cska32_fa14_15_xor1[0]), .cin(u_csamul_cska32_fa13_15_or0[0]), .fa_xor1(u_csamul_cska32_fa13_16_xor1), .fa_or0(u_csamul_cska32_fa13_16_or0));
  and_gate and_gate_u_csamul_cska32_and14_16(.a(a[14]), .b(b[16]), .out(u_csamul_cska32_and14_16));
  fa fa_u_csamul_cska32_fa14_16_out(.a(u_csamul_cska32_and14_16[0]), .b(u_csamul_cska32_fa15_15_xor1[0]), .cin(u_csamul_cska32_fa14_15_or0[0]), .fa_xor1(u_csamul_cska32_fa14_16_xor1), .fa_or0(u_csamul_cska32_fa14_16_or0));
  and_gate and_gate_u_csamul_cska32_and15_16(.a(a[15]), .b(b[16]), .out(u_csamul_cska32_and15_16));
  fa fa_u_csamul_cska32_fa15_16_out(.a(u_csamul_cska32_and15_16[0]), .b(u_csamul_cska32_fa16_15_xor1[0]), .cin(u_csamul_cska32_fa15_15_or0[0]), .fa_xor1(u_csamul_cska32_fa15_16_xor1), .fa_or0(u_csamul_cska32_fa15_16_or0));
  and_gate and_gate_u_csamul_cska32_and16_16(.a(a[16]), .b(b[16]), .out(u_csamul_cska32_and16_16));
  fa fa_u_csamul_cska32_fa16_16_out(.a(u_csamul_cska32_and16_16[0]), .b(u_csamul_cska32_fa17_15_xor1[0]), .cin(u_csamul_cska32_fa16_15_or0[0]), .fa_xor1(u_csamul_cska32_fa16_16_xor1), .fa_or0(u_csamul_cska32_fa16_16_or0));
  and_gate and_gate_u_csamul_cska32_and17_16(.a(a[17]), .b(b[16]), .out(u_csamul_cska32_and17_16));
  fa fa_u_csamul_cska32_fa17_16_out(.a(u_csamul_cska32_and17_16[0]), .b(u_csamul_cska32_fa18_15_xor1[0]), .cin(u_csamul_cska32_fa17_15_or0[0]), .fa_xor1(u_csamul_cska32_fa17_16_xor1), .fa_or0(u_csamul_cska32_fa17_16_or0));
  and_gate and_gate_u_csamul_cska32_and18_16(.a(a[18]), .b(b[16]), .out(u_csamul_cska32_and18_16));
  fa fa_u_csamul_cska32_fa18_16_out(.a(u_csamul_cska32_and18_16[0]), .b(u_csamul_cska32_fa19_15_xor1[0]), .cin(u_csamul_cska32_fa18_15_or0[0]), .fa_xor1(u_csamul_cska32_fa18_16_xor1), .fa_or0(u_csamul_cska32_fa18_16_or0));
  and_gate and_gate_u_csamul_cska32_and19_16(.a(a[19]), .b(b[16]), .out(u_csamul_cska32_and19_16));
  fa fa_u_csamul_cska32_fa19_16_out(.a(u_csamul_cska32_and19_16[0]), .b(u_csamul_cska32_fa20_15_xor1[0]), .cin(u_csamul_cska32_fa19_15_or0[0]), .fa_xor1(u_csamul_cska32_fa19_16_xor1), .fa_or0(u_csamul_cska32_fa19_16_or0));
  and_gate and_gate_u_csamul_cska32_and20_16(.a(a[20]), .b(b[16]), .out(u_csamul_cska32_and20_16));
  fa fa_u_csamul_cska32_fa20_16_out(.a(u_csamul_cska32_and20_16[0]), .b(u_csamul_cska32_fa21_15_xor1[0]), .cin(u_csamul_cska32_fa20_15_or0[0]), .fa_xor1(u_csamul_cska32_fa20_16_xor1), .fa_or0(u_csamul_cska32_fa20_16_or0));
  and_gate and_gate_u_csamul_cska32_and21_16(.a(a[21]), .b(b[16]), .out(u_csamul_cska32_and21_16));
  fa fa_u_csamul_cska32_fa21_16_out(.a(u_csamul_cska32_and21_16[0]), .b(u_csamul_cska32_fa22_15_xor1[0]), .cin(u_csamul_cska32_fa21_15_or0[0]), .fa_xor1(u_csamul_cska32_fa21_16_xor1), .fa_or0(u_csamul_cska32_fa21_16_or0));
  and_gate and_gate_u_csamul_cska32_and22_16(.a(a[22]), .b(b[16]), .out(u_csamul_cska32_and22_16));
  fa fa_u_csamul_cska32_fa22_16_out(.a(u_csamul_cska32_and22_16[0]), .b(u_csamul_cska32_fa23_15_xor1[0]), .cin(u_csamul_cska32_fa22_15_or0[0]), .fa_xor1(u_csamul_cska32_fa22_16_xor1), .fa_or0(u_csamul_cska32_fa22_16_or0));
  and_gate and_gate_u_csamul_cska32_and23_16(.a(a[23]), .b(b[16]), .out(u_csamul_cska32_and23_16));
  fa fa_u_csamul_cska32_fa23_16_out(.a(u_csamul_cska32_and23_16[0]), .b(u_csamul_cska32_fa24_15_xor1[0]), .cin(u_csamul_cska32_fa23_15_or0[0]), .fa_xor1(u_csamul_cska32_fa23_16_xor1), .fa_or0(u_csamul_cska32_fa23_16_or0));
  and_gate and_gate_u_csamul_cska32_and24_16(.a(a[24]), .b(b[16]), .out(u_csamul_cska32_and24_16));
  fa fa_u_csamul_cska32_fa24_16_out(.a(u_csamul_cska32_and24_16[0]), .b(u_csamul_cska32_fa25_15_xor1[0]), .cin(u_csamul_cska32_fa24_15_or0[0]), .fa_xor1(u_csamul_cska32_fa24_16_xor1), .fa_or0(u_csamul_cska32_fa24_16_or0));
  and_gate and_gate_u_csamul_cska32_and25_16(.a(a[25]), .b(b[16]), .out(u_csamul_cska32_and25_16));
  fa fa_u_csamul_cska32_fa25_16_out(.a(u_csamul_cska32_and25_16[0]), .b(u_csamul_cska32_fa26_15_xor1[0]), .cin(u_csamul_cska32_fa25_15_or0[0]), .fa_xor1(u_csamul_cska32_fa25_16_xor1), .fa_or0(u_csamul_cska32_fa25_16_or0));
  and_gate and_gate_u_csamul_cska32_and26_16(.a(a[26]), .b(b[16]), .out(u_csamul_cska32_and26_16));
  fa fa_u_csamul_cska32_fa26_16_out(.a(u_csamul_cska32_and26_16[0]), .b(u_csamul_cska32_fa27_15_xor1[0]), .cin(u_csamul_cska32_fa26_15_or0[0]), .fa_xor1(u_csamul_cska32_fa26_16_xor1), .fa_or0(u_csamul_cska32_fa26_16_or0));
  and_gate and_gate_u_csamul_cska32_and27_16(.a(a[27]), .b(b[16]), .out(u_csamul_cska32_and27_16));
  fa fa_u_csamul_cska32_fa27_16_out(.a(u_csamul_cska32_and27_16[0]), .b(u_csamul_cska32_fa28_15_xor1[0]), .cin(u_csamul_cska32_fa27_15_or0[0]), .fa_xor1(u_csamul_cska32_fa27_16_xor1), .fa_or0(u_csamul_cska32_fa27_16_or0));
  and_gate and_gate_u_csamul_cska32_and28_16(.a(a[28]), .b(b[16]), .out(u_csamul_cska32_and28_16));
  fa fa_u_csamul_cska32_fa28_16_out(.a(u_csamul_cska32_and28_16[0]), .b(u_csamul_cska32_fa29_15_xor1[0]), .cin(u_csamul_cska32_fa28_15_or0[0]), .fa_xor1(u_csamul_cska32_fa28_16_xor1), .fa_or0(u_csamul_cska32_fa28_16_or0));
  and_gate and_gate_u_csamul_cska32_and29_16(.a(a[29]), .b(b[16]), .out(u_csamul_cska32_and29_16));
  fa fa_u_csamul_cska32_fa29_16_out(.a(u_csamul_cska32_and29_16[0]), .b(u_csamul_cska32_fa30_15_xor1[0]), .cin(u_csamul_cska32_fa29_15_or0[0]), .fa_xor1(u_csamul_cska32_fa29_16_xor1), .fa_or0(u_csamul_cska32_fa29_16_or0));
  and_gate and_gate_u_csamul_cska32_and30_16(.a(a[30]), .b(b[16]), .out(u_csamul_cska32_and30_16));
  fa fa_u_csamul_cska32_fa30_16_out(.a(u_csamul_cska32_and30_16[0]), .b(u_csamul_cska32_and31_15[0]), .cin(u_csamul_cska32_fa30_15_or0[0]), .fa_xor1(u_csamul_cska32_fa30_16_xor1), .fa_or0(u_csamul_cska32_fa30_16_or0));
  and_gate and_gate_u_csamul_cska32_and31_16(.a(a[31]), .b(b[16]), .out(u_csamul_cska32_and31_16));
  and_gate and_gate_u_csamul_cska32_and0_17(.a(a[0]), .b(b[17]), .out(u_csamul_cska32_and0_17));
  fa fa_u_csamul_cska32_fa0_17_out(.a(u_csamul_cska32_and0_17[0]), .b(u_csamul_cska32_fa1_16_xor1[0]), .cin(u_csamul_cska32_fa0_16_or0[0]), .fa_xor1(u_csamul_cska32_fa0_17_xor1), .fa_or0(u_csamul_cska32_fa0_17_or0));
  and_gate and_gate_u_csamul_cska32_and1_17(.a(a[1]), .b(b[17]), .out(u_csamul_cska32_and1_17));
  fa fa_u_csamul_cska32_fa1_17_out(.a(u_csamul_cska32_and1_17[0]), .b(u_csamul_cska32_fa2_16_xor1[0]), .cin(u_csamul_cska32_fa1_16_or0[0]), .fa_xor1(u_csamul_cska32_fa1_17_xor1), .fa_or0(u_csamul_cska32_fa1_17_or0));
  and_gate and_gate_u_csamul_cska32_and2_17(.a(a[2]), .b(b[17]), .out(u_csamul_cska32_and2_17));
  fa fa_u_csamul_cska32_fa2_17_out(.a(u_csamul_cska32_and2_17[0]), .b(u_csamul_cska32_fa3_16_xor1[0]), .cin(u_csamul_cska32_fa2_16_or0[0]), .fa_xor1(u_csamul_cska32_fa2_17_xor1), .fa_or0(u_csamul_cska32_fa2_17_or0));
  and_gate and_gate_u_csamul_cska32_and3_17(.a(a[3]), .b(b[17]), .out(u_csamul_cska32_and3_17));
  fa fa_u_csamul_cska32_fa3_17_out(.a(u_csamul_cska32_and3_17[0]), .b(u_csamul_cska32_fa4_16_xor1[0]), .cin(u_csamul_cska32_fa3_16_or0[0]), .fa_xor1(u_csamul_cska32_fa3_17_xor1), .fa_or0(u_csamul_cska32_fa3_17_or0));
  and_gate and_gate_u_csamul_cska32_and4_17(.a(a[4]), .b(b[17]), .out(u_csamul_cska32_and4_17));
  fa fa_u_csamul_cska32_fa4_17_out(.a(u_csamul_cska32_and4_17[0]), .b(u_csamul_cska32_fa5_16_xor1[0]), .cin(u_csamul_cska32_fa4_16_or0[0]), .fa_xor1(u_csamul_cska32_fa4_17_xor1), .fa_or0(u_csamul_cska32_fa4_17_or0));
  and_gate and_gate_u_csamul_cska32_and5_17(.a(a[5]), .b(b[17]), .out(u_csamul_cska32_and5_17));
  fa fa_u_csamul_cska32_fa5_17_out(.a(u_csamul_cska32_and5_17[0]), .b(u_csamul_cska32_fa6_16_xor1[0]), .cin(u_csamul_cska32_fa5_16_or0[0]), .fa_xor1(u_csamul_cska32_fa5_17_xor1), .fa_or0(u_csamul_cska32_fa5_17_or0));
  and_gate and_gate_u_csamul_cska32_and6_17(.a(a[6]), .b(b[17]), .out(u_csamul_cska32_and6_17));
  fa fa_u_csamul_cska32_fa6_17_out(.a(u_csamul_cska32_and6_17[0]), .b(u_csamul_cska32_fa7_16_xor1[0]), .cin(u_csamul_cska32_fa6_16_or0[0]), .fa_xor1(u_csamul_cska32_fa6_17_xor1), .fa_or0(u_csamul_cska32_fa6_17_or0));
  and_gate and_gate_u_csamul_cska32_and7_17(.a(a[7]), .b(b[17]), .out(u_csamul_cska32_and7_17));
  fa fa_u_csamul_cska32_fa7_17_out(.a(u_csamul_cska32_and7_17[0]), .b(u_csamul_cska32_fa8_16_xor1[0]), .cin(u_csamul_cska32_fa7_16_or0[0]), .fa_xor1(u_csamul_cska32_fa7_17_xor1), .fa_or0(u_csamul_cska32_fa7_17_or0));
  and_gate and_gate_u_csamul_cska32_and8_17(.a(a[8]), .b(b[17]), .out(u_csamul_cska32_and8_17));
  fa fa_u_csamul_cska32_fa8_17_out(.a(u_csamul_cska32_and8_17[0]), .b(u_csamul_cska32_fa9_16_xor1[0]), .cin(u_csamul_cska32_fa8_16_or0[0]), .fa_xor1(u_csamul_cska32_fa8_17_xor1), .fa_or0(u_csamul_cska32_fa8_17_or0));
  and_gate and_gate_u_csamul_cska32_and9_17(.a(a[9]), .b(b[17]), .out(u_csamul_cska32_and9_17));
  fa fa_u_csamul_cska32_fa9_17_out(.a(u_csamul_cska32_and9_17[0]), .b(u_csamul_cska32_fa10_16_xor1[0]), .cin(u_csamul_cska32_fa9_16_or0[0]), .fa_xor1(u_csamul_cska32_fa9_17_xor1), .fa_or0(u_csamul_cska32_fa9_17_or0));
  and_gate and_gate_u_csamul_cska32_and10_17(.a(a[10]), .b(b[17]), .out(u_csamul_cska32_and10_17));
  fa fa_u_csamul_cska32_fa10_17_out(.a(u_csamul_cska32_and10_17[0]), .b(u_csamul_cska32_fa11_16_xor1[0]), .cin(u_csamul_cska32_fa10_16_or0[0]), .fa_xor1(u_csamul_cska32_fa10_17_xor1), .fa_or0(u_csamul_cska32_fa10_17_or0));
  and_gate and_gate_u_csamul_cska32_and11_17(.a(a[11]), .b(b[17]), .out(u_csamul_cska32_and11_17));
  fa fa_u_csamul_cska32_fa11_17_out(.a(u_csamul_cska32_and11_17[0]), .b(u_csamul_cska32_fa12_16_xor1[0]), .cin(u_csamul_cska32_fa11_16_or0[0]), .fa_xor1(u_csamul_cska32_fa11_17_xor1), .fa_or0(u_csamul_cska32_fa11_17_or0));
  and_gate and_gate_u_csamul_cska32_and12_17(.a(a[12]), .b(b[17]), .out(u_csamul_cska32_and12_17));
  fa fa_u_csamul_cska32_fa12_17_out(.a(u_csamul_cska32_and12_17[0]), .b(u_csamul_cska32_fa13_16_xor1[0]), .cin(u_csamul_cska32_fa12_16_or0[0]), .fa_xor1(u_csamul_cska32_fa12_17_xor1), .fa_or0(u_csamul_cska32_fa12_17_or0));
  and_gate and_gate_u_csamul_cska32_and13_17(.a(a[13]), .b(b[17]), .out(u_csamul_cska32_and13_17));
  fa fa_u_csamul_cska32_fa13_17_out(.a(u_csamul_cska32_and13_17[0]), .b(u_csamul_cska32_fa14_16_xor1[0]), .cin(u_csamul_cska32_fa13_16_or0[0]), .fa_xor1(u_csamul_cska32_fa13_17_xor1), .fa_or0(u_csamul_cska32_fa13_17_or0));
  and_gate and_gate_u_csamul_cska32_and14_17(.a(a[14]), .b(b[17]), .out(u_csamul_cska32_and14_17));
  fa fa_u_csamul_cska32_fa14_17_out(.a(u_csamul_cska32_and14_17[0]), .b(u_csamul_cska32_fa15_16_xor1[0]), .cin(u_csamul_cska32_fa14_16_or0[0]), .fa_xor1(u_csamul_cska32_fa14_17_xor1), .fa_or0(u_csamul_cska32_fa14_17_or0));
  and_gate and_gate_u_csamul_cska32_and15_17(.a(a[15]), .b(b[17]), .out(u_csamul_cska32_and15_17));
  fa fa_u_csamul_cska32_fa15_17_out(.a(u_csamul_cska32_and15_17[0]), .b(u_csamul_cska32_fa16_16_xor1[0]), .cin(u_csamul_cska32_fa15_16_or0[0]), .fa_xor1(u_csamul_cska32_fa15_17_xor1), .fa_or0(u_csamul_cska32_fa15_17_or0));
  and_gate and_gate_u_csamul_cska32_and16_17(.a(a[16]), .b(b[17]), .out(u_csamul_cska32_and16_17));
  fa fa_u_csamul_cska32_fa16_17_out(.a(u_csamul_cska32_and16_17[0]), .b(u_csamul_cska32_fa17_16_xor1[0]), .cin(u_csamul_cska32_fa16_16_or0[0]), .fa_xor1(u_csamul_cska32_fa16_17_xor1), .fa_or0(u_csamul_cska32_fa16_17_or0));
  and_gate and_gate_u_csamul_cska32_and17_17(.a(a[17]), .b(b[17]), .out(u_csamul_cska32_and17_17));
  fa fa_u_csamul_cska32_fa17_17_out(.a(u_csamul_cska32_and17_17[0]), .b(u_csamul_cska32_fa18_16_xor1[0]), .cin(u_csamul_cska32_fa17_16_or0[0]), .fa_xor1(u_csamul_cska32_fa17_17_xor1), .fa_or0(u_csamul_cska32_fa17_17_or0));
  and_gate and_gate_u_csamul_cska32_and18_17(.a(a[18]), .b(b[17]), .out(u_csamul_cska32_and18_17));
  fa fa_u_csamul_cska32_fa18_17_out(.a(u_csamul_cska32_and18_17[0]), .b(u_csamul_cska32_fa19_16_xor1[0]), .cin(u_csamul_cska32_fa18_16_or0[0]), .fa_xor1(u_csamul_cska32_fa18_17_xor1), .fa_or0(u_csamul_cska32_fa18_17_or0));
  and_gate and_gate_u_csamul_cska32_and19_17(.a(a[19]), .b(b[17]), .out(u_csamul_cska32_and19_17));
  fa fa_u_csamul_cska32_fa19_17_out(.a(u_csamul_cska32_and19_17[0]), .b(u_csamul_cska32_fa20_16_xor1[0]), .cin(u_csamul_cska32_fa19_16_or0[0]), .fa_xor1(u_csamul_cska32_fa19_17_xor1), .fa_or0(u_csamul_cska32_fa19_17_or0));
  and_gate and_gate_u_csamul_cska32_and20_17(.a(a[20]), .b(b[17]), .out(u_csamul_cska32_and20_17));
  fa fa_u_csamul_cska32_fa20_17_out(.a(u_csamul_cska32_and20_17[0]), .b(u_csamul_cska32_fa21_16_xor1[0]), .cin(u_csamul_cska32_fa20_16_or0[0]), .fa_xor1(u_csamul_cska32_fa20_17_xor1), .fa_or0(u_csamul_cska32_fa20_17_or0));
  and_gate and_gate_u_csamul_cska32_and21_17(.a(a[21]), .b(b[17]), .out(u_csamul_cska32_and21_17));
  fa fa_u_csamul_cska32_fa21_17_out(.a(u_csamul_cska32_and21_17[0]), .b(u_csamul_cska32_fa22_16_xor1[0]), .cin(u_csamul_cska32_fa21_16_or0[0]), .fa_xor1(u_csamul_cska32_fa21_17_xor1), .fa_or0(u_csamul_cska32_fa21_17_or0));
  and_gate and_gate_u_csamul_cska32_and22_17(.a(a[22]), .b(b[17]), .out(u_csamul_cska32_and22_17));
  fa fa_u_csamul_cska32_fa22_17_out(.a(u_csamul_cska32_and22_17[0]), .b(u_csamul_cska32_fa23_16_xor1[0]), .cin(u_csamul_cska32_fa22_16_or0[0]), .fa_xor1(u_csamul_cska32_fa22_17_xor1), .fa_or0(u_csamul_cska32_fa22_17_or0));
  and_gate and_gate_u_csamul_cska32_and23_17(.a(a[23]), .b(b[17]), .out(u_csamul_cska32_and23_17));
  fa fa_u_csamul_cska32_fa23_17_out(.a(u_csamul_cska32_and23_17[0]), .b(u_csamul_cska32_fa24_16_xor1[0]), .cin(u_csamul_cska32_fa23_16_or0[0]), .fa_xor1(u_csamul_cska32_fa23_17_xor1), .fa_or0(u_csamul_cska32_fa23_17_or0));
  and_gate and_gate_u_csamul_cska32_and24_17(.a(a[24]), .b(b[17]), .out(u_csamul_cska32_and24_17));
  fa fa_u_csamul_cska32_fa24_17_out(.a(u_csamul_cska32_and24_17[0]), .b(u_csamul_cska32_fa25_16_xor1[0]), .cin(u_csamul_cska32_fa24_16_or0[0]), .fa_xor1(u_csamul_cska32_fa24_17_xor1), .fa_or0(u_csamul_cska32_fa24_17_or0));
  and_gate and_gate_u_csamul_cska32_and25_17(.a(a[25]), .b(b[17]), .out(u_csamul_cska32_and25_17));
  fa fa_u_csamul_cska32_fa25_17_out(.a(u_csamul_cska32_and25_17[0]), .b(u_csamul_cska32_fa26_16_xor1[0]), .cin(u_csamul_cska32_fa25_16_or0[0]), .fa_xor1(u_csamul_cska32_fa25_17_xor1), .fa_or0(u_csamul_cska32_fa25_17_or0));
  and_gate and_gate_u_csamul_cska32_and26_17(.a(a[26]), .b(b[17]), .out(u_csamul_cska32_and26_17));
  fa fa_u_csamul_cska32_fa26_17_out(.a(u_csamul_cska32_and26_17[0]), .b(u_csamul_cska32_fa27_16_xor1[0]), .cin(u_csamul_cska32_fa26_16_or0[0]), .fa_xor1(u_csamul_cska32_fa26_17_xor1), .fa_or0(u_csamul_cska32_fa26_17_or0));
  and_gate and_gate_u_csamul_cska32_and27_17(.a(a[27]), .b(b[17]), .out(u_csamul_cska32_and27_17));
  fa fa_u_csamul_cska32_fa27_17_out(.a(u_csamul_cska32_and27_17[0]), .b(u_csamul_cska32_fa28_16_xor1[0]), .cin(u_csamul_cska32_fa27_16_or0[0]), .fa_xor1(u_csamul_cska32_fa27_17_xor1), .fa_or0(u_csamul_cska32_fa27_17_or0));
  and_gate and_gate_u_csamul_cska32_and28_17(.a(a[28]), .b(b[17]), .out(u_csamul_cska32_and28_17));
  fa fa_u_csamul_cska32_fa28_17_out(.a(u_csamul_cska32_and28_17[0]), .b(u_csamul_cska32_fa29_16_xor1[0]), .cin(u_csamul_cska32_fa28_16_or0[0]), .fa_xor1(u_csamul_cska32_fa28_17_xor1), .fa_or0(u_csamul_cska32_fa28_17_or0));
  and_gate and_gate_u_csamul_cska32_and29_17(.a(a[29]), .b(b[17]), .out(u_csamul_cska32_and29_17));
  fa fa_u_csamul_cska32_fa29_17_out(.a(u_csamul_cska32_and29_17[0]), .b(u_csamul_cska32_fa30_16_xor1[0]), .cin(u_csamul_cska32_fa29_16_or0[0]), .fa_xor1(u_csamul_cska32_fa29_17_xor1), .fa_or0(u_csamul_cska32_fa29_17_or0));
  and_gate and_gate_u_csamul_cska32_and30_17(.a(a[30]), .b(b[17]), .out(u_csamul_cska32_and30_17));
  fa fa_u_csamul_cska32_fa30_17_out(.a(u_csamul_cska32_and30_17[0]), .b(u_csamul_cska32_and31_16[0]), .cin(u_csamul_cska32_fa30_16_or0[0]), .fa_xor1(u_csamul_cska32_fa30_17_xor1), .fa_or0(u_csamul_cska32_fa30_17_or0));
  and_gate and_gate_u_csamul_cska32_and31_17(.a(a[31]), .b(b[17]), .out(u_csamul_cska32_and31_17));
  and_gate and_gate_u_csamul_cska32_and0_18(.a(a[0]), .b(b[18]), .out(u_csamul_cska32_and0_18));
  fa fa_u_csamul_cska32_fa0_18_out(.a(u_csamul_cska32_and0_18[0]), .b(u_csamul_cska32_fa1_17_xor1[0]), .cin(u_csamul_cska32_fa0_17_or0[0]), .fa_xor1(u_csamul_cska32_fa0_18_xor1), .fa_or0(u_csamul_cska32_fa0_18_or0));
  and_gate and_gate_u_csamul_cska32_and1_18(.a(a[1]), .b(b[18]), .out(u_csamul_cska32_and1_18));
  fa fa_u_csamul_cska32_fa1_18_out(.a(u_csamul_cska32_and1_18[0]), .b(u_csamul_cska32_fa2_17_xor1[0]), .cin(u_csamul_cska32_fa1_17_or0[0]), .fa_xor1(u_csamul_cska32_fa1_18_xor1), .fa_or0(u_csamul_cska32_fa1_18_or0));
  and_gate and_gate_u_csamul_cska32_and2_18(.a(a[2]), .b(b[18]), .out(u_csamul_cska32_and2_18));
  fa fa_u_csamul_cska32_fa2_18_out(.a(u_csamul_cska32_and2_18[0]), .b(u_csamul_cska32_fa3_17_xor1[0]), .cin(u_csamul_cska32_fa2_17_or0[0]), .fa_xor1(u_csamul_cska32_fa2_18_xor1), .fa_or0(u_csamul_cska32_fa2_18_or0));
  and_gate and_gate_u_csamul_cska32_and3_18(.a(a[3]), .b(b[18]), .out(u_csamul_cska32_and3_18));
  fa fa_u_csamul_cska32_fa3_18_out(.a(u_csamul_cska32_and3_18[0]), .b(u_csamul_cska32_fa4_17_xor1[0]), .cin(u_csamul_cska32_fa3_17_or0[0]), .fa_xor1(u_csamul_cska32_fa3_18_xor1), .fa_or0(u_csamul_cska32_fa3_18_or0));
  and_gate and_gate_u_csamul_cska32_and4_18(.a(a[4]), .b(b[18]), .out(u_csamul_cska32_and4_18));
  fa fa_u_csamul_cska32_fa4_18_out(.a(u_csamul_cska32_and4_18[0]), .b(u_csamul_cska32_fa5_17_xor1[0]), .cin(u_csamul_cska32_fa4_17_or0[0]), .fa_xor1(u_csamul_cska32_fa4_18_xor1), .fa_or0(u_csamul_cska32_fa4_18_or0));
  and_gate and_gate_u_csamul_cska32_and5_18(.a(a[5]), .b(b[18]), .out(u_csamul_cska32_and5_18));
  fa fa_u_csamul_cska32_fa5_18_out(.a(u_csamul_cska32_and5_18[0]), .b(u_csamul_cska32_fa6_17_xor1[0]), .cin(u_csamul_cska32_fa5_17_or0[0]), .fa_xor1(u_csamul_cska32_fa5_18_xor1), .fa_or0(u_csamul_cska32_fa5_18_or0));
  and_gate and_gate_u_csamul_cska32_and6_18(.a(a[6]), .b(b[18]), .out(u_csamul_cska32_and6_18));
  fa fa_u_csamul_cska32_fa6_18_out(.a(u_csamul_cska32_and6_18[0]), .b(u_csamul_cska32_fa7_17_xor1[0]), .cin(u_csamul_cska32_fa6_17_or0[0]), .fa_xor1(u_csamul_cska32_fa6_18_xor1), .fa_or0(u_csamul_cska32_fa6_18_or0));
  and_gate and_gate_u_csamul_cska32_and7_18(.a(a[7]), .b(b[18]), .out(u_csamul_cska32_and7_18));
  fa fa_u_csamul_cska32_fa7_18_out(.a(u_csamul_cska32_and7_18[0]), .b(u_csamul_cska32_fa8_17_xor1[0]), .cin(u_csamul_cska32_fa7_17_or0[0]), .fa_xor1(u_csamul_cska32_fa7_18_xor1), .fa_or0(u_csamul_cska32_fa7_18_or0));
  and_gate and_gate_u_csamul_cska32_and8_18(.a(a[8]), .b(b[18]), .out(u_csamul_cska32_and8_18));
  fa fa_u_csamul_cska32_fa8_18_out(.a(u_csamul_cska32_and8_18[0]), .b(u_csamul_cska32_fa9_17_xor1[0]), .cin(u_csamul_cska32_fa8_17_or0[0]), .fa_xor1(u_csamul_cska32_fa8_18_xor1), .fa_or0(u_csamul_cska32_fa8_18_or0));
  and_gate and_gate_u_csamul_cska32_and9_18(.a(a[9]), .b(b[18]), .out(u_csamul_cska32_and9_18));
  fa fa_u_csamul_cska32_fa9_18_out(.a(u_csamul_cska32_and9_18[0]), .b(u_csamul_cska32_fa10_17_xor1[0]), .cin(u_csamul_cska32_fa9_17_or0[0]), .fa_xor1(u_csamul_cska32_fa9_18_xor1), .fa_or0(u_csamul_cska32_fa9_18_or0));
  and_gate and_gate_u_csamul_cska32_and10_18(.a(a[10]), .b(b[18]), .out(u_csamul_cska32_and10_18));
  fa fa_u_csamul_cska32_fa10_18_out(.a(u_csamul_cska32_and10_18[0]), .b(u_csamul_cska32_fa11_17_xor1[0]), .cin(u_csamul_cska32_fa10_17_or0[0]), .fa_xor1(u_csamul_cska32_fa10_18_xor1), .fa_or0(u_csamul_cska32_fa10_18_or0));
  and_gate and_gate_u_csamul_cska32_and11_18(.a(a[11]), .b(b[18]), .out(u_csamul_cska32_and11_18));
  fa fa_u_csamul_cska32_fa11_18_out(.a(u_csamul_cska32_and11_18[0]), .b(u_csamul_cska32_fa12_17_xor1[0]), .cin(u_csamul_cska32_fa11_17_or0[0]), .fa_xor1(u_csamul_cska32_fa11_18_xor1), .fa_or0(u_csamul_cska32_fa11_18_or0));
  and_gate and_gate_u_csamul_cska32_and12_18(.a(a[12]), .b(b[18]), .out(u_csamul_cska32_and12_18));
  fa fa_u_csamul_cska32_fa12_18_out(.a(u_csamul_cska32_and12_18[0]), .b(u_csamul_cska32_fa13_17_xor1[0]), .cin(u_csamul_cska32_fa12_17_or0[0]), .fa_xor1(u_csamul_cska32_fa12_18_xor1), .fa_or0(u_csamul_cska32_fa12_18_or0));
  and_gate and_gate_u_csamul_cska32_and13_18(.a(a[13]), .b(b[18]), .out(u_csamul_cska32_and13_18));
  fa fa_u_csamul_cska32_fa13_18_out(.a(u_csamul_cska32_and13_18[0]), .b(u_csamul_cska32_fa14_17_xor1[0]), .cin(u_csamul_cska32_fa13_17_or0[0]), .fa_xor1(u_csamul_cska32_fa13_18_xor1), .fa_or0(u_csamul_cska32_fa13_18_or0));
  and_gate and_gate_u_csamul_cska32_and14_18(.a(a[14]), .b(b[18]), .out(u_csamul_cska32_and14_18));
  fa fa_u_csamul_cska32_fa14_18_out(.a(u_csamul_cska32_and14_18[0]), .b(u_csamul_cska32_fa15_17_xor1[0]), .cin(u_csamul_cska32_fa14_17_or0[0]), .fa_xor1(u_csamul_cska32_fa14_18_xor1), .fa_or0(u_csamul_cska32_fa14_18_or0));
  and_gate and_gate_u_csamul_cska32_and15_18(.a(a[15]), .b(b[18]), .out(u_csamul_cska32_and15_18));
  fa fa_u_csamul_cska32_fa15_18_out(.a(u_csamul_cska32_and15_18[0]), .b(u_csamul_cska32_fa16_17_xor1[0]), .cin(u_csamul_cska32_fa15_17_or0[0]), .fa_xor1(u_csamul_cska32_fa15_18_xor1), .fa_or0(u_csamul_cska32_fa15_18_or0));
  and_gate and_gate_u_csamul_cska32_and16_18(.a(a[16]), .b(b[18]), .out(u_csamul_cska32_and16_18));
  fa fa_u_csamul_cska32_fa16_18_out(.a(u_csamul_cska32_and16_18[0]), .b(u_csamul_cska32_fa17_17_xor1[0]), .cin(u_csamul_cska32_fa16_17_or0[0]), .fa_xor1(u_csamul_cska32_fa16_18_xor1), .fa_or0(u_csamul_cska32_fa16_18_or0));
  and_gate and_gate_u_csamul_cska32_and17_18(.a(a[17]), .b(b[18]), .out(u_csamul_cska32_and17_18));
  fa fa_u_csamul_cska32_fa17_18_out(.a(u_csamul_cska32_and17_18[0]), .b(u_csamul_cska32_fa18_17_xor1[0]), .cin(u_csamul_cska32_fa17_17_or0[0]), .fa_xor1(u_csamul_cska32_fa17_18_xor1), .fa_or0(u_csamul_cska32_fa17_18_or0));
  and_gate and_gate_u_csamul_cska32_and18_18(.a(a[18]), .b(b[18]), .out(u_csamul_cska32_and18_18));
  fa fa_u_csamul_cska32_fa18_18_out(.a(u_csamul_cska32_and18_18[0]), .b(u_csamul_cska32_fa19_17_xor1[0]), .cin(u_csamul_cska32_fa18_17_or0[0]), .fa_xor1(u_csamul_cska32_fa18_18_xor1), .fa_or0(u_csamul_cska32_fa18_18_or0));
  and_gate and_gate_u_csamul_cska32_and19_18(.a(a[19]), .b(b[18]), .out(u_csamul_cska32_and19_18));
  fa fa_u_csamul_cska32_fa19_18_out(.a(u_csamul_cska32_and19_18[0]), .b(u_csamul_cska32_fa20_17_xor1[0]), .cin(u_csamul_cska32_fa19_17_or0[0]), .fa_xor1(u_csamul_cska32_fa19_18_xor1), .fa_or0(u_csamul_cska32_fa19_18_or0));
  and_gate and_gate_u_csamul_cska32_and20_18(.a(a[20]), .b(b[18]), .out(u_csamul_cska32_and20_18));
  fa fa_u_csamul_cska32_fa20_18_out(.a(u_csamul_cska32_and20_18[0]), .b(u_csamul_cska32_fa21_17_xor1[0]), .cin(u_csamul_cska32_fa20_17_or0[0]), .fa_xor1(u_csamul_cska32_fa20_18_xor1), .fa_or0(u_csamul_cska32_fa20_18_or0));
  and_gate and_gate_u_csamul_cska32_and21_18(.a(a[21]), .b(b[18]), .out(u_csamul_cska32_and21_18));
  fa fa_u_csamul_cska32_fa21_18_out(.a(u_csamul_cska32_and21_18[0]), .b(u_csamul_cska32_fa22_17_xor1[0]), .cin(u_csamul_cska32_fa21_17_or0[0]), .fa_xor1(u_csamul_cska32_fa21_18_xor1), .fa_or0(u_csamul_cska32_fa21_18_or0));
  and_gate and_gate_u_csamul_cska32_and22_18(.a(a[22]), .b(b[18]), .out(u_csamul_cska32_and22_18));
  fa fa_u_csamul_cska32_fa22_18_out(.a(u_csamul_cska32_and22_18[0]), .b(u_csamul_cska32_fa23_17_xor1[0]), .cin(u_csamul_cska32_fa22_17_or0[0]), .fa_xor1(u_csamul_cska32_fa22_18_xor1), .fa_or0(u_csamul_cska32_fa22_18_or0));
  and_gate and_gate_u_csamul_cska32_and23_18(.a(a[23]), .b(b[18]), .out(u_csamul_cska32_and23_18));
  fa fa_u_csamul_cska32_fa23_18_out(.a(u_csamul_cska32_and23_18[0]), .b(u_csamul_cska32_fa24_17_xor1[0]), .cin(u_csamul_cska32_fa23_17_or0[0]), .fa_xor1(u_csamul_cska32_fa23_18_xor1), .fa_or0(u_csamul_cska32_fa23_18_or0));
  and_gate and_gate_u_csamul_cska32_and24_18(.a(a[24]), .b(b[18]), .out(u_csamul_cska32_and24_18));
  fa fa_u_csamul_cska32_fa24_18_out(.a(u_csamul_cska32_and24_18[0]), .b(u_csamul_cska32_fa25_17_xor1[0]), .cin(u_csamul_cska32_fa24_17_or0[0]), .fa_xor1(u_csamul_cska32_fa24_18_xor1), .fa_or0(u_csamul_cska32_fa24_18_or0));
  and_gate and_gate_u_csamul_cska32_and25_18(.a(a[25]), .b(b[18]), .out(u_csamul_cska32_and25_18));
  fa fa_u_csamul_cska32_fa25_18_out(.a(u_csamul_cska32_and25_18[0]), .b(u_csamul_cska32_fa26_17_xor1[0]), .cin(u_csamul_cska32_fa25_17_or0[0]), .fa_xor1(u_csamul_cska32_fa25_18_xor1), .fa_or0(u_csamul_cska32_fa25_18_or0));
  and_gate and_gate_u_csamul_cska32_and26_18(.a(a[26]), .b(b[18]), .out(u_csamul_cska32_and26_18));
  fa fa_u_csamul_cska32_fa26_18_out(.a(u_csamul_cska32_and26_18[0]), .b(u_csamul_cska32_fa27_17_xor1[0]), .cin(u_csamul_cska32_fa26_17_or0[0]), .fa_xor1(u_csamul_cska32_fa26_18_xor1), .fa_or0(u_csamul_cska32_fa26_18_or0));
  and_gate and_gate_u_csamul_cska32_and27_18(.a(a[27]), .b(b[18]), .out(u_csamul_cska32_and27_18));
  fa fa_u_csamul_cska32_fa27_18_out(.a(u_csamul_cska32_and27_18[0]), .b(u_csamul_cska32_fa28_17_xor1[0]), .cin(u_csamul_cska32_fa27_17_or0[0]), .fa_xor1(u_csamul_cska32_fa27_18_xor1), .fa_or0(u_csamul_cska32_fa27_18_or0));
  and_gate and_gate_u_csamul_cska32_and28_18(.a(a[28]), .b(b[18]), .out(u_csamul_cska32_and28_18));
  fa fa_u_csamul_cska32_fa28_18_out(.a(u_csamul_cska32_and28_18[0]), .b(u_csamul_cska32_fa29_17_xor1[0]), .cin(u_csamul_cska32_fa28_17_or0[0]), .fa_xor1(u_csamul_cska32_fa28_18_xor1), .fa_or0(u_csamul_cska32_fa28_18_or0));
  and_gate and_gate_u_csamul_cska32_and29_18(.a(a[29]), .b(b[18]), .out(u_csamul_cska32_and29_18));
  fa fa_u_csamul_cska32_fa29_18_out(.a(u_csamul_cska32_and29_18[0]), .b(u_csamul_cska32_fa30_17_xor1[0]), .cin(u_csamul_cska32_fa29_17_or0[0]), .fa_xor1(u_csamul_cska32_fa29_18_xor1), .fa_or0(u_csamul_cska32_fa29_18_or0));
  and_gate and_gate_u_csamul_cska32_and30_18(.a(a[30]), .b(b[18]), .out(u_csamul_cska32_and30_18));
  fa fa_u_csamul_cska32_fa30_18_out(.a(u_csamul_cska32_and30_18[0]), .b(u_csamul_cska32_and31_17[0]), .cin(u_csamul_cska32_fa30_17_or0[0]), .fa_xor1(u_csamul_cska32_fa30_18_xor1), .fa_or0(u_csamul_cska32_fa30_18_or0));
  and_gate and_gate_u_csamul_cska32_and31_18(.a(a[31]), .b(b[18]), .out(u_csamul_cska32_and31_18));
  and_gate and_gate_u_csamul_cska32_and0_19(.a(a[0]), .b(b[19]), .out(u_csamul_cska32_and0_19));
  fa fa_u_csamul_cska32_fa0_19_out(.a(u_csamul_cska32_and0_19[0]), .b(u_csamul_cska32_fa1_18_xor1[0]), .cin(u_csamul_cska32_fa0_18_or0[0]), .fa_xor1(u_csamul_cska32_fa0_19_xor1), .fa_or0(u_csamul_cska32_fa0_19_or0));
  and_gate and_gate_u_csamul_cska32_and1_19(.a(a[1]), .b(b[19]), .out(u_csamul_cska32_and1_19));
  fa fa_u_csamul_cska32_fa1_19_out(.a(u_csamul_cska32_and1_19[0]), .b(u_csamul_cska32_fa2_18_xor1[0]), .cin(u_csamul_cska32_fa1_18_or0[0]), .fa_xor1(u_csamul_cska32_fa1_19_xor1), .fa_or0(u_csamul_cska32_fa1_19_or0));
  and_gate and_gate_u_csamul_cska32_and2_19(.a(a[2]), .b(b[19]), .out(u_csamul_cska32_and2_19));
  fa fa_u_csamul_cska32_fa2_19_out(.a(u_csamul_cska32_and2_19[0]), .b(u_csamul_cska32_fa3_18_xor1[0]), .cin(u_csamul_cska32_fa2_18_or0[0]), .fa_xor1(u_csamul_cska32_fa2_19_xor1), .fa_or0(u_csamul_cska32_fa2_19_or0));
  and_gate and_gate_u_csamul_cska32_and3_19(.a(a[3]), .b(b[19]), .out(u_csamul_cska32_and3_19));
  fa fa_u_csamul_cska32_fa3_19_out(.a(u_csamul_cska32_and3_19[0]), .b(u_csamul_cska32_fa4_18_xor1[0]), .cin(u_csamul_cska32_fa3_18_or0[0]), .fa_xor1(u_csamul_cska32_fa3_19_xor1), .fa_or0(u_csamul_cska32_fa3_19_or0));
  and_gate and_gate_u_csamul_cska32_and4_19(.a(a[4]), .b(b[19]), .out(u_csamul_cska32_and4_19));
  fa fa_u_csamul_cska32_fa4_19_out(.a(u_csamul_cska32_and4_19[0]), .b(u_csamul_cska32_fa5_18_xor1[0]), .cin(u_csamul_cska32_fa4_18_or0[0]), .fa_xor1(u_csamul_cska32_fa4_19_xor1), .fa_or0(u_csamul_cska32_fa4_19_or0));
  and_gate and_gate_u_csamul_cska32_and5_19(.a(a[5]), .b(b[19]), .out(u_csamul_cska32_and5_19));
  fa fa_u_csamul_cska32_fa5_19_out(.a(u_csamul_cska32_and5_19[0]), .b(u_csamul_cska32_fa6_18_xor1[0]), .cin(u_csamul_cska32_fa5_18_or0[0]), .fa_xor1(u_csamul_cska32_fa5_19_xor1), .fa_or0(u_csamul_cska32_fa5_19_or0));
  and_gate and_gate_u_csamul_cska32_and6_19(.a(a[6]), .b(b[19]), .out(u_csamul_cska32_and6_19));
  fa fa_u_csamul_cska32_fa6_19_out(.a(u_csamul_cska32_and6_19[0]), .b(u_csamul_cska32_fa7_18_xor1[0]), .cin(u_csamul_cska32_fa6_18_or0[0]), .fa_xor1(u_csamul_cska32_fa6_19_xor1), .fa_or0(u_csamul_cska32_fa6_19_or0));
  and_gate and_gate_u_csamul_cska32_and7_19(.a(a[7]), .b(b[19]), .out(u_csamul_cska32_and7_19));
  fa fa_u_csamul_cska32_fa7_19_out(.a(u_csamul_cska32_and7_19[0]), .b(u_csamul_cska32_fa8_18_xor1[0]), .cin(u_csamul_cska32_fa7_18_or0[0]), .fa_xor1(u_csamul_cska32_fa7_19_xor1), .fa_or0(u_csamul_cska32_fa7_19_or0));
  and_gate and_gate_u_csamul_cska32_and8_19(.a(a[8]), .b(b[19]), .out(u_csamul_cska32_and8_19));
  fa fa_u_csamul_cska32_fa8_19_out(.a(u_csamul_cska32_and8_19[0]), .b(u_csamul_cska32_fa9_18_xor1[0]), .cin(u_csamul_cska32_fa8_18_or0[0]), .fa_xor1(u_csamul_cska32_fa8_19_xor1), .fa_or0(u_csamul_cska32_fa8_19_or0));
  and_gate and_gate_u_csamul_cska32_and9_19(.a(a[9]), .b(b[19]), .out(u_csamul_cska32_and9_19));
  fa fa_u_csamul_cska32_fa9_19_out(.a(u_csamul_cska32_and9_19[0]), .b(u_csamul_cska32_fa10_18_xor1[0]), .cin(u_csamul_cska32_fa9_18_or0[0]), .fa_xor1(u_csamul_cska32_fa9_19_xor1), .fa_or0(u_csamul_cska32_fa9_19_or0));
  and_gate and_gate_u_csamul_cska32_and10_19(.a(a[10]), .b(b[19]), .out(u_csamul_cska32_and10_19));
  fa fa_u_csamul_cska32_fa10_19_out(.a(u_csamul_cska32_and10_19[0]), .b(u_csamul_cska32_fa11_18_xor1[0]), .cin(u_csamul_cska32_fa10_18_or0[0]), .fa_xor1(u_csamul_cska32_fa10_19_xor1), .fa_or0(u_csamul_cska32_fa10_19_or0));
  and_gate and_gate_u_csamul_cska32_and11_19(.a(a[11]), .b(b[19]), .out(u_csamul_cska32_and11_19));
  fa fa_u_csamul_cska32_fa11_19_out(.a(u_csamul_cska32_and11_19[0]), .b(u_csamul_cska32_fa12_18_xor1[0]), .cin(u_csamul_cska32_fa11_18_or0[0]), .fa_xor1(u_csamul_cska32_fa11_19_xor1), .fa_or0(u_csamul_cska32_fa11_19_or0));
  and_gate and_gate_u_csamul_cska32_and12_19(.a(a[12]), .b(b[19]), .out(u_csamul_cska32_and12_19));
  fa fa_u_csamul_cska32_fa12_19_out(.a(u_csamul_cska32_and12_19[0]), .b(u_csamul_cska32_fa13_18_xor1[0]), .cin(u_csamul_cska32_fa12_18_or0[0]), .fa_xor1(u_csamul_cska32_fa12_19_xor1), .fa_or0(u_csamul_cska32_fa12_19_or0));
  and_gate and_gate_u_csamul_cska32_and13_19(.a(a[13]), .b(b[19]), .out(u_csamul_cska32_and13_19));
  fa fa_u_csamul_cska32_fa13_19_out(.a(u_csamul_cska32_and13_19[0]), .b(u_csamul_cska32_fa14_18_xor1[0]), .cin(u_csamul_cska32_fa13_18_or0[0]), .fa_xor1(u_csamul_cska32_fa13_19_xor1), .fa_or0(u_csamul_cska32_fa13_19_or0));
  and_gate and_gate_u_csamul_cska32_and14_19(.a(a[14]), .b(b[19]), .out(u_csamul_cska32_and14_19));
  fa fa_u_csamul_cska32_fa14_19_out(.a(u_csamul_cska32_and14_19[0]), .b(u_csamul_cska32_fa15_18_xor1[0]), .cin(u_csamul_cska32_fa14_18_or0[0]), .fa_xor1(u_csamul_cska32_fa14_19_xor1), .fa_or0(u_csamul_cska32_fa14_19_or0));
  and_gate and_gate_u_csamul_cska32_and15_19(.a(a[15]), .b(b[19]), .out(u_csamul_cska32_and15_19));
  fa fa_u_csamul_cska32_fa15_19_out(.a(u_csamul_cska32_and15_19[0]), .b(u_csamul_cska32_fa16_18_xor1[0]), .cin(u_csamul_cska32_fa15_18_or0[0]), .fa_xor1(u_csamul_cska32_fa15_19_xor1), .fa_or0(u_csamul_cska32_fa15_19_or0));
  and_gate and_gate_u_csamul_cska32_and16_19(.a(a[16]), .b(b[19]), .out(u_csamul_cska32_and16_19));
  fa fa_u_csamul_cska32_fa16_19_out(.a(u_csamul_cska32_and16_19[0]), .b(u_csamul_cska32_fa17_18_xor1[0]), .cin(u_csamul_cska32_fa16_18_or0[0]), .fa_xor1(u_csamul_cska32_fa16_19_xor1), .fa_or0(u_csamul_cska32_fa16_19_or0));
  and_gate and_gate_u_csamul_cska32_and17_19(.a(a[17]), .b(b[19]), .out(u_csamul_cska32_and17_19));
  fa fa_u_csamul_cska32_fa17_19_out(.a(u_csamul_cska32_and17_19[0]), .b(u_csamul_cska32_fa18_18_xor1[0]), .cin(u_csamul_cska32_fa17_18_or0[0]), .fa_xor1(u_csamul_cska32_fa17_19_xor1), .fa_or0(u_csamul_cska32_fa17_19_or0));
  and_gate and_gate_u_csamul_cska32_and18_19(.a(a[18]), .b(b[19]), .out(u_csamul_cska32_and18_19));
  fa fa_u_csamul_cska32_fa18_19_out(.a(u_csamul_cska32_and18_19[0]), .b(u_csamul_cska32_fa19_18_xor1[0]), .cin(u_csamul_cska32_fa18_18_or0[0]), .fa_xor1(u_csamul_cska32_fa18_19_xor1), .fa_or0(u_csamul_cska32_fa18_19_or0));
  and_gate and_gate_u_csamul_cska32_and19_19(.a(a[19]), .b(b[19]), .out(u_csamul_cska32_and19_19));
  fa fa_u_csamul_cska32_fa19_19_out(.a(u_csamul_cska32_and19_19[0]), .b(u_csamul_cska32_fa20_18_xor1[0]), .cin(u_csamul_cska32_fa19_18_or0[0]), .fa_xor1(u_csamul_cska32_fa19_19_xor1), .fa_or0(u_csamul_cska32_fa19_19_or0));
  and_gate and_gate_u_csamul_cska32_and20_19(.a(a[20]), .b(b[19]), .out(u_csamul_cska32_and20_19));
  fa fa_u_csamul_cska32_fa20_19_out(.a(u_csamul_cska32_and20_19[0]), .b(u_csamul_cska32_fa21_18_xor1[0]), .cin(u_csamul_cska32_fa20_18_or0[0]), .fa_xor1(u_csamul_cska32_fa20_19_xor1), .fa_or0(u_csamul_cska32_fa20_19_or0));
  and_gate and_gate_u_csamul_cska32_and21_19(.a(a[21]), .b(b[19]), .out(u_csamul_cska32_and21_19));
  fa fa_u_csamul_cska32_fa21_19_out(.a(u_csamul_cska32_and21_19[0]), .b(u_csamul_cska32_fa22_18_xor1[0]), .cin(u_csamul_cska32_fa21_18_or0[0]), .fa_xor1(u_csamul_cska32_fa21_19_xor1), .fa_or0(u_csamul_cska32_fa21_19_or0));
  and_gate and_gate_u_csamul_cska32_and22_19(.a(a[22]), .b(b[19]), .out(u_csamul_cska32_and22_19));
  fa fa_u_csamul_cska32_fa22_19_out(.a(u_csamul_cska32_and22_19[0]), .b(u_csamul_cska32_fa23_18_xor1[0]), .cin(u_csamul_cska32_fa22_18_or0[0]), .fa_xor1(u_csamul_cska32_fa22_19_xor1), .fa_or0(u_csamul_cska32_fa22_19_or0));
  and_gate and_gate_u_csamul_cska32_and23_19(.a(a[23]), .b(b[19]), .out(u_csamul_cska32_and23_19));
  fa fa_u_csamul_cska32_fa23_19_out(.a(u_csamul_cska32_and23_19[0]), .b(u_csamul_cska32_fa24_18_xor1[0]), .cin(u_csamul_cska32_fa23_18_or0[0]), .fa_xor1(u_csamul_cska32_fa23_19_xor1), .fa_or0(u_csamul_cska32_fa23_19_or0));
  and_gate and_gate_u_csamul_cska32_and24_19(.a(a[24]), .b(b[19]), .out(u_csamul_cska32_and24_19));
  fa fa_u_csamul_cska32_fa24_19_out(.a(u_csamul_cska32_and24_19[0]), .b(u_csamul_cska32_fa25_18_xor1[0]), .cin(u_csamul_cska32_fa24_18_or0[0]), .fa_xor1(u_csamul_cska32_fa24_19_xor1), .fa_or0(u_csamul_cska32_fa24_19_or0));
  and_gate and_gate_u_csamul_cska32_and25_19(.a(a[25]), .b(b[19]), .out(u_csamul_cska32_and25_19));
  fa fa_u_csamul_cska32_fa25_19_out(.a(u_csamul_cska32_and25_19[0]), .b(u_csamul_cska32_fa26_18_xor1[0]), .cin(u_csamul_cska32_fa25_18_or0[0]), .fa_xor1(u_csamul_cska32_fa25_19_xor1), .fa_or0(u_csamul_cska32_fa25_19_or0));
  and_gate and_gate_u_csamul_cska32_and26_19(.a(a[26]), .b(b[19]), .out(u_csamul_cska32_and26_19));
  fa fa_u_csamul_cska32_fa26_19_out(.a(u_csamul_cska32_and26_19[0]), .b(u_csamul_cska32_fa27_18_xor1[0]), .cin(u_csamul_cska32_fa26_18_or0[0]), .fa_xor1(u_csamul_cska32_fa26_19_xor1), .fa_or0(u_csamul_cska32_fa26_19_or0));
  and_gate and_gate_u_csamul_cska32_and27_19(.a(a[27]), .b(b[19]), .out(u_csamul_cska32_and27_19));
  fa fa_u_csamul_cska32_fa27_19_out(.a(u_csamul_cska32_and27_19[0]), .b(u_csamul_cska32_fa28_18_xor1[0]), .cin(u_csamul_cska32_fa27_18_or0[0]), .fa_xor1(u_csamul_cska32_fa27_19_xor1), .fa_or0(u_csamul_cska32_fa27_19_or0));
  and_gate and_gate_u_csamul_cska32_and28_19(.a(a[28]), .b(b[19]), .out(u_csamul_cska32_and28_19));
  fa fa_u_csamul_cska32_fa28_19_out(.a(u_csamul_cska32_and28_19[0]), .b(u_csamul_cska32_fa29_18_xor1[0]), .cin(u_csamul_cska32_fa28_18_or0[0]), .fa_xor1(u_csamul_cska32_fa28_19_xor1), .fa_or0(u_csamul_cska32_fa28_19_or0));
  and_gate and_gate_u_csamul_cska32_and29_19(.a(a[29]), .b(b[19]), .out(u_csamul_cska32_and29_19));
  fa fa_u_csamul_cska32_fa29_19_out(.a(u_csamul_cska32_and29_19[0]), .b(u_csamul_cska32_fa30_18_xor1[0]), .cin(u_csamul_cska32_fa29_18_or0[0]), .fa_xor1(u_csamul_cska32_fa29_19_xor1), .fa_or0(u_csamul_cska32_fa29_19_or0));
  and_gate and_gate_u_csamul_cska32_and30_19(.a(a[30]), .b(b[19]), .out(u_csamul_cska32_and30_19));
  fa fa_u_csamul_cska32_fa30_19_out(.a(u_csamul_cska32_and30_19[0]), .b(u_csamul_cska32_and31_18[0]), .cin(u_csamul_cska32_fa30_18_or0[0]), .fa_xor1(u_csamul_cska32_fa30_19_xor1), .fa_or0(u_csamul_cska32_fa30_19_or0));
  and_gate and_gate_u_csamul_cska32_and31_19(.a(a[31]), .b(b[19]), .out(u_csamul_cska32_and31_19));
  and_gate and_gate_u_csamul_cska32_and0_20(.a(a[0]), .b(b[20]), .out(u_csamul_cska32_and0_20));
  fa fa_u_csamul_cska32_fa0_20_out(.a(u_csamul_cska32_and0_20[0]), .b(u_csamul_cska32_fa1_19_xor1[0]), .cin(u_csamul_cska32_fa0_19_or0[0]), .fa_xor1(u_csamul_cska32_fa0_20_xor1), .fa_or0(u_csamul_cska32_fa0_20_or0));
  and_gate and_gate_u_csamul_cska32_and1_20(.a(a[1]), .b(b[20]), .out(u_csamul_cska32_and1_20));
  fa fa_u_csamul_cska32_fa1_20_out(.a(u_csamul_cska32_and1_20[0]), .b(u_csamul_cska32_fa2_19_xor1[0]), .cin(u_csamul_cska32_fa1_19_or0[0]), .fa_xor1(u_csamul_cska32_fa1_20_xor1), .fa_or0(u_csamul_cska32_fa1_20_or0));
  and_gate and_gate_u_csamul_cska32_and2_20(.a(a[2]), .b(b[20]), .out(u_csamul_cska32_and2_20));
  fa fa_u_csamul_cska32_fa2_20_out(.a(u_csamul_cska32_and2_20[0]), .b(u_csamul_cska32_fa3_19_xor1[0]), .cin(u_csamul_cska32_fa2_19_or0[0]), .fa_xor1(u_csamul_cska32_fa2_20_xor1), .fa_or0(u_csamul_cska32_fa2_20_or0));
  and_gate and_gate_u_csamul_cska32_and3_20(.a(a[3]), .b(b[20]), .out(u_csamul_cska32_and3_20));
  fa fa_u_csamul_cska32_fa3_20_out(.a(u_csamul_cska32_and3_20[0]), .b(u_csamul_cska32_fa4_19_xor1[0]), .cin(u_csamul_cska32_fa3_19_or0[0]), .fa_xor1(u_csamul_cska32_fa3_20_xor1), .fa_or0(u_csamul_cska32_fa3_20_or0));
  and_gate and_gate_u_csamul_cska32_and4_20(.a(a[4]), .b(b[20]), .out(u_csamul_cska32_and4_20));
  fa fa_u_csamul_cska32_fa4_20_out(.a(u_csamul_cska32_and4_20[0]), .b(u_csamul_cska32_fa5_19_xor1[0]), .cin(u_csamul_cska32_fa4_19_or0[0]), .fa_xor1(u_csamul_cska32_fa4_20_xor1), .fa_or0(u_csamul_cska32_fa4_20_or0));
  and_gate and_gate_u_csamul_cska32_and5_20(.a(a[5]), .b(b[20]), .out(u_csamul_cska32_and5_20));
  fa fa_u_csamul_cska32_fa5_20_out(.a(u_csamul_cska32_and5_20[0]), .b(u_csamul_cska32_fa6_19_xor1[0]), .cin(u_csamul_cska32_fa5_19_or0[0]), .fa_xor1(u_csamul_cska32_fa5_20_xor1), .fa_or0(u_csamul_cska32_fa5_20_or0));
  and_gate and_gate_u_csamul_cska32_and6_20(.a(a[6]), .b(b[20]), .out(u_csamul_cska32_and6_20));
  fa fa_u_csamul_cska32_fa6_20_out(.a(u_csamul_cska32_and6_20[0]), .b(u_csamul_cska32_fa7_19_xor1[0]), .cin(u_csamul_cska32_fa6_19_or0[0]), .fa_xor1(u_csamul_cska32_fa6_20_xor1), .fa_or0(u_csamul_cska32_fa6_20_or0));
  and_gate and_gate_u_csamul_cska32_and7_20(.a(a[7]), .b(b[20]), .out(u_csamul_cska32_and7_20));
  fa fa_u_csamul_cska32_fa7_20_out(.a(u_csamul_cska32_and7_20[0]), .b(u_csamul_cska32_fa8_19_xor1[0]), .cin(u_csamul_cska32_fa7_19_or0[0]), .fa_xor1(u_csamul_cska32_fa7_20_xor1), .fa_or0(u_csamul_cska32_fa7_20_or0));
  and_gate and_gate_u_csamul_cska32_and8_20(.a(a[8]), .b(b[20]), .out(u_csamul_cska32_and8_20));
  fa fa_u_csamul_cska32_fa8_20_out(.a(u_csamul_cska32_and8_20[0]), .b(u_csamul_cska32_fa9_19_xor1[0]), .cin(u_csamul_cska32_fa8_19_or0[0]), .fa_xor1(u_csamul_cska32_fa8_20_xor1), .fa_or0(u_csamul_cska32_fa8_20_or0));
  and_gate and_gate_u_csamul_cska32_and9_20(.a(a[9]), .b(b[20]), .out(u_csamul_cska32_and9_20));
  fa fa_u_csamul_cska32_fa9_20_out(.a(u_csamul_cska32_and9_20[0]), .b(u_csamul_cska32_fa10_19_xor1[0]), .cin(u_csamul_cska32_fa9_19_or0[0]), .fa_xor1(u_csamul_cska32_fa9_20_xor1), .fa_or0(u_csamul_cska32_fa9_20_or0));
  and_gate and_gate_u_csamul_cska32_and10_20(.a(a[10]), .b(b[20]), .out(u_csamul_cska32_and10_20));
  fa fa_u_csamul_cska32_fa10_20_out(.a(u_csamul_cska32_and10_20[0]), .b(u_csamul_cska32_fa11_19_xor1[0]), .cin(u_csamul_cska32_fa10_19_or0[0]), .fa_xor1(u_csamul_cska32_fa10_20_xor1), .fa_or0(u_csamul_cska32_fa10_20_or0));
  and_gate and_gate_u_csamul_cska32_and11_20(.a(a[11]), .b(b[20]), .out(u_csamul_cska32_and11_20));
  fa fa_u_csamul_cska32_fa11_20_out(.a(u_csamul_cska32_and11_20[0]), .b(u_csamul_cska32_fa12_19_xor1[0]), .cin(u_csamul_cska32_fa11_19_or0[0]), .fa_xor1(u_csamul_cska32_fa11_20_xor1), .fa_or0(u_csamul_cska32_fa11_20_or0));
  and_gate and_gate_u_csamul_cska32_and12_20(.a(a[12]), .b(b[20]), .out(u_csamul_cska32_and12_20));
  fa fa_u_csamul_cska32_fa12_20_out(.a(u_csamul_cska32_and12_20[0]), .b(u_csamul_cska32_fa13_19_xor1[0]), .cin(u_csamul_cska32_fa12_19_or0[0]), .fa_xor1(u_csamul_cska32_fa12_20_xor1), .fa_or0(u_csamul_cska32_fa12_20_or0));
  and_gate and_gate_u_csamul_cska32_and13_20(.a(a[13]), .b(b[20]), .out(u_csamul_cska32_and13_20));
  fa fa_u_csamul_cska32_fa13_20_out(.a(u_csamul_cska32_and13_20[0]), .b(u_csamul_cska32_fa14_19_xor1[0]), .cin(u_csamul_cska32_fa13_19_or0[0]), .fa_xor1(u_csamul_cska32_fa13_20_xor1), .fa_or0(u_csamul_cska32_fa13_20_or0));
  and_gate and_gate_u_csamul_cska32_and14_20(.a(a[14]), .b(b[20]), .out(u_csamul_cska32_and14_20));
  fa fa_u_csamul_cska32_fa14_20_out(.a(u_csamul_cska32_and14_20[0]), .b(u_csamul_cska32_fa15_19_xor1[0]), .cin(u_csamul_cska32_fa14_19_or0[0]), .fa_xor1(u_csamul_cska32_fa14_20_xor1), .fa_or0(u_csamul_cska32_fa14_20_or0));
  and_gate and_gate_u_csamul_cska32_and15_20(.a(a[15]), .b(b[20]), .out(u_csamul_cska32_and15_20));
  fa fa_u_csamul_cska32_fa15_20_out(.a(u_csamul_cska32_and15_20[0]), .b(u_csamul_cska32_fa16_19_xor1[0]), .cin(u_csamul_cska32_fa15_19_or0[0]), .fa_xor1(u_csamul_cska32_fa15_20_xor1), .fa_or0(u_csamul_cska32_fa15_20_or0));
  and_gate and_gate_u_csamul_cska32_and16_20(.a(a[16]), .b(b[20]), .out(u_csamul_cska32_and16_20));
  fa fa_u_csamul_cska32_fa16_20_out(.a(u_csamul_cska32_and16_20[0]), .b(u_csamul_cska32_fa17_19_xor1[0]), .cin(u_csamul_cska32_fa16_19_or0[0]), .fa_xor1(u_csamul_cska32_fa16_20_xor1), .fa_or0(u_csamul_cska32_fa16_20_or0));
  and_gate and_gate_u_csamul_cska32_and17_20(.a(a[17]), .b(b[20]), .out(u_csamul_cska32_and17_20));
  fa fa_u_csamul_cska32_fa17_20_out(.a(u_csamul_cska32_and17_20[0]), .b(u_csamul_cska32_fa18_19_xor1[0]), .cin(u_csamul_cska32_fa17_19_or0[0]), .fa_xor1(u_csamul_cska32_fa17_20_xor1), .fa_or0(u_csamul_cska32_fa17_20_or0));
  and_gate and_gate_u_csamul_cska32_and18_20(.a(a[18]), .b(b[20]), .out(u_csamul_cska32_and18_20));
  fa fa_u_csamul_cska32_fa18_20_out(.a(u_csamul_cska32_and18_20[0]), .b(u_csamul_cska32_fa19_19_xor1[0]), .cin(u_csamul_cska32_fa18_19_or0[0]), .fa_xor1(u_csamul_cska32_fa18_20_xor1), .fa_or0(u_csamul_cska32_fa18_20_or0));
  and_gate and_gate_u_csamul_cska32_and19_20(.a(a[19]), .b(b[20]), .out(u_csamul_cska32_and19_20));
  fa fa_u_csamul_cska32_fa19_20_out(.a(u_csamul_cska32_and19_20[0]), .b(u_csamul_cska32_fa20_19_xor1[0]), .cin(u_csamul_cska32_fa19_19_or0[0]), .fa_xor1(u_csamul_cska32_fa19_20_xor1), .fa_or0(u_csamul_cska32_fa19_20_or0));
  and_gate and_gate_u_csamul_cska32_and20_20(.a(a[20]), .b(b[20]), .out(u_csamul_cska32_and20_20));
  fa fa_u_csamul_cska32_fa20_20_out(.a(u_csamul_cska32_and20_20[0]), .b(u_csamul_cska32_fa21_19_xor1[0]), .cin(u_csamul_cska32_fa20_19_or0[0]), .fa_xor1(u_csamul_cska32_fa20_20_xor1), .fa_or0(u_csamul_cska32_fa20_20_or0));
  and_gate and_gate_u_csamul_cska32_and21_20(.a(a[21]), .b(b[20]), .out(u_csamul_cska32_and21_20));
  fa fa_u_csamul_cska32_fa21_20_out(.a(u_csamul_cska32_and21_20[0]), .b(u_csamul_cska32_fa22_19_xor1[0]), .cin(u_csamul_cska32_fa21_19_or0[0]), .fa_xor1(u_csamul_cska32_fa21_20_xor1), .fa_or0(u_csamul_cska32_fa21_20_or0));
  and_gate and_gate_u_csamul_cska32_and22_20(.a(a[22]), .b(b[20]), .out(u_csamul_cska32_and22_20));
  fa fa_u_csamul_cska32_fa22_20_out(.a(u_csamul_cska32_and22_20[0]), .b(u_csamul_cska32_fa23_19_xor1[0]), .cin(u_csamul_cska32_fa22_19_or0[0]), .fa_xor1(u_csamul_cska32_fa22_20_xor1), .fa_or0(u_csamul_cska32_fa22_20_or0));
  and_gate and_gate_u_csamul_cska32_and23_20(.a(a[23]), .b(b[20]), .out(u_csamul_cska32_and23_20));
  fa fa_u_csamul_cska32_fa23_20_out(.a(u_csamul_cska32_and23_20[0]), .b(u_csamul_cska32_fa24_19_xor1[0]), .cin(u_csamul_cska32_fa23_19_or0[0]), .fa_xor1(u_csamul_cska32_fa23_20_xor1), .fa_or0(u_csamul_cska32_fa23_20_or0));
  and_gate and_gate_u_csamul_cska32_and24_20(.a(a[24]), .b(b[20]), .out(u_csamul_cska32_and24_20));
  fa fa_u_csamul_cska32_fa24_20_out(.a(u_csamul_cska32_and24_20[0]), .b(u_csamul_cska32_fa25_19_xor1[0]), .cin(u_csamul_cska32_fa24_19_or0[0]), .fa_xor1(u_csamul_cska32_fa24_20_xor1), .fa_or0(u_csamul_cska32_fa24_20_or0));
  and_gate and_gate_u_csamul_cska32_and25_20(.a(a[25]), .b(b[20]), .out(u_csamul_cska32_and25_20));
  fa fa_u_csamul_cska32_fa25_20_out(.a(u_csamul_cska32_and25_20[0]), .b(u_csamul_cska32_fa26_19_xor1[0]), .cin(u_csamul_cska32_fa25_19_or0[0]), .fa_xor1(u_csamul_cska32_fa25_20_xor1), .fa_or0(u_csamul_cska32_fa25_20_or0));
  and_gate and_gate_u_csamul_cska32_and26_20(.a(a[26]), .b(b[20]), .out(u_csamul_cska32_and26_20));
  fa fa_u_csamul_cska32_fa26_20_out(.a(u_csamul_cska32_and26_20[0]), .b(u_csamul_cska32_fa27_19_xor1[0]), .cin(u_csamul_cska32_fa26_19_or0[0]), .fa_xor1(u_csamul_cska32_fa26_20_xor1), .fa_or0(u_csamul_cska32_fa26_20_or0));
  and_gate and_gate_u_csamul_cska32_and27_20(.a(a[27]), .b(b[20]), .out(u_csamul_cska32_and27_20));
  fa fa_u_csamul_cska32_fa27_20_out(.a(u_csamul_cska32_and27_20[0]), .b(u_csamul_cska32_fa28_19_xor1[0]), .cin(u_csamul_cska32_fa27_19_or0[0]), .fa_xor1(u_csamul_cska32_fa27_20_xor1), .fa_or0(u_csamul_cska32_fa27_20_or0));
  and_gate and_gate_u_csamul_cska32_and28_20(.a(a[28]), .b(b[20]), .out(u_csamul_cska32_and28_20));
  fa fa_u_csamul_cska32_fa28_20_out(.a(u_csamul_cska32_and28_20[0]), .b(u_csamul_cska32_fa29_19_xor1[0]), .cin(u_csamul_cska32_fa28_19_or0[0]), .fa_xor1(u_csamul_cska32_fa28_20_xor1), .fa_or0(u_csamul_cska32_fa28_20_or0));
  and_gate and_gate_u_csamul_cska32_and29_20(.a(a[29]), .b(b[20]), .out(u_csamul_cska32_and29_20));
  fa fa_u_csamul_cska32_fa29_20_out(.a(u_csamul_cska32_and29_20[0]), .b(u_csamul_cska32_fa30_19_xor1[0]), .cin(u_csamul_cska32_fa29_19_or0[0]), .fa_xor1(u_csamul_cska32_fa29_20_xor1), .fa_or0(u_csamul_cska32_fa29_20_or0));
  and_gate and_gate_u_csamul_cska32_and30_20(.a(a[30]), .b(b[20]), .out(u_csamul_cska32_and30_20));
  fa fa_u_csamul_cska32_fa30_20_out(.a(u_csamul_cska32_and30_20[0]), .b(u_csamul_cska32_and31_19[0]), .cin(u_csamul_cska32_fa30_19_or0[0]), .fa_xor1(u_csamul_cska32_fa30_20_xor1), .fa_or0(u_csamul_cska32_fa30_20_or0));
  and_gate and_gate_u_csamul_cska32_and31_20(.a(a[31]), .b(b[20]), .out(u_csamul_cska32_and31_20));
  and_gate and_gate_u_csamul_cska32_and0_21(.a(a[0]), .b(b[21]), .out(u_csamul_cska32_and0_21));
  fa fa_u_csamul_cska32_fa0_21_out(.a(u_csamul_cska32_and0_21[0]), .b(u_csamul_cska32_fa1_20_xor1[0]), .cin(u_csamul_cska32_fa0_20_or0[0]), .fa_xor1(u_csamul_cska32_fa0_21_xor1), .fa_or0(u_csamul_cska32_fa0_21_or0));
  and_gate and_gate_u_csamul_cska32_and1_21(.a(a[1]), .b(b[21]), .out(u_csamul_cska32_and1_21));
  fa fa_u_csamul_cska32_fa1_21_out(.a(u_csamul_cska32_and1_21[0]), .b(u_csamul_cska32_fa2_20_xor1[0]), .cin(u_csamul_cska32_fa1_20_or0[0]), .fa_xor1(u_csamul_cska32_fa1_21_xor1), .fa_or0(u_csamul_cska32_fa1_21_or0));
  and_gate and_gate_u_csamul_cska32_and2_21(.a(a[2]), .b(b[21]), .out(u_csamul_cska32_and2_21));
  fa fa_u_csamul_cska32_fa2_21_out(.a(u_csamul_cska32_and2_21[0]), .b(u_csamul_cska32_fa3_20_xor1[0]), .cin(u_csamul_cska32_fa2_20_or0[0]), .fa_xor1(u_csamul_cska32_fa2_21_xor1), .fa_or0(u_csamul_cska32_fa2_21_or0));
  and_gate and_gate_u_csamul_cska32_and3_21(.a(a[3]), .b(b[21]), .out(u_csamul_cska32_and3_21));
  fa fa_u_csamul_cska32_fa3_21_out(.a(u_csamul_cska32_and3_21[0]), .b(u_csamul_cska32_fa4_20_xor1[0]), .cin(u_csamul_cska32_fa3_20_or0[0]), .fa_xor1(u_csamul_cska32_fa3_21_xor1), .fa_or0(u_csamul_cska32_fa3_21_or0));
  and_gate and_gate_u_csamul_cska32_and4_21(.a(a[4]), .b(b[21]), .out(u_csamul_cska32_and4_21));
  fa fa_u_csamul_cska32_fa4_21_out(.a(u_csamul_cska32_and4_21[0]), .b(u_csamul_cska32_fa5_20_xor1[0]), .cin(u_csamul_cska32_fa4_20_or0[0]), .fa_xor1(u_csamul_cska32_fa4_21_xor1), .fa_or0(u_csamul_cska32_fa4_21_or0));
  and_gate and_gate_u_csamul_cska32_and5_21(.a(a[5]), .b(b[21]), .out(u_csamul_cska32_and5_21));
  fa fa_u_csamul_cska32_fa5_21_out(.a(u_csamul_cska32_and5_21[0]), .b(u_csamul_cska32_fa6_20_xor1[0]), .cin(u_csamul_cska32_fa5_20_or0[0]), .fa_xor1(u_csamul_cska32_fa5_21_xor1), .fa_or0(u_csamul_cska32_fa5_21_or0));
  and_gate and_gate_u_csamul_cska32_and6_21(.a(a[6]), .b(b[21]), .out(u_csamul_cska32_and6_21));
  fa fa_u_csamul_cska32_fa6_21_out(.a(u_csamul_cska32_and6_21[0]), .b(u_csamul_cska32_fa7_20_xor1[0]), .cin(u_csamul_cska32_fa6_20_or0[0]), .fa_xor1(u_csamul_cska32_fa6_21_xor1), .fa_or0(u_csamul_cska32_fa6_21_or0));
  and_gate and_gate_u_csamul_cska32_and7_21(.a(a[7]), .b(b[21]), .out(u_csamul_cska32_and7_21));
  fa fa_u_csamul_cska32_fa7_21_out(.a(u_csamul_cska32_and7_21[0]), .b(u_csamul_cska32_fa8_20_xor1[0]), .cin(u_csamul_cska32_fa7_20_or0[0]), .fa_xor1(u_csamul_cska32_fa7_21_xor1), .fa_or0(u_csamul_cska32_fa7_21_or0));
  and_gate and_gate_u_csamul_cska32_and8_21(.a(a[8]), .b(b[21]), .out(u_csamul_cska32_and8_21));
  fa fa_u_csamul_cska32_fa8_21_out(.a(u_csamul_cska32_and8_21[0]), .b(u_csamul_cska32_fa9_20_xor1[0]), .cin(u_csamul_cska32_fa8_20_or0[0]), .fa_xor1(u_csamul_cska32_fa8_21_xor1), .fa_or0(u_csamul_cska32_fa8_21_or0));
  and_gate and_gate_u_csamul_cska32_and9_21(.a(a[9]), .b(b[21]), .out(u_csamul_cska32_and9_21));
  fa fa_u_csamul_cska32_fa9_21_out(.a(u_csamul_cska32_and9_21[0]), .b(u_csamul_cska32_fa10_20_xor1[0]), .cin(u_csamul_cska32_fa9_20_or0[0]), .fa_xor1(u_csamul_cska32_fa9_21_xor1), .fa_or0(u_csamul_cska32_fa9_21_or0));
  and_gate and_gate_u_csamul_cska32_and10_21(.a(a[10]), .b(b[21]), .out(u_csamul_cska32_and10_21));
  fa fa_u_csamul_cska32_fa10_21_out(.a(u_csamul_cska32_and10_21[0]), .b(u_csamul_cska32_fa11_20_xor1[0]), .cin(u_csamul_cska32_fa10_20_or0[0]), .fa_xor1(u_csamul_cska32_fa10_21_xor1), .fa_or0(u_csamul_cska32_fa10_21_or0));
  and_gate and_gate_u_csamul_cska32_and11_21(.a(a[11]), .b(b[21]), .out(u_csamul_cska32_and11_21));
  fa fa_u_csamul_cska32_fa11_21_out(.a(u_csamul_cska32_and11_21[0]), .b(u_csamul_cska32_fa12_20_xor1[0]), .cin(u_csamul_cska32_fa11_20_or0[0]), .fa_xor1(u_csamul_cska32_fa11_21_xor1), .fa_or0(u_csamul_cska32_fa11_21_or0));
  and_gate and_gate_u_csamul_cska32_and12_21(.a(a[12]), .b(b[21]), .out(u_csamul_cska32_and12_21));
  fa fa_u_csamul_cska32_fa12_21_out(.a(u_csamul_cska32_and12_21[0]), .b(u_csamul_cska32_fa13_20_xor1[0]), .cin(u_csamul_cska32_fa12_20_or0[0]), .fa_xor1(u_csamul_cska32_fa12_21_xor1), .fa_or0(u_csamul_cska32_fa12_21_or0));
  and_gate and_gate_u_csamul_cska32_and13_21(.a(a[13]), .b(b[21]), .out(u_csamul_cska32_and13_21));
  fa fa_u_csamul_cska32_fa13_21_out(.a(u_csamul_cska32_and13_21[0]), .b(u_csamul_cska32_fa14_20_xor1[0]), .cin(u_csamul_cska32_fa13_20_or0[0]), .fa_xor1(u_csamul_cska32_fa13_21_xor1), .fa_or0(u_csamul_cska32_fa13_21_or0));
  and_gate and_gate_u_csamul_cska32_and14_21(.a(a[14]), .b(b[21]), .out(u_csamul_cska32_and14_21));
  fa fa_u_csamul_cska32_fa14_21_out(.a(u_csamul_cska32_and14_21[0]), .b(u_csamul_cska32_fa15_20_xor1[0]), .cin(u_csamul_cska32_fa14_20_or0[0]), .fa_xor1(u_csamul_cska32_fa14_21_xor1), .fa_or0(u_csamul_cska32_fa14_21_or0));
  and_gate and_gate_u_csamul_cska32_and15_21(.a(a[15]), .b(b[21]), .out(u_csamul_cska32_and15_21));
  fa fa_u_csamul_cska32_fa15_21_out(.a(u_csamul_cska32_and15_21[0]), .b(u_csamul_cska32_fa16_20_xor1[0]), .cin(u_csamul_cska32_fa15_20_or0[0]), .fa_xor1(u_csamul_cska32_fa15_21_xor1), .fa_or0(u_csamul_cska32_fa15_21_or0));
  and_gate and_gate_u_csamul_cska32_and16_21(.a(a[16]), .b(b[21]), .out(u_csamul_cska32_and16_21));
  fa fa_u_csamul_cska32_fa16_21_out(.a(u_csamul_cska32_and16_21[0]), .b(u_csamul_cska32_fa17_20_xor1[0]), .cin(u_csamul_cska32_fa16_20_or0[0]), .fa_xor1(u_csamul_cska32_fa16_21_xor1), .fa_or0(u_csamul_cska32_fa16_21_or0));
  and_gate and_gate_u_csamul_cska32_and17_21(.a(a[17]), .b(b[21]), .out(u_csamul_cska32_and17_21));
  fa fa_u_csamul_cska32_fa17_21_out(.a(u_csamul_cska32_and17_21[0]), .b(u_csamul_cska32_fa18_20_xor1[0]), .cin(u_csamul_cska32_fa17_20_or0[0]), .fa_xor1(u_csamul_cska32_fa17_21_xor1), .fa_or0(u_csamul_cska32_fa17_21_or0));
  and_gate and_gate_u_csamul_cska32_and18_21(.a(a[18]), .b(b[21]), .out(u_csamul_cska32_and18_21));
  fa fa_u_csamul_cska32_fa18_21_out(.a(u_csamul_cska32_and18_21[0]), .b(u_csamul_cska32_fa19_20_xor1[0]), .cin(u_csamul_cska32_fa18_20_or0[0]), .fa_xor1(u_csamul_cska32_fa18_21_xor1), .fa_or0(u_csamul_cska32_fa18_21_or0));
  and_gate and_gate_u_csamul_cska32_and19_21(.a(a[19]), .b(b[21]), .out(u_csamul_cska32_and19_21));
  fa fa_u_csamul_cska32_fa19_21_out(.a(u_csamul_cska32_and19_21[0]), .b(u_csamul_cska32_fa20_20_xor1[0]), .cin(u_csamul_cska32_fa19_20_or0[0]), .fa_xor1(u_csamul_cska32_fa19_21_xor1), .fa_or0(u_csamul_cska32_fa19_21_or0));
  and_gate and_gate_u_csamul_cska32_and20_21(.a(a[20]), .b(b[21]), .out(u_csamul_cska32_and20_21));
  fa fa_u_csamul_cska32_fa20_21_out(.a(u_csamul_cska32_and20_21[0]), .b(u_csamul_cska32_fa21_20_xor1[0]), .cin(u_csamul_cska32_fa20_20_or0[0]), .fa_xor1(u_csamul_cska32_fa20_21_xor1), .fa_or0(u_csamul_cska32_fa20_21_or0));
  and_gate and_gate_u_csamul_cska32_and21_21(.a(a[21]), .b(b[21]), .out(u_csamul_cska32_and21_21));
  fa fa_u_csamul_cska32_fa21_21_out(.a(u_csamul_cska32_and21_21[0]), .b(u_csamul_cska32_fa22_20_xor1[0]), .cin(u_csamul_cska32_fa21_20_or0[0]), .fa_xor1(u_csamul_cska32_fa21_21_xor1), .fa_or0(u_csamul_cska32_fa21_21_or0));
  and_gate and_gate_u_csamul_cska32_and22_21(.a(a[22]), .b(b[21]), .out(u_csamul_cska32_and22_21));
  fa fa_u_csamul_cska32_fa22_21_out(.a(u_csamul_cska32_and22_21[0]), .b(u_csamul_cska32_fa23_20_xor1[0]), .cin(u_csamul_cska32_fa22_20_or0[0]), .fa_xor1(u_csamul_cska32_fa22_21_xor1), .fa_or0(u_csamul_cska32_fa22_21_or0));
  and_gate and_gate_u_csamul_cska32_and23_21(.a(a[23]), .b(b[21]), .out(u_csamul_cska32_and23_21));
  fa fa_u_csamul_cska32_fa23_21_out(.a(u_csamul_cska32_and23_21[0]), .b(u_csamul_cska32_fa24_20_xor1[0]), .cin(u_csamul_cska32_fa23_20_or0[0]), .fa_xor1(u_csamul_cska32_fa23_21_xor1), .fa_or0(u_csamul_cska32_fa23_21_or0));
  and_gate and_gate_u_csamul_cska32_and24_21(.a(a[24]), .b(b[21]), .out(u_csamul_cska32_and24_21));
  fa fa_u_csamul_cska32_fa24_21_out(.a(u_csamul_cska32_and24_21[0]), .b(u_csamul_cska32_fa25_20_xor1[0]), .cin(u_csamul_cska32_fa24_20_or0[0]), .fa_xor1(u_csamul_cska32_fa24_21_xor1), .fa_or0(u_csamul_cska32_fa24_21_or0));
  and_gate and_gate_u_csamul_cska32_and25_21(.a(a[25]), .b(b[21]), .out(u_csamul_cska32_and25_21));
  fa fa_u_csamul_cska32_fa25_21_out(.a(u_csamul_cska32_and25_21[0]), .b(u_csamul_cska32_fa26_20_xor1[0]), .cin(u_csamul_cska32_fa25_20_or0[0]), .fa_xor1(u_csamul_cska32_fa25_21_xor1), .fa_or0(u_csamul_cska32_fa25_21_or0));
  and_gate and_gate_u_csamul_cska32_and26_21(.a(a[26]), .b(b[21]), .out(u_csamul_cska32_and26_21));
  fa fa_u_csamul_cska32_fa26_21_out(.a(u_csamul_cska32_and26_21[0]), .b(u_csamul_cska32_fa27_20_xor1[0]), .cin(u_csamul_cska32_fa26_20_or0[0]), .fa_xor1(u_csamul_cska32_fa26_21_xor1), .fa_or0(u_csamul_cska32_fa26_21_or0));
  and_gate and_gate_u_csamul_cska32_and27_21(.a(a[27]), .b(b[21]), .out(u_csamul_cska32_and27_21));
  fa fa_u_csamul_cska32_fa27_21_out(.a(u_csamul_cska32_and27_21[0]), .b(u_csamul_cska32_fa28_20_xor1[0]), .cin(u_csamul_cska32_fa27_20_or0[0]), .fa_xor1(u_csamul_cska32_fa27_21_xor1), .fa_or0(u_csamul_cska32_fa27_21_or0));
  and_gate and_gate_u_csamul_cska32_and28_21(.a(a[28]), .b(b[21]), .out(u_csamul_cska32_and28_21));
  fa fa_u_csamul_cska32_fa28_21_out(.a(u_csamul_cska32_and28_21[0]), .b(u_csamul_cska32_fa29_20_xor1[0]), .cin(u_csamul_cska32_fa28_20_or0[0]), .fa_xor1(u_csamul_cska32_fa28_21_xor1), .fa_or0(u_csamul_cska32_fa28_21_or0));
  and_gate and_gate_u_csamul_cska32_and29_21(.a(a[29]), .b(b[21]), .out(u_csamul_cska32_and29_21));
  fa fa_u_csamul_cska32_fa29_21_out(.a(u_csamul_cska32_and29_21[0]), .b(u_csamul_cska32_fa30_20_xor1[0]), .cin(u_csamul_cska32_fa29_20_or0[0]), .fa_xor1(u_csamul_cska32_fa29_21_xor1), .fa_or0(u_csamul_cska32_fa29_21_or0));
  and_gate and_gate_u_csamul_cska32_and30_21(.a(a[30]), .b(b[21]), .out(u_csamul_cska32_and30_21));
  fa fa_u_csamul_cska32_fa30_21_out(.a(u_csamul_cska32_and30_21[0]), .b(u_csamul_cska32_and31_20[0]), .cin(u_csamul_cska32_fa30_20_or0[0]), .fa_xor1(u_csamul_cska32_fa30_21_xor1), .fa_or0(u_csamul_cska32_fa30_21_or0));
  and_gate and_gate_u_csamul_cska32_and31_21(.a(a[31]), .b(b[21]), .out(u_csamul_cska32_and31_21));
  and_gate and_gate_u_csamul_cska32_and0_22(.a(a[0]), .b(b[22]), .out(u_csamul_cska32_and0_22));
  fa fa_u_csamul_cska32_fa0_22_out(.a(u_csamul_cska32_and0_22[0]), .b(u_csamul_cska32_fa1_21_xor1[0]), .cin(u_csamul_cska32_fa0_21_or0[0]), .fa_xor1(u_csamul_cska32_fa0_22_xor1), .fa_or0(u_csamul_cska32_fa0_22_or0));
  and_gate and_gate_u_csamul_cska32_and1_22(.a(a[1]), .b(b[22]), .out(u_csamul_cska32_and1_22));
  fa fa_u_csamul_cska32_fa1_22_out(.a(u_csamul_cska32_and1_22[0]), .b(u_csamul_cska32_fa2_21_xor1[0]), .cin(u_csamul_cska32_fa1_21_or0[0]), .fa_xor1(u_csamul_cska32_fa1_22_xor1), .fa_or0(u_csamul_cska32_fa1_22_or0));
  and_gate and_gate_u_csamul_cska32_and2_22(.a(a[2]), .b(b[22]), .out(u_csamul_cska32_and2_22));
  fa fa_u_csamul_cska32_fa2_22_out(.a(u_csamul_cska32_and2_22[0]), .b(u_csamul_cska32_fa3_21_xor1[0]), .cin(u_csamul_cska32_fa2_21_or0[0]), .fa_xor1(u_csamul_cska32_fa2_22_xor1), .fa_or0(u_csamul_cska32_fa2_22_or0));
  and_gate and_gate_u_csamul_cska32_and3_22(.a(a[3]), .b(b[22]), .out(u_csamul_cska32_and3_22));
  fa fa_u_csamul_cska32_fa3_22_out(.a(u_csamul_cska32_and3_22[0]), .b(u_csamul_cska32_fa4_21_xor1[0]), .cin(u_csamul_cska32_fa3_21_or0[0]), .fa_xor1(u_csamul_cska32_fa3_22_xor1), .fa_or0(u_csamul_cska32_fa3_22_or0));
  and_gate and_gate_u_csamul_cska32_and4_22(.a(a[4]), .b(b[22]), .out(u_csamul_cska32_and4_22));
  fa fa_u_csamul_cska32_fa4_22_out(.a(u_csamul_cska32_and4_22[0]), .b(u_csamul_cska32_fa5_21_xor1[0]), .cin(u_csamul_cska32_fa4_21_or0[0]), .fa_xor1(u_csamul_cska32_fa4_22_xor1), .fa_or0(u_csamul_cska32_fa4_22_or0));
  and_gate and_gate_u_csamul_cska32_and5_22(.a(a[5]), .b(b[22]), .out(u_csamul_cska32_and5_22));
  fa fa_u_csamul_cska32_fa5_22_out(.a(u_csamul_cska32_and5_22[0]), .b(u_csamul_cska32_fa6_21_xor1[0]), .cin(u_csamul_cska32_fa5_21_or0[0]), .fa_xor1(u_csamul_cska32_fa5_22_xor1), .fa_or0(u_csamul_cska32_fa5_22_or0));
  and_gate and_gate_u_csamul_cska32_and6_22(.a(a[6]), .b(b[22]), .out(u_csamul_cska32_and6_22));
  fa fa_u_csamul_cska32_fa6_22_out(.a(u_csamul_cska32_and6_22[0]), .b(u_csamul_cska32_fa7_21_xor1[0]), .cin(u_csamul_cska32_fa6_21_or0[0]), .fa_xor1(u_csamul_cska32_fa6_22_xor1), .fa_or0(u_csamul_cska32_fa6_22_or0));
  and_gate and_gate_u_csamul_cska32_and7_22(.a(a[7]), .b(b[22]), .out(u_csamul_cska32_and7_22));
  fa fa_u_csamul_cska32_fa7_22_out(.a(u_csamul_cska32_and7_22[0]), .b(u_csamul_cska32_fa8_21_xor1[0]), .cin(u_csamul_cska32_fa7_21_or0[0]), .fa_xor1(u_csamul_cska32_fa7_22_xor1), .fa_or0(u_csamul_cska32_fa7_22_or0));
  and_gate and_gate_u_csamul_cska32_and8_22(.a(a[8]), .b(b[22]), .out(u_csamul_cska32_and8_22));
  fa fa_u_csamul_cska32_fa8_22_out(.a(u_csamul_cska32_and8_22[0]), .b(u_csamul_cska32_fa9_21_xor1[0]), .cin(u_csamul_cska32_fa8_21_or0[0]), .fa_xor1(u_csamul_cska32_fa8_22_xor1), .fa_or0(u_csamul_cska32_fa8_22_or0));
  and_gate and_gate_u_csamul_cska32_and9_22(.a(a[9]), .b(b[22]), .out(u_csamul_cska32_and9_22));
  fa fa_u_csamul_cska32_fa9_22_out(.a(u_csamul_cska32_and9_22[0]), .b(u_csamul_cska32_fa10_21_xor1[0]), .cin(u_csamul_cska32_fa9_21_or0[0]), .fa_xor1(u_csamul_cska32_fa9_22_xor1), .fa_or0(u_csamul_cska32_fa9_22_or0));
  and_gate and_gate_u_csamul_cska32_and10_22(.a(a[10]), .b(b[22]), .out(u_csamul_cska32_and10_22));
  fa fa_u_csamul_cska32_fa10_22_out(.a(u_csamul_cska32_and10_22[0]), .b(u_csamul_cska32_fa11_21_xor1[0]), .cin(u_csamul_cska32_fa10_21_or0[0]), .fa_xor1(u_csamul_cska32_fa10_22_xor1), .fa_or0(u_csamul_cska32_fa10_22_or0));
  and_gate and_gate_u_csamul_cska32_and11_22(.a(a[11]), .b(b[22]), .out(u_csamul_cska32_and11_22));
  fa fa_u_csamul_cska32_fa11_22_out(.a(u_csamul_cska32_and11_22[0]), .b(u_csamul_cska32_fa12_21_xor1[0]), .cin(u_csamul_cska32_fa11_21_or0[0]), .fa_xor1(u_csamul_cska32_fa11_22_xor1), .fa_or0(u_csamul_cska32_fa11_22_or0));
  and_gate and_gate_u_csamul_cska32_and12_22(.a(a[12]), .b(b[22]), .out(u_csamul_cska32_and12_22));
  fa fa_u_csamul_cska32_fa12_22_out(.a(u_csamul_cska32_and12_22[0]), .b(u_csamul_cska32_fa13_21_xor1[0]), .cin(u_csamul_cska32_fa12_21_or0[0]), .fa_xor1(u_csamul_cska32_fa12_22_xor1), .fa_or0(u_csamul_cska32_fa12_22_or0));
  and_gate and_gate_u_csamul_cska32_and13_22(.a(a[13]), .b(b[22]), .out(u_csamul_cska32_and13_22));
  fa fa_u_csamul_cska32_fa13_22_out(.a(u_csamul_cska32_and13_22[0]), .b(u_csamul_cska32_fa14_21_xor1[0]), .cin(u_csamul_cska32_fa13_21_or0[0]), .fa_xor1(u_csamul_cska32_fa13_22_xor1), .fa_or0(u_csamul_cska32_fa13_22_or0));
  and_gate and_gate_u_csamul_cska32_and14_22(.a(a[14]), .b(b[22]), .out(u_csamul_cska32_and14_22));
  fa fa_u_csamul_cska32_fa14_22_out(.a(u_csamul_cska32_and14_22[0]), .b(u_csamul_cska32_fa15_21_xor1[0]), .cin(u_csamul_cska32_fa14_21_or0[0]), .fa_xor1(u_csamul_cska32_fa14_22_xor1), .fa_or0(u_csamul_cska32_fa14_22_or0));
  and_gate and_gate_u_csamul_cska32_and15_22(.a(a[15]), .b(b[22]), .out(u_csamul_cska32_and15_22));
  fa fa_u_csamul_cska32_fa15_22_out(.a(u_csamul_cska32_and15_22[0]), .b(u_csamul_cska32_fa16_21_xor1[0]), .cin(u_csamul_cska32_fa15_21_or0[0]), .fa_xor1(u_csamul_cska32_fa15_22_xor1), .fa_or0(u_csamul_cska32_fa15_22_or0));
  and_gate and_gate_u_csamul_cska32_and16_22(.a(a[16]), .b(b[22]), .out(u_csamul_cska32_and16_22));
  fa fa_u_csamul_cska32_fa16_22_out(.a(u_csamul_cska32_and16_22[0]), .b(u_csamul_cska32_fa17_21_xor1[0]), .cin(u_csamul_cska32_fa16_21_or0[0]), .fa_xor1(u_csamul_cska32_fa16_22_xor1), .fa_or0(u_csamul_cska32_fa16_22_or0));
  and_gate and_gate_u_csamul_cska32_and17_22(.a(a[17]), .b(b[22]), .out(u_csamul_cska32_and17_22));
  fa fa_u_csamul_cska32_fa17_22_out(.a(u_csamul_cska32_and17_22[0]), .b(u_csamul_cska32_fa18_21_xor1[0]), .cin(u_csamul_cska32_fa17_21_or0[0]), .fa_xor1(u_csamul_cska32_fa17_22_xor1), .fa_or0(u_csamul_cska32_fa17_22_or0));
  and_gate and_gate_u_csamul_cska32_and18_22(.a(a[18]), .b(b[22]), .out(u_csamul_cska32_and18_22));
  fa fa_u_csamul_cska32_fa18_22_out(.a(u_csamul_cska32_and18_22[0]), .b(u_csamul_cska32_fa19_21_xor1[0]), .cin(u_csamul_cska32_fa18_21_or0[0]), .fa_xor1(u_csamul_cska32_fa18_22_xor1), .fa_or0(u_csamul_cska32_fa18_22_or0));
  and_gate and_gate_u_csamul_cska32_and19_22(.a(a[19]), .b(b[22]), .out(u_csamul_cska32_and19_22));
  fa fa_u_csamul_cska32_fa19_22_out(.a(u_csamul_cska32_and19_22[0]), .b(u_csamul_cska32_fa20_21_xor1[0]), .cin(u_csamul_cska32_fa19_21_or0[0]), .fa_xor1(u_csamul_cska32_fa19_22_xor1), .fa_or0(u_csamul_cska32_fa19_22_or0));
  and_gate and_gate_u_csamul_cska32_and20_22(.a(a[20]), .b(b[22]), .out(u_csamul_cska32_and20_22));
  fa fa_u_csamul_cska32_fa20_22_out(.a(u_csamul_cska32_and20_22[0]), .b(u_csamul_cska32_fa21_21_xor1[0]), .cin(u_csamul_cska32_fa20_21_or0[0]), .fa_xor1(u_csamul_cska32_fa20_22_xor1), .fa_or0(u_csamul_cska32_fa20_22_or0));
  and_gate and_gate_u_csamul_cska32_and21_22(.a(a[21]), .b(b[22]), .out(u_csamul_cska32_and21_22));
  fa fa_u_csamul_cska32_fa21_22_out(.a(u_csamul_cska32_and21_22[0]), .b(u_csamul_cska32_fa22_21_xor1[0]), .cin(u_csamul_cska32_fa21_21_or0[0]), .fa_xor1(u_csamul_cska32_fa21_22_xor1), .fa_or0(u_csamul_cska32_fa21_22_or0));
  and_gate and_gate_u_csamul_cska32_and22_22(.a(a[22]), .b(b[22]), .out(u_csamul_cska32_and22_22));
  fa fa_u_csamul_cska32_fa22_22_out(.a(u_csamul_cska32_and22_22[0]), .b(u_csamul_cska32_fa23_21_xor1[0]), .cin(u_csamul_cska32_fa22_21_or0[0]), .fa_xor1(u_csamul_cska32_fa22_22_xor1), .fa_or0(u_csamul_cska32_fa22_22_or0));
  and_gate and_gate_u_csamul_cska32_and23_22(.a(a[23]), .b(b[22]), .out(u_csamul_cska32_and23_22));
  fa fa_u_csamul_cska32_fa23_22_out(.a(u_csamul_cska32_and23_22[0]), .b(u_csamul_cska32_fa24_21_xor1[0]), .cin(u_csamul_cska32_fa23_21_or0[0]), .fa_xor1(u_csamul_cska32_fa23_22_xor1), .fa_or0(u_csamul_cska32_fa23_22_or0));
  and_gate and_gate_u_csamul_cska32_and24_22(.a(a[24]), .b(b[22]), .out(u_csamul_cska32_and24_22));
  fa fa_u_csamul_cska32_fa24_22_out(.a(u_csamul_cska32_and24_22[0]), .b(u_csamul_cska32_fa25_21_xor1[0]), .cin(u_csamul_cska32_fa24_21_or0[0]), .fa_xor1(u_csamul_cska32_fa24_22_xor1), .fa_or0(u_csamul_cska32_fa24_22_or0));
  and_gate and_gate_u_csamul_cska32_and25_22(.a(a[25]), .b(b[22]), .out(u_csamul_cska32_and25_22));
  fa fa_u_csamul_cska32_fa25_22_out(.a(u_csamul_cska32_and25_22[0]), .b(u_csamul_cska32_fa26_21_xor1[0]), .cin(u_csamul_cska32_fa25_21_or0[0]), .fa_xor1(u_csamul_cska32_fa25_22_xor1), .fa_or0(u_csamul_cska32_fa25_22_or0));
  and_gate and_gate_u_csamul_cska32_and26_22(.a(a[26]), .b(b[22]), .out(u_csamul_cska32_and26_22));
  fa fa_u_csamul_cska32_fa26_22_out(.a(u_csamul_cska32_and26_22[0]), .b(u_csamul_cska32_fa27_21_xor1[0]), .cin(u_csamul_cska32_fa26_21_or0[0]), .fa_xor1(u_csamul_cska32_fa26_22_xor1), .fa_or0(u_csamul_cska32_fa26_22_or0));
  and_gate and_gate_u_csamul_cska32_and27_22(.a(a[27]), .b(b[22]), .out(u_csamul_cska32_and27_22));
  fa fa_u_csamul_cska32_fa27_22_out(.a(u_csamul_cska32_and27_22[0]), .b(u_csamul_cska32_fa28_21_xor1[0]), .cin(u_csamul_cska32_fa27_21_or0[0]), .fa_xor1(u_csamul_cska32_fa27_22_xor1), .fa_or0(u_csamul_cska32_fa27_22_or0));
  and_gate and_gate_u_csamul_cska32_and28_22(.a(a[28]), .b(b[22]), .out(u_csamul_cska32_and28_22));
  fa fa_u_csamul_cska32_fa28_22_out(.a(u_csamul_cska32_and28_22[0]), .b(u_csamul_cska32_fa29_21_xor1[0]), .cin(u_csamul_cska32_fa28_21_or0[0]), .fa_xor1(u_csamul_cska32_fa28_22_xor1), .fa_or0(u_csamul_cska32_fa28_22_or0));
  and_gate and_gate_u_csamul_cska32_and29_22(.a(a[29]), .b(b[22]), .out(u_csamul_cska32_and29_22));
  fa fa_u_csamul_cska32_fa29_22_out(.a(u_csamul_cska32_and29_22[0]), .b(u_csamul_cska32_fa30_21_xor1[0]), .cin(u_csamul_cska32_fa29_21_or0[0]), .fa_xor1(u_csamul_cska32_fa29_22_xor1), .fa_or0(u_csamul_cska32_fa29_22_or0));
  and_gate and_gate_u_csamul_cska32_and30_22(.a(a[30]), .b(b[22]), .out(u_csamul_cska32_and30_22));
  fa fa_u_csamul_cska32_fa30_22_out(.a(u_csamul_cska32_and30_22[0]), .b(u_csamul_cska32_and31_21[0]), .cin(u_csamul_cska32_fa30_21_or0[0]), .fa_xor1(u_csamul_cska32_fa30_22_xor1), .fa_or0(u_csamul_cska32_fa30_22_or0));
  and_gate and_gate_u_csamul_cska32_and31_22(.a(a[31]), .b(b[22]), .out(u_csamul_cska32_and31_22));
  and_gate and_gate_u_csamul_cska32_and0_23(.a(a[0]), .b(b[23]), .out(u_csamul_cska32_and0_23));
  fa fa_u_csamul_cska32_fa0_23_out(.a(u_csamul_cska32_and0_23[0]), .b(u_csamul_cska32_fa1_22_xor1[0]), .cin(u_csamul_cska32_fa0_22_or0[0]), .fa_xor1(u_csamul_cska32_fa0_23_xor1), .fa_or0(u_csamul_cska32_fa0_23_or0));
  and_gate and_gate_u_csamul_cska32_and1_23(.a(a[1]), .b(b[23]), .out(u_csamul_cska32_and1_23));
  fa fa_u_csamul_cska32_fa1_23_out(.a(u_csamul_cska32_and1_23[0]), .b(u_csamul_cska32_fa2_22_xor1[0]), .cin(u_csamul_cska32_fa1_22_or0[0]), .fa_xor1(u_csamul_cska32_fa1_23_xor1), .fa_or0(u_csamul_cska32_fa1_23_or0));
  and_gate and_gate_u_csamul_cska32_and2_23(.a(a[2]), .b(b[23]), .out(u_csamul_cska32_and2_23));
  fa fa_u_csamul_cska32_fa2_23_out(.a(u_csamul_cska32_and2_23[0]), .b(u_csamul_cska32_fa3_22_xor1[0]), .cin(u_csamul_cska32_fa2_22_or0[0]), .fa_xor1(u_csamul_cska32_fa2_23_xor1), .fa_or0(u_csamul_cska32_fa2_23_or0));
  and_gate and_gate_u_csamul_cska32_and3_23(.a(a[3]), .b(b[23]), .out(u_csamul_cska32_and3_23));
  fa fa_u_csamul_cska32_fa3_23_out(.a(u_csamul_cska32_and3_23[0]), .b(u_csamul_cska32_fa4_22_xor1[0]), .cin(u_csamul_cska32_fa3_22_or0[0]), .fa_xor1(u_csamul_cska32_fa3_23_xor1), .fa_or0(u_csamul_cska32_fa3_23_or0));
  and_gate and_gate_u_csamul_cska32_and4_23(.a(a[4]), .b(b[23]), .out(u_csamul_cska32_and4_23));
  fa fa_u_csamul_cska32_fa4_23_out(.a(u_csamul_cska32_and4_23[0]), .b(u_csamul_cska32_fa5_22_xor1[0]), .cin(u_csamul_cska32_fa4_22_or0[0]), .fa_xor1(u_csamul_cska32_fa4_23_xor1), .fa_or0(u_csamul_cska32_fa4_23_or0));
  and_gate and_gate_u_csamul_cska32_and5_23(.a(a[5]), .b(b[23]), .out(u_csamul_cska32_and5_23));
  fa fa_u_csamul_cska32_fa5_23_out(.a(u_csamul_cska32_and5_23[0]), .b(u_csamul_cska32_fa6_22_xor1[0]), .cin(u_csamul_cska32_fa5_22_or0[0]), .fa_xor1(u_csamul_cska32_fa5_23_xor1), .fa_or0(u_csamul_cska32_fa5_23_or0));
  and_gate and_gate_u_csamul_cska32_and6_23(.a(a[6]), .b(b[23]), .out(u_csamul_cska32_and6_23));
  fa fa_u_csamul_cska32_fa6_23_out(.a(u_csamul_cska32_and6_23[0]), .b(u_csamul_cska32_fa7_22_xor1[0]), .cin(u_csamul_cska32_fa6_22_or0[0]), .fa_xor1(u_csamul_cska32_fa6_23_xor1), .fa_or0(u_csamul_cska32_fa6_23_or0));
  and_gate and_gate_u_csamul_cska32_and7_23(.a(a[7]), .b(b[23]), .out(u_csamul_cska32_and7_23));
  fa fa_u_csamul_cska32_fa7_23_out(.a(u_csamul_cska32_and7_23[0]), .b(u_csamul_cska32_fa8_22_xor1[0]), .cin(u_csamul_cska32_fa7_22_or0[0]), .fa_xor1(u_csamul_cska32_fa7_23_xor1), .fa_or0(u_csamul_cska32_fa7_23_or0));
  and_gate and_gate_u_csamul_cska32_and8_23(.a(a[8]), .b(b[23]), .out(u_csamul_cska32_and8_23));
  fa fa_u_csamul_cska32_fa8_23_out(.a(u_csamul_cska32_and8_23[0]), .b(u_csamul_cska32_fa9_22_xor1[0]), .cin(u_csamul_cska32_fa8_22_or0[0]), .fa_xor1(u_csamul_cska32_fa8_23_xor1), .fa_or0(u_csamul_cska32_fa8_23_or0));
  and_gate and_gate_u_csamul_cska32_and9_23(.a(a[9]), .b(b[23]), .out(u_csamul_cska32_and9_23));
  fa fa_u_csamul_cska32_fa9_23_out(.a(u_csamul_cska32_and9_23[0]), .b(u_csamul_cska32_fa10_22_xor1[0]), .cin(u_csamul_cska32_fa9_22_or0[0]), .fa_xor1(u_csamul_cska32_fa9_23_xor1), .fa_or0(u_csamul_cska32_fa9_23_or0));
  and_gate and_gate_u_csamul_cska32_and10_23(.a(a[10]), .b(b[23]), .out(u_csamul_cska32_and10_23));
  fa fa_u_csamul_cska32_fa10_23_out(.a(u_csamul_cska32_and10_23[0]), .b(u_csamul_cska32_fa11_22_xor1[0]), .cin(u_csamul_cska32_fa10_22_or0[0]), .fa_xor1(u_csamul_cska32_fa10_23_xor1), .fa_or0(u_csamul_cska32_fa10_23_or0));
  and_gate and_gate_u_csamul_cska32_and11_23(.a(a[11]), .b(b[23]), .out(u_csamul_cska32_and11_23));
  fa fa_u_csamul_cska32_fa11_23_out(.a(u_csamul_cska32_and11_23[0]), .b(u_csamul_cska32_fa12_22_xor1[0]), .cin(u_csamul_cska32_fa11_22_or0[0]), .fa_xor1(u_csamul_cska32_fa11_23_xor1), .fa_or0(u_csamul_cska32_fa11_23_or0));
  and_gate and_gate_u_csamul_cska32_and12_23(.a(a[12]), .b(b[23]), .out(u_csamul_cska32_and12_23));
  fa fa_u_csamul_cska32_fa12_23_out(.a(u_csamul_cska32_and12_23[0]), .b(u_csamul_cska32_fa13_22_xor1[0]), .cin(u_csamul_cska32_fa12_22_or0[0]), .fa_xor1(u_csamul_cska32_fa12_23_xor1), .fa_or0(u_csamul_cska32_fa12_23_or0));
  and_gate and_gate_u_csamul_cska32_and13_23(.a(a[13]), .b(b[23]), .out(u_csamul_cska32_and13_23));
  fa fa_u_csamul_cska32_fa13_23_out(.a(u_csamul_cska32_and13_23[0]), .b(u_csamul_cska32_fa14_22_xor1[0]), .cin(u_csamul_cska32_fa13_22_or0[0]), .fa_xor1(u_csamul_cska32_fa13_23_xor1), .fa_or0(u_csamul_cska32_fa13_23_or0));
  and_gate and_gate_u_csamul_cska32_and14_23(.a(a[14]), .b(b[23]), .out(u_csamul_cska32_and14_23));
  fa fa_u_csamul_cska32_fa14_23_out(.a(u_csamul_cska32_and14_23[0]), .b(u_csamul_cska32_fa15_22_xor1[0]), .cin(u_csamul_cska32_fa14_22_or0[0]), .fa_xor1(u_csamul_cska32_fa14_23_xor1), .fa_or0(u_csamul_cska32_fa14_23_or0));
  and_gate and_gate_u_csamul_cska32_and15_23(.a(a[15]), .b(b[23]), .out(u_csamul_cska32_and15_23));
  fa fa_u_csamul_cska32_fa15_23_out(.a(u_csamul_cska32_and15_23[0]), .b(u_csamul_cska32_fa16_22_xor1[0]), .cin(u_csamul_cska32_fa15_22_or0[0]), .fa_xor1(u_csamul_cska32_fa15_23_xor1), .fa_or0(u_csamul_cska32_fa15_23_or0));
  and_gate and_gate_u_csamul_cska32_and16_23(.a(a[16]), .b(b[23]), .out(u_csamul_cska32_and16_23));
  fa fa_u_csamul_cska32_fa16_23_out(.a(u_csamul_cska32_and16_23[0]), .b(u_csamul_cska32_fa17_22_xor1[0]), .cin(u_csamul_cska32_fa16_22_or0[0]), .fa_xor1(u_csamul_cska32_fa16_23_xor1), .fa_or0(u_csamul_cska32_fa16_23_or0));
  and_gate and_gate_u_csamul_cska32_and17_23(.a(a[17]), .b(b[23]), .out(u_csamul_cska32_and17_23));
  fa fa_u_csamul_cska32_fa17_23_out(.a(u_csamul_cska32_and17_23[0]), .b(u_csamul_cska32_fa18_22_xor1[0]), .cin(u_csamul_cska32_fa17_22_or0[0]), .fa_xor1(u_csamul_cska32_fa17_23_xor1), .fa_or0(u_csamul_cska32_fa17_23_or0));
  and_gate and_gate_u_csamul_cska32_and18_23(.a(a[18]), .b(b[23]), .out(u_csamul_cska32_and18_23));
  fa fa_u_csamul_cska32_fa18_23_out(.a(u_csamul_cska32_and18_23[0]), .b(u_csamul_cska32_fa19_22_xor1[0]), .cin(u_csamul_cska32_fa18_22_or0[0]), .fa_xor1(u_csamul_cska32_fa18_23_xor1), .fa_or0(u_csamul_cska32_fa18_23_or0));
  and_gate and_gate_u_csamul_cska32_and19_23(.a(a[19]), .b(b[23]), .out(u_csamul_cska32_and19_23));
  fa fa_u_csamul_cska32_fa19_23_out(.a(u_csamul_cska32_and19_23[0]), .b(u_csamul_cska32_fa20_22_xor1[0]), .cin(u_csamul_cska32_fa19_22_or0[0]), .fa_xor1(u_csamul_cska32_fa19_23_xor1), .fa_or0(u_csamul_cska32_fa19_23_or0));
  and_gate and_gate_u_csamul_cska32_and20_23(.a(a[20]), .b(b[23]), .out(u_csamul_cska32_and20_23));
  fa fa_u_csamul_cska32_fa20_23_out(.a(u_csamul_cska32_and20_23[0]), .b(u_csamul_cska32_fa21_22_xor1[0]), .cin(u_csamul_cska32_fa20_22_or0[0]), .fa_xor1(u_csamul_cska32_fa20_23_xor1), .fa_or0(u_csamul_cska32_fa20_23_or0));
  and_gate and_gate_u_csamul_cska32_and21_23(.a(a[21]), .b(b[23]), .out(u_csamul_cska32_and21_23));
  fa fa_u_csamul_cska32_fa21_23_out(.a(u_csamul_cska32_and21_23[0]), .b(u_csamul_cska32_fa22_22_xor1[0]), .cin(u_csamul_cska32_fa21_22_or0[0]), .fa_xor1(u_csamul_cska32_fa21_23_xor1), .fa_or0(u_csamul_cska32_fa21_23_or0));
  and_gate and_gate_u_csamul_cska32_and22_23(.a(a[22]), .b(b[23]), .out(u_csamul_cska32_and22_23));
  fa fa_u_csamul_cska32_fa22_23_out(.a(u_csamul_cska32_and22_23[0]), .b(u_csamul_cska32_fa23_22_xor1[0]), .cin(u_csamul_cska32_fa22_22_or0[0]), .fa_xor1(u_csamul_cska32_fa22_23_xor1), .fa_or0(u_csamul_cska32_fa22_23_or0));
  and_gate and_gate_u_csamul_cska32_and23_23(.a(a[23]), .b(b[23]), .out(u_csamul_cska32_and23_23));
  fa fa_u_csamul_cska32_fa23_23_out(.a(u_csamul_cska32_and23_23[0]), .b(u_csamul_cska32_fa24_22_xor1[0]), .cin(u_csamul_cska32_fa23_22_or0[0]), .fa_xor1(u_csamul_cska32_fa23_23_xor1), .fa_or0(u_csamul_cska32_fa23_23_or0));
  and_gate and_gate_u_csamul_cska32_and24_23(.a(a[24]), .b(b[23]), .out(u_csamul_cska32_and24_23));
  fa fa_u_csamul_cska32_fa24_23_out(.a(u_csamul_cska32_and24_23[0]), .b(u_csamul_cska32_fa25_22_xor1[0]), .cin(u_csamul_cska32_fa24_22_or0[0]), .fa_xor1(u_csamul_cska32_fa24_23_xor1), .fa_or0(u_csamul_cska32_fa24_23_or0));
  and_gate and_gate_u_csamul_cska32_and25_23(.a(a[25]), .b(b[23]), .out(u_csamul_cska32_and25_23));
  fa fa_u_csamul_cska32_fa25_23_out(.a(u_csamul_cska32_and25_23[0]), .b(u_csamul_cska32_fa26_22_xor1[0]), .cin(u_csamul_cska32_fa25_22_or0[0]), .fa_xor1(u_csamul_cska32_fa25_23_xor1), .fa_or0(u_csamul_cska32_fa25_23_or0));
  and_gate and_gate_u_csamul_cska32_and26_23(.a(a[26]), .b(b[23]), .out(u_csamul_cska32_and26_23));
  fa fa_u_csamul_cska32_fa26_23_out(.a(u_csamul_cska32_and26_23[0]), .b(u_csamul_cska32_fa27_22_xor1[0]), .cin(u_csamul_cska32_fa26_22_or0[0]), .fa_xor1(u_csamul_cska32_fa26_23_xor1), .fa_or0(u_csamul_cska32_fa26_23_or0));
  and_gate and_gate_u_csamul_cska32_and27_23(.a(a[27]), .b(b[23]), .out(u_csamul_cska32_and27_23));
  fa fa_u_csamul_cska32_fa27_23_out(.a(u_csamul_cska32_and27_23[0]), .b(u_csamul_cska32_fa28_22_xor1[0]), .cin(u_csamul_cska32_fa27_22_or0[0]), .fa_xor1(u_csamul_cska32_fa27_23_xor1), .fa_or0(u_csamul_cska32_fa27_23_or0));
  and_gate and_gate_u_csamul_cska32_and28_23(.a(a[28]), .b(b[23]), .out(u_csamul_cska32_and28_23));
  fa fa_u_csamul_cska32_fa28_23_out(.a(u_csamul_cska32_and28_23[0]), .b(u_csamul_cska32_fa29_22_xor1[0]), .cin(u_csamul_cska32_fa28_22_or0[0]), .fa_xor1(u_csamul_cska32_fa28_23_xor1), .fa_or0(u_csamul_cska32_fa28_23_or0));
  and_gate and_gate_u_csamul_cska32_and29_23(.a(a[29]), .b(b[23]), .out(u_csamul_cska32_and29_23));
  fa fa_u_csamul_cska32_fa29_23_out(.a(u_csamul_cska32_and29_23[0]), .b(u_csamul_cska32_fa30_22_xor1[0]), .cin(u_csamul_cska32_fa29_22_or0[0]), .fa_xor1(u_csamul_cska32_fa29_23_xor1), .fa_or0(u_csamul_cska32_fa29_23_or0));
  and_gate and_gate_u_csamul_cska32_and30_23(.a(a[30]), .b(b[23]), .out(u_csamul_cska32_and30_23));
  fa fa_u_csamul_cska32_fa30_23_out(.a(u_csamul_cska32_and30_23[0]), .b(u_csamul_cska32_and31_22[0]), .cin(u_csamul_cska32_fa30_22_or0[0]), .fa_xor1(u_csamul_cska32_fa30_23_xor1), .fa_or0(u_csamul_cska32_fa30_23_or0));
  and_gate and_gate_u_csamul_cska32_and31_23(.a(a[31]), .b(b[23]), .out(u_csamul_cska32_and31_23));
  and_gate and_gate_u_csamul_cska32_and0_24(.a(a[0]), .b(b[24]), .out(u_csamul_cska32_and0_24));
  fa fa_u_csamul_cska32_fa0_24_out(.a(u_csamul_cska32_and0_24[0]), .b(u_csamul_cska32_fa1_23_xor1[0]), .cin(u_csamul_cska32_fa0_23_or0[0]), .fa_xor1(u_csamul_cska32_fa0_24_xor1), .fa_or0(u_csamul_cska32_fa0_24_or0));
  and_gate and_gate_u_csamul_cska32_and1_24(.a(a[1]), .b(b[24]), .out(u_csamul_cska32_and1_24));
  fa fa_u_csamul_cska32_fa1_24_out(.a(u_csamul_cska32_and1_24[0]), .b(u_csamul_cska32_fa2_23_xor1[0]), .cin(u_csamul_cska32_fa1_23_or0[0]), .fa_xor1(u_csamul_cska32_fa1_24_xor1), .fa_or0(u_csamul_cska32_fa1_24_or0));
  and_gate and_gate_u_csamul_cska32_and2_24(.a(a[2]), .b(b[24]), .out(u_csamul_cska32_and2_24));
  fa fa_u_csamul_cska32_fa2_24_out(.a(u_csamul_cska32_and2_24[0]), .b(u_csamul_cska32_fa3_23_xor1[0]), .cin(u_csamul_cska32_fa2_23_or0[0]), .fa_xor1(u_csamul_cska32_fa2_24_xor1), .fa_or0(u_csamul_cska32_fa2_24_or0));
  and_gate and_gate_u_csamul_cska32_and3_24(.a(a[3]), .b(b[24]), .out(u_csamul_cska32_and3_24));
  fa fa_u_csamul_cska32_fa3_24_out(.a(u_csamul_cska32_and3_24[0]), .b(u_csamul_cska32_fa4_23_xor1[0]), .cin(u_csamul_cska32_fa3_23_or0[0]), .fa_xor1(u_csamul_cska32_fa3_24_xor1), .fa_or0(u_csamul_cska32_fa3_24_or0));
  and_gate and_gate_u_csamul_cska32_and4_24(.a(a[4]), .b(b[24]), .out(u_csamul_cska32_and4_24));
  fa fa_u_csamul_cska32_fa4_24_out(.a(u_csamul_cska32_and4_24[0]), .b(u_csamul_cska32_fa5_23_xor1[0]), .cin(u_csamul_cska32_fa4_23_or0[0]), .fa_xor1(u_csamul_cska32_fa4_24_xor1), .fa_or0(u_csamul_cska32_fa4_24_or0));
  and_gate and_gate_u_csamul_cska32_and5_24(.a(a[5]), .b(b[24]), .out(u_csamul_cska32_and5_24));
  fa fa_u_csamul_cska32_fa5_24_out(.a(u_csamul_cska32_and5_24[0]), .b(u_csamul_cska32_fa6_23_xor1[0]), .cin(u_csamul_cska32_fa5_23_or0[0]), .fa_xor1(u_csamul_cska32_fa5_24_xor1), .fa_or0(u_csamul_cska32_fa5_24_or0));
  and_gate and_gate_u_csamul_cska32_and6_24(.a(a[6]), .b(b[24]), .out(u_csamul_cska32_and6_24));
  fa fa_u_csamul_cska32_fa6_24_out(.a(u_csamul_cska32_and6_24[0]), .b(u_csamul_cska32_fa7_23_xor1[0]), .cin(u_csamul_cska32_fa6_23_or0[0]), .fa_xor1(u_csamul_cska32_fa6_24_xor1), .fa_or0(u_csamul_cska32_fa6_24_or0));
  and_gate and_gate_u_csamul_cska32_and7_24(.a(a[7]), .b(b[24]), .out(u_csamul_cska32_and7_24));
  fa fa_u_csamul_cska32_fa7_24_out(.a(u_csamul_cska32_and7_24[0]), .b(u_csamul_cska32_fa8_23_xor1[0]), .cin(u_csamul_cska32_fa7_23_or0[0]), .fa_xor1(u_csamul_cska32_fa7_24_xor1), .fa_or0(u_csamul_cska32_fa7_24_or0));
  and_gate and_gate_u_csamul_cska32_and8_24(.a(a[8]), .b(b[24]), .out(u_csamul_cska32_and8_24));
  fa fa_u_csamul_cska32_fa8_24_out(.a(u_csamul_cska32_and8_24[0]), .b(u_csamul_cska32_fa9_23_xor1[0]), .cin(u_csamul_cska32_fa8_23_or0[0]), .fa_xor1(u_csamul_cska32_fa8_24_xor1), .fa_or0(u_csamul_cska32_fa8_24_or0));
  and_gate and_gate_u_csamul_cska32_and9_24(.a(a[9]), .b(b[24]), .out(u_csamul_cska32_and9_24));
  fa fa_u_csamul_cska32_fa9_24_out(.a(u_csamul_cska32_and9_24[0]), .b(u_csamul_cska32_fa10_23_xor1[0]), .cin(u_csamul_cska32_fa9_23_or0[0]), .fa_xor1(u_csamul_cska32_fa9_24_xor1), .fa_or0(u_csamul_cska32_fa9_24_or0));
  and_gate and_gate_u_csamul_cska32_and10_24(.a(a[10]), .b(b[24]), .out(u_csamul_cska32_and10_24));
  fa fa_u_csamul_cska32_fa10_24_out(.a(u_csamul_cska32_and10_24[0]), .b(u_csamul_cska32_fa11_23_xor1[0]), .cin(u_csamul_cska32_fa10_23_or0[0]), .fa_xor1(u_csamul_cska32_fa10_24_xor1), .fa_or0(u_csamul_cska32_fa10_24_or0));
  and_gate and_gate_u_csamul_cska32_and11_24(.a(a[11]), .b(b[24]), .out(u_csamul_cska32_and11_24));
  fa fa_u_csamul_cska32_fa11_24_out(.a(u_csamul_cska32_and11_24[0]), .b(u_csamul_cska32_fa12_23_xor1[0]), .cin(u_csamul_cska32_fa11_23_or0[0]), .fa_xor1(u_csamul_cska32_fa11_24_xor1), .fa_or0(u_csamul_cska32_fa11_24_or0));
  and_gate and_gate_u_csamul_cska32_and12_24(.a(a[12]), .b(b[24]), .out(u_csamul_cska32_and12_24));
  fa fa_u_csamul_cska32_fa12_24_out(.a(u_csamul_cska32_and12_24[0]), .b(u_csamul_cska32_fa13_23_xor1[0]), .cin(u_csamul_cska32_fa12_23_or0[0]), .fa_xor1(u_csamul_cska32_fa12_24_xor1), .fa_or0(u_csamul_cska32_fa12_24_or0));
  and_gate and_gate_u_csamul_cska32_and13_24(.a(a[13]), .b(b[24]), .out(u_csamul_cska32_and13_24));
  fa fa_u_csamul_cska32_fa13_24_out(.a(u_csamul_cska32_and13_24[0]), .b(u_csamul_cska32_fa14_23_xor1[0]), .cin(u_csamul_cska32_fa13_23_or0[0]), .fa_xor1(u_csamul_cska32_fa13_24_xor1), .fa_or0(u_csamul_cska32_fa13_24_or0));
  and_gate and_gate_u_csamul_cska32_and14_24(.a(a[14]), .b(b[24]), .out(u_csamul_cska32_and14_24));
  fa fa_u_csamul_cska32_fa14_24_out(.a(u_csamul_cska32_and14_24[0]), .b(u_csamul_cska32_fa15_23_xor1[0]), .cin(u_csamul_cska32_fa14_23_or0[0]), .fa_xor1(u_csamul_cska32_fa14_24_xor1), .fa_or0(u_csamul_cska32_fa14_24_or0));
  and_gate and_gate_u_csamul_cska32_and15_24(.a(a[15]), .b(b[24]), .out(u_csamul_cska32_and15_24));
  fa fa_u_csamul_cska32_fa15_24_out(.a(u_csamul_cska32_and15_24[0]), .b(u_csamul_cska32_fa16_23_xor1[0]), .cin(u_csamul_cska32_fa15_23_or0[0]), .fa_xor1(u_csamul_cska32_fa15_24_xor1), .fa_or0(u_csamul_cska32_fa15_24_or0));
  and_gate and_gate_u_csamul_cska32_and16_24(.a(a[16]), .b(b[24]), .out(u_csamul_cska32_and16_24));
  fa fa_u_csamul_cska32_fa16_24_out(.a(u_csamul_cska32_and16_24[0]), .b(u_csamul_cska32_fa17_23_xor1[0]), .cin(u_csamul_cska32_fa16_23_or0[0]), .fa_xor1(u_csamul_cska32_fa16_24_xor1), .fa_or0(u_csamul_cska32_fa16_24_or0));
  and_gate and_gate_u_csamul_cska32_and17_24(.a(a[17]), .b(b[24]), .out(u_csamul_cska32_and17_24));
  fa fa_u_csamul_cska32_fa17_24_out(.a(u_csamul_cska32_and17_24[0]), .b(u_csamul_cska32_fa18_23_xor1[0]), .cin(u_csamul_cska32_fa17_23_or0[0]), .fa_xor1(u_csamul_cska32_fa17_24_xor1), .fa_or0(u_csamul_cska32_fa17_24_or0));
  and_gate and_gate_u_csamul_cska32_and18_24(.a(a[18]), .b(b[24]), .out(u_csamul_cska32_and18_24));
  fa fa_u_csamul_cska32_fa18_24_out(.a(u_csamul_cska32_and18_24[0]), .b(u_csamul_cska32_fa19_23_xor1[0]), .cin(u_csamul_cska32_fa18_23_or0[0]), .fa_xor1(u_csamul_cska32_fa18_24_xor1), .fa_or0(u_csamul_cska32_fa18_24_or0));
  and_gate and_gate_u_csamul_cska32_and19_24(.a(a[19]), .b(b[24]), .out(u_csamul_cska32_and19_24));
  fa fa_u_csamul_cska32_fa19_24_out(.a(u_csamul_cska32_and19_24[0]), .b(u_csamul_cska32_fa20_23_xor1[0]), .cin(u_csamul_cska32_fa19_23_or0[0]), .fa_xor1(u_csamul_cska32_fa19_24_xor1), .fa_or0(u_csamul_cska32_fa19_24_or0));
  and_gate and_gate_u_csamul_cska32_and20_24(.a(a[20]), .b(b[24]), .out(u_csamul_cska32_and20_24));
  fa fa_u_csamul_cska32_fa20_24_out(.a(u_csamul_cska32_and20_24[0]), .b(u_csamul_cska32_fa21_23_xor1[0]), .cin(u_csamul_cska32_fa20_23_or0[0]), .fa_xor1(u_csamul_cska32_fa20_24_xor1), .fa_or0(u_csamul_cska32_fa20_24_or0));
  and_gate and_gate_u_csamul_cska32_and21_24(.a(a[21]), .b(b[24]), .out(u_csamul_cska32_and21_24));
  fa fa_u_csamul_cska32_fa21_24_out(.a(u_csamul_cska32_and21_24[0]), .b(u_csamul_cska32_fa22_23_xor1[0]), .cin(u_csamul_cska32_fa21_23_or0[0]), .fa_xor1(u_csamul_cska32_fa21_24_xor1), .fa_or0(u_csamul_cska32_fa21_24_or0));
  and_gate and_gate_u_csamul_cska32_and22_24(.a(a[22]), .b(b[24]), .out(u_csamul_cska32_and22_24));
  fa fa_u_csamul_cska32_fa22_24_out(.a(u_csamul_cska32_and22_24[0]), .b(u_csamul_cska32_fa23_23_xor1[0]), .cin(u_csamul_cska32_fa22_23_or0[0]), .fa_xor1(u_csamul_cska32_fa22_24_xor1), .fa_or0(u_csamul_cska32_fa22_24_or0));
  and_gate and_gate_u_csamul_cska32_and23_24(.a(a[23]), .b(b[24]), .out(u_csamul_cska32_and23_24));
  fa fa_u_csamul_cska32_fa23_24_out(.a(u_csamul_cska32_and23_24[0]), .b(u_csamul_cska32_fa24_23_xor1[0]), .cin(u_csamul_cska32_fa23_23_or0[0]), .fa_xor1(u_csamul_cska32_fa23_24_xor1), .fa_or0(u_csamul_cska32_fa23_24_or0));
  and_gate and_gate_u_csamul_cska32_and24_24(.a(a[24]), .b(b[24]), .out(u_csamul_cska32_and24_24));
  fa fa_u_csamul_cska32_fa24_24_out(.a(u_csamul_cska32_and24_24[0]), .b(u_csamul_cska32_fa25_23_xor1[0]), .cin(u_csamul_cska32_fa24_23_or0[0]), .fa_xor1(u_csamul_cska32_fa24_24_xor1), .fa_or0(u_csamul_cska32_fa24_24_or0));
  and_gate and_gate_u_csamul_cska32_and25_24(.a(a[25]), .b(b[24]), .out(u_csamul_cska32_and25_24));
  fa fa_u_csamul_cska32_fa25_24_out(.a(u_csamul_cska32_and25_24[0]), .b(u_csamul_cska32_fa26_23_xor1[0]), .cin(u_csamul_cska32_fa25_23_or0[0]), .fa_xor1(u_csamul_cska32_fa25_24_xor1), .fa_or0(u_csamul_cska32_fa25_24_or0));
  and_gate and_gate_u_csamul_cska32_and26_24(.a(a[26]), .b(b[24]), .out(u_csamul_cska32_and26_24));
  fa fa_u_csamul_cska32_fa26_24_out(.a(u_csamul_cska32_and26_24[0]), .b(u_csamul_cska32_fa27_23_xor1[0]), .cin(u_csamul_cska32_fa26_23_or0[0]), .fa_xor1(u_csamul_cska32_fa26_24_xor1), .fa_or0(u_csamul_cska32_fa26_24_or0));
  and_gate and_gate_u_csamul_cska32_and27_24(.a(a[27]), .b(b[24]), .out(u_csamul_cska32_and27_24));
  fa fa_u_csamul_cska32_fa27_24_out(.a(u_csamul_cska32_and27_24[0]), .b(u_csamul_cska32_fa28_23_xor1[0]), .cin(u_csamul_cska32_fa27_23_or0[0]), .fa_xor1(u_csamul_cska32_fa27_24_xor1), .fa_or0(u_csamul_cska32_fa27_24_or0));
  and_gate and_gate_u_csamul_cska32_and28_24(.a(a[28]), .b(b[24]), .out(u_csamul_cska32_and28_24));
  fa fa_u_csamul_cska32_fa28_24_out(.a(u_csamul_cska32_and28_24[0]), .b(u_csamul_cska32_fa29_23_xor1[0]), .cin(u_csamul_cska32_fa28_23_or0[0]), .fa_xor1(u_csamul_cska32_fa28_24_xor1), .fa_or0(u_csamul_cska32_fa28_24_or0));
  and_gate and_gate_u_csamul_cska32_and29_24(.a(a[29]), .b(b[24]), .out(u_csamul_cska32_and29_24));
  fa fa_u_csamul_cska32_fa29_24_out(.a(u_csamul_cska32_and29_24[0]), .b(u_csamul_cska32_fa30_23_xor1[0]), .cin(u_csamul_cska32_fa29_23_or0[0]), .fa_xor1(u_csamul_cska32_fa29_24_xor1), .fa_or0(u_csamul_cska32_fa29_24_or0));
  and_gate and_gate_u_csamul_cska32_and30_24(.a(a[30]), .b(b[24]), .out(u_csamul_cska32_and30_24));
  fa fa_u_csamul_cska32_fa30_24_out(.a(u_csamul_cska32_and30_24[0]), .b(u_csamul_cska32_and31_23[0]), .cin(u_csamul_cska32_fa30_23_or0[0]), .fa_xor1(u_csamul_cska32_fa30_24_xor1), .fa_or0(u_csamul_cska32_fa30_24_or0));
  and_gate and_gate_u_csamul_cska32_and31_24(.a(a[31]), .b(b[24]), .out(u_csamul_cska32_and31_24));
  and_gate and_gate_u_csamul_cska32_and0_25(.a(a[0]), .b(b[25]), .out(u_csamul_cska32_and0_25));
  fa fa_u_csamul_cska32_fa0_25_out(.a(u_csamul_cska32_and0_25[0]), .b(u_csamul_cska32_fa1_24_xor1[0]), .cin(u_csamul_cska32_fa0_24_or0[0]), .fa_xor1(u_csamul_cska32_fa0_25_xor1), .fa_or0(u_csamul_cska32_fa0_25_or0));
  and_gate and_gate_u_csamul_cska32_and1_25(.a(a[1]), .b(b[25]), .out(u_csamul_cska32_and1_25));
  fa fa_u_csamul_cska32_fa1_25_out(.a(u_csamul_cska32_and1_25[0]), .b(u_csamul_cska32_fa2_24_xor1[0]), .cin(u_csamul_cska32_fa1_24_or0[0]), .fa_xor1(u_csamul_cska32_fa1_25_xor1), .fa_or0(u_csamul_cska32_fa1_25_or0));
  and_gate and_gate_u_csamul_cska32_and2_25(.a(a[2]), .b(b[25]), .out(u_csamul_cska32_and2_25));
  fa fa_u_csamul_cska32_fa2_25_out(.a(u_csamul_cska32_and2_25[0]), .b(u_csamul_cska32_fa3_24_xor1[0]), .cin(u_csamul_cska32_fa2_24_or0[0]), .fa_xor1(u_csamul_cska32_fa2_25_xor1), .fa_or0(u_csamul_cska32_fa2_25_or0));
  and_gate and_gate_u_csamul_cska32_and3_25(.a(a[3]), .b(b[25]), .out(u_csamul_cska32_and3_25));
  fa fa_u_csamul_cska32_fa3_25_out(.a(u_csamul_cska32_and3_25[0]), .b(u_csamul_cska32_fa4_24_xor1[0]), .cin(u_csamul_cska32_fa3_24_or0[0]), .fa_xor1(u_csamul_cska32_fa3_25_xor1), .fa_or0(u_csamul_cska32_fa3_25_or0));
  and_gate and_gate_u_csamul_cska32_and4_25(.a(a[4]), .b(b[25]), .out(u_csamul_cska32_and4_25));
  fa fa_u_csamul_cska32_fa4_25_out(.a(u_csamul_cska32_and4_25[0]), .b(u_csamul_cska32_fa5_24_xor1[0]), .cin(u_csamul_cska32_fa4_24_or0[0]), .fa_xor1(u_csamul_cska32_fa4_25_xor1), .fa_or0(u_csamul_cska32_fa4_25_or0));
  and_gate and_gate_u_csamul_cska32_and5_25(.a(a[5]), .b(b[25]), .out(u_csamul_cska32_and5_25));
  fa fa_u_csamul_cska32_fa5_25_out(.a(u_csamul_cska32_and5_25[0]), .b(u_csamul_cska32_fa6_24_xor1[0]), .cin(u_csamul_cska32_fa5_24_or0[0]), .fa_xor1(u_csamul_cska32_fa5_25_xor1), .fa_or0(u_csamul_cska32_fa5_25_or0));
  and_gate and_gate_u_csamul_cska32_and6_25(.a(a[6]), .b(b[25]), .out(u_csamul_cska32_and6_25));
  fa fa_u_csamul_cska32_fa6_25_out(.a(u_csamul_cska32_and6_25[0]), .b(u_csamul_cska32_fa7_24_xor1[0]), .cin(u_csamul_cska32_fa6_24_or0[0]), .fa_xor1(u_csamul_cska32_fa6_25_xor1), .fa_or0(u_csamul_cska32_fa6_25_or0));
  and_gate and_gate_u_csamul_cska32_and7_25(.a(a[7]), .b(b[25]), .out(u_csamul_cska32_and7_25));
  fa fa_u_csamul_cska32_fa7_25_out(.a(u_csamul_cska32_and7_25[0]), .b(u_csamul_cska32_fa8_24_xor1[0]), .cin(u_csamul_cska32_fa7_24_or0[0]), .fa_xor1(u_csamul_cska32_fa7_25_xor1), .fa_or0(u_csamul_cska32_fa7_25_or0));
  and_gate and_gate_u_csamul_cska32_and8_25(.a(a[8]), .b(b[25]), .out(u_csamul_cska32_and8_25));
  fa fa_u_csamul_cska32_fa8_25_out(.a(u_csamul_cska32_and8_25[0]), .b(u_csamul_cska32_fa9_24_xor1[0]), .cin(u_csamul_cska32_fa8_24_or0[0]), .fa_xor1(u_csamul_cska32_fa8_25_xor1), .fa_or0(u_csamul_cska32_fa8_25_or0));
  and_gate and_gate_u_csamul_cska32_and9_25(.a(a[9]), .b(b[25]), .out(u_csamul_cska32_and9_25));
  fa fa_u_csamul_cska32_fa9_25_out(.a(u_csamul_cska32_and9_25[0]), .b(u_csamul_cska32_fa10_24_xor1[0]), .cin(u_csamul_cska32_fa9_24_or0[0]), .fa_xor1(u_csamul_cska32_fa9_25_xor1), .fa_or0(u_csamul_cska32_fa9_25_or0));
  and_gate and_gate_u_csamul_cska32_and10_25(.a(a[10]), .b(b[25]), .out(u_csamul_cska32_and10_25));
  fa fa_u_csamul_cska32_fa10_25_out(.a(u_csamul_cska32_and10_25[0]), .b(u_csamul_cska32_fa11_24_xor1[0]), .cin(u_csamul_cska32_fa10_24_or0[0]), .fa_xor1(u_csamul_cska32_fa10_25_xor1), .fa_or0(u_csamul_cska32_fa10_25_or0));
  and_gate and_gate_u_csamul_cska32_and11_25(.a(a[11]), .b(b[25]), .out(u_csamul_cska32_and11_25));
  fa fa_u_csamul_cska32_fa11_25_out(.a(u_csamul_cska32_and11_25[0]), .b(u_csamul_cska32_fa12_24_xor1[0]), .cin(u_csamul_cska32_fa11_24_or0[0]), .fa_xor1(u_csamul_cska32_fa11_25_xor1), .fa_or0(u_csamul_cska32_fa11_25_or0));
  and_gate and_gate_u_csamul_cska32_and12_25(.a(a[12]), .b(b[25]), .out(u_csamul_cska32_and12_25));
  fa fa_u_csamul_cska32_fa12_25_out(.a(u_csamul_cska32_and12_25[0]), .b(u_csamul_cska32_fa13_24_xor1[0]), .cin(u_csamul_cska32_fa12_24_or0[0]), .fa_xor1(u_csamul_cska32_fa12_25_xor1), .fa_or0(u_csamul_cska32_fa12_25_or0));
  and_gate and_gate_u_csamul_cska32_and13_25(.a(a[13]), .b(b[25]), .out(u_csamul_cska32_and13_25));
  fa fa_u_csamul_cska32_fa13_25_out(.a(u_csamul_cska32_and13_25[0]), .b(u_csamul_cska32_fa14_24_xor1[0]), .cin(u_csamul_cska32_fa13_24_or0[0]), .fa_xor1(u_csamul_cska32_fa13_25_xor1), .fa_or0(u_csamul_cska32_fa13_25_or0));
  and_gate and_gate_u_csamul_cska32_and14_25(.a(a[14]), .b(b[25]), .out(u_csamul_cska32_and14_25));
  fa fa_u_csamul_cska32_fa14_25_out(.a(u_csamul_cska32_and14_25[0]), .b(u_csamul_cska32_fa15_24_xor1[0]), .cin(u_csamul_cska32_fa14_24_or0[0]), .fa_xor1(u_csamul_cska32_fa14_25_xor1), .fa_or0(u_csamul_cska32_fa14_25_or0));
  and_gate and_gate_u_csamul_cska32_and15_25(.a(a[15]), .b(b[25]), .out(u_csamul_cska32_and15_25));
  fa fa_u_csamul_cska32_fa15_25_out(.a(u_csamul_cska32_and15_25[0]), .b(u_csamul_cska32_fa16_24_xor1[0]), .cin(u_csamul_cska32_fa15_24_or0[0]), .fa_xor1(u_csamul_cska32_fa15_25_xor1), .fa_or0(u_csamul_cska32_fa15_25_or0));
  and_gate and_gate_u_csamul_cska32_and16_25(.a(a[16]), .b(b[25]), .out(u_csamul_cska32_and16_25));
  fa fa_u_csamul_cska32_fa16_25_out(.a(u_csamul_cska32_and16_25[0]), .b(u_csamul_cska32_fa17_24_xor1[0]), .cin(u_csamul_cska32_fa16_24_or0[0]), .fa_xor1(u_csamul_cska32_fa16_25_xor1), .fa_or0(u_csamul_cska32_fa16_25_or0));
  and_gate and_gate_u_csamul_cska32_and17_25(.a(a[17]), .b(b[25]), .out(u_csamul_cska32_and17_25));
  fa fa_u_csamul_cska32_fa17_25_out(.a(u_csamul_cska32_and17_25[0]), .b(u_csamul_cska32_fa18_24_xor1[0]), .cin(u_csamul_cska32_fa17_24_or0[0]), .fa_xor1(u_csamul_cska32_fa17_25_xor1), .fa_or0(u_csamul_cska32_fa17_25_or0));
  and_gate and_gate_u_csamul_cska32_and18_25(.a(a[18]), .b(b[25]), .out(u_csamul_cska32_and18_25));
  fa fa_u_csamul_cska32_fa18_25_out(.a(u_csamul_cska32_and18_25[0]), .b(u_csamul_cska32_fa19_24_xor1[0]), .cin(u_csamul_cska32_fa18_24_or0[0]), .fa_xor1(u_csamul_cska32_fa18_25_xor1), .fa_or0(u_csamul_cska32_fa18_25_or0));
  and_gate and_gate_u_csamul_cska32_and19_25(.a(a[19]), .b(b[25]), .out(u_csamul_cska32_and19_25));
  fa fa_u_csamul_cska32_fa19_25_out(.a(u_csamul_cska32_and19_25[0]), .b(u_csamul_cska32_fa20_24_xor1[0]), .cin(u_csamul_cska32_fa19_24_or0[0]), .fa_xor1(u_csamul_cska32_fa19_25_xor1), .fa_or0(u_csamul_cska32_fa19_25_or0));
  and_gate and_gate_u_csamul_cska32_and20_25(.a(a[20]), .b(b[25]), .out(u_csamul_cska32_and20_25));
  fa fa_u_csamul_cska32_fa20_25_out(.a(u_csamul_cska32_and20_25[0]), .b(u_csamul_cska32_fa21_24_xor1[0]), .cin(u_csamul_cska32_fa20_24_or0[0]), .fa_xor1(u_csamul_cska32_fa20_25_xor1), .fa_or0(u_csamul_cska32_fa20_25_or0));
  and_gate and_gate_u_csamul_cska32_and21_25(.a(a[21]), .b(b[25]), .out(u_csamul_cska32_and21_25));
  fa fa_u_csamul_cska32_fa21_25_out(.a(u_csamul_cska32_and21_25[0]), .b(u_csamul_cska32_fa22_24_xor1[0]), .cin(u_csamul_cska32_fa21_24_or0[0]), .fa_xor1(u_csamul_cska32_fa21_25_xor1), .fa_or0(u_csamul_cska32_fa21_25_or0));
  and_gate and_gate_u_csamul_cska32_and22_25(.a(a[22]), .b(b[25]), .out(u_csamul_cska32_and22_25));
  fa fa_u_csamul_cska32_fa22_25_out(.a(u_csamul_cska32_and22_25[0]), .b(u_csamul_cska32_fa23_24_xor1[0]), .cin(u_csamul_cska32_fa22_24_or0[0]), .fa_xor1(u_csamul_cska32_fa22_25_xor1), .fa_or0(u_csamul_cska32_fa22_25_or0));
  and_gate and_gate_u_csamul_cska32_and23_25(.a(a[23]), .b(b[25]), .out(u_csamul_cska32_and23_25));
  fa fa_u_csamul_cska32_fa23_25_out(.a(u_csamul_cska32_and23_25[0]), .b(u_csamul_cska32_fa24_24_xor1[0]), .cin(u_csamul_cska32_fa23_24_or0[0]), .fa_xor1(u_csamul_cska32_fa23_25_xor1), .fa_or0(u_csamul_cska32_fa23_25_or0));
  and_gate and_gate_u_csamul_cska32_and24_25(.a(a[24]), .b(b[25]), .out(u_csamul_cska32_and24_25));
  fa fa_u_csamul_cska32_fa24_25_out(.a(u_csamul_cska32_and24_25[0]), .b(u_csamul_cska32_fa25_24_xor1[0]), .cin(u_csamul_cska32_fa24_24_or0[0]), .fa_xor1(u_csamul_cska32_fa24_25_xor1), .fa_or0(u_csamul_cska32_fa24_25_or0));
  and_gate and_gate_u_csamul_cska32_and25_25(.a(a[25]), .b(b[25]), .out(u_csamul_cska32_and25_25));
  fa fa_u_csamul_cska32_fa25_25_out(.a(u_csamul_cska32_and25_25[0]), .b(u_csamul_cska32_fa26_24_xor1[0]), .cin(u_csamul_cska32_fa25_24_or0[0]), .fa_xor1(u_csamul_cska32_fa25_25_xor1), .fa_or0(u_csamul_cska32_fa25_25_or0));
  and_gate and_gate_u_csamul_cska32_and26_25(.a(a[26]), .b(b[25]), .out(u_csamul_cska32_and26_25));
  fa fa_u_csamul_cska32_fa26_25_out(.a(u_csamul_cska32_and26_25[0]), .b(u_csamul_cska32_fa27_24_xor1[0]), .cin(u_csamul_cska32_fa26_24_or0[0]), .fa_xor1(u_csamul_cska32_fa26_25_xor1), .fa_or0(u_csamul_cska32_fa26_25_or0));
  and_gate and_gate_u_csamul_cska32_and27_25(.a(a[27]), .b(b[25]), .out(u_csamul_cska32_and27_25));
  fa fa_u_csamul_cska32_fa27_25_out(.a(u_csamul_cska32_and27_25[0]), .b(u_csamul_cska32_fa28_24_xor1[0]), .cin(u_csamul_cska32_fa27_24_or0[0]), .fa_xor1(u_csamul_cska32_fa27_25_xor1), .fa_or0(u_csamul_cska32_fa27_25_or0));
  and_gate and_gate_u_csamul_cska32_and28_25(.a(a[28]), .b(b[25]), .out(u_csamul_cska32_and28_25));
  fa fa_u_csamul_cska32_fa28_25_out(.a(u_csamul_cska32_and28_25[0]), .b(u_csamul_cska32_fa29_24_xor1[0]), .cin(u_csamul_cska32_fa28_24_or0[0]), .fa_xor1(u_csamul_cska32_fa28_25_xor1), .fa_or0(u_csamul_cska32_fa28_25_or0));
  and_gate and_gate_u_csamul_cska32_and29_25(.a(a[29]), .b(b[25]), .out(u_csamul_cska32_and29_25));
  fa fa_u_csamul_cska32_fa29_25_out(.a(u_csamul_cska32_and29_25[0]), .b(u_csamul_cska32_fa30_24_xor1[0]), .cin(u_csamul_cska32_fa29_24_or0[0]), .fa_xor1(u_csamul_cska32_fa29_25_xor1), .fa_or0(u_csamul_cska32_fa29_25_or0));
  and_gate and_gate_u_csamul_cska32_and30_25(.a(a[30]), .b(b[25]), .out(u_csamul_cska32_and30_25));
  fa fa_u_csamul_cska32_fa30_25_out(.a(u_csamul_cska32_and30_25[0]), .b(u_csamul_cska32_and31_24[0]), .cin(u_csamul_cska32_fa30_24_or0[0]), .fa_xor1(u_csamul_cska32_fa30_25_xor1), .fa_or0(u_csamul_cska32_fa30_25_or0));
  and_gate and_gate_u_csamul_cska32_and31_25(.a(a[31]), .b(b[25]), .out(u_csamul_cska32_and31_25));
  and_gate and_gate_u_csamul_cska32_and0_26(.a(a[0]), .b(b[26]), .out(u_csamul_cska32_and0_26));
  fa fa_u_csamul_cska32_fa0_26_out(.a(u_csamul_cska32_and0_26[0]), .b(u_csamul_cska32_fa1_25_xor1[0]), .cin(u_csamul_cska32_fa0_25_or0[0]), .fa_xor1(u_csamul_cska32_fa0_26_xor1), .fa_or0(u_csamul_cska32_fa0_26_or0));
  and_gate and_gate_u_csamul_cska32_and1_26(.a(a[1]), .b(b[26]), .out(u_csamul_cska32_and1_26));
  fa fa_u_csamul_cska32_fa1_26_out(.a(u_csamul_cska32_and1_26[0]), .b(u_csamul_cska32_fa2_25_xor1[0]), .cin(u_csamul_cska32_fa1_25_or0[0]), .fa_xor1(u_csamul_cska32_fa1_26_xor1), .fa_or0(u_csamul_cska32_fa1_26_or0));
  and_gate and_gate_u_csamul_cska32_and2_26(.a(a[2]), .b(b[26]), .out(u_csamul_cska32_and2_26));
  fa fa_u_csamul_cska32_fa2_26_out(.a(u_csamul_cska32_and2_26[0]), .b(u_csamul_cska32_fa3_25_xor1[0]), .cin(u_csamul_cska32_fa2_25_or0[0]), .fa_xor1(u_csamul_cska32_fa2_26_xor1), .fa_or0(u_csamul_cska32_fa2_26_or0));
  and_gate and_gate_u_csamul_cska32_and3_26(.a(a[3]), .b(b[26]), .out(u_csamul_cska32_and3_26));
  fa fa_u_csamul_cska32_fa3_26_out(.a(u_csamul_cska32_and3_26[0]), .b(u_csamul_cska32_fa4_25_xor1[0]), .cin(u_csamul_cska32_fa3_25_or0[0]), .fa_xor1(u_csamul_cska32_fa3_26_xor1), .fa_or0(u_csamul_cska32_fa3_26_or0));
  and_gate and_gate_u_csamul_cska32_and4_26(.a(a[4]), .b(b[26]), .out(u_csamul_cska32_and4_26));
  fa fa_u_csamul_cska32_fa4_26_out(.a(u_csamul_cska32_and4_26[0]), .b(u_csamul_cska32_fa5_25_xor1[0]), .cin(u_csamul_cska32_fa4_25_or0[0]), .fa_xor1(u_csamul_cska32_fa4_26_xor1), .fa_or0(u_csamul_cska32_fa4_26_or0));
  and_gate and_gate_u_csamul_cska32_and5_26(.a(a[5]), .b(b[26]), .out(u_csamul_cska32_and5_26));
  fa fa_u_csamul_cska32_fa5_26_out(.a(u_csamul_cska32_and5_26[0]), .b(u_csamul_cska32_fa6_25_xor1[0]), .cin(u_csamul_cska32_fa5_25_or0[0]), .fa_xor1(u_csamul_cska32_fa5_26_xor1), .fa_or0(u_csamul_cska32_fa5_26_or0));
  and_gate and_gate_u_csamul_cska32_and6_26(.a(a[6]), .b(b[26]), .out(u_csamul_cska32_and6_26));
  fa fa_u_csamul_cska32_fa6_26_out(.a(u_csamul_cska32_and6_26[0]), .b(u_csamul_cska32_fa7_25_xor1[0]), .cin(u_csamul_cska32_fa6_25_or0[0]), .fa_xor1(u_csamul_cska32_fa6_26_xor1), .fa_or0(u_csamul_cska32_fa6_26_or0));
  and_gate and_gate_u_csamul_cska32_and7_26(.a(a[7]), .b(b[26]), .out(u_csamul_cska32_and7_26));
  fa fa_u_csamul_cska32_fa7_26_out(.a(u_csamul_cska32_and7_26[0]), .b(u_csamul_cska32_fa8_25_xor1[0]), .cin(u_csamul_cska32_fa7_25_or0[0]), .fa_xor1(u_csamul_cska32_fa7_26_xor1), .fa_or0(u_csamul_cska32_fa7_26_or0));
  and_gate and_gate_u_csamul_cska32_and8_26(.a(a[8]), .b(b[26]), .out(u_csamul_cska32_and8_26));
  fa fa_u_csamul_cska32_fa8_26_out(.a(u_csamul_cska32_and8_26[0]), .b(u_csamul_cska32_fa9_25_xor1[0]), .cin(u_csamul_cska32_fa8_25_or0[0]), .fa_xor1(u_csamul_cska32_fa8_26_xor1), .fa_or0(u_csamul_cska32_fa8_26_or0));
  and_gate and_gate_u_csamul_cska32_and9_26(.a(a[9]), .b(b[26]), .out(u_csamul_cska32_and9_26));
  fa fa_u_csamul_cska32_fa9_26_out(.a(u_csamul_cska32_and9_26[0]), .b(u_csamul_cska32_fa10_25_xor1[0]), .cin(u_csamul_cska32_fa9_25_or0[0]), .fa_xor1(u_csamul_cska32_fa9_26_xor1), .fa_or0(u_csamul_cska32_fa9_26_or0));
  and_gate and_gate_u_csamul_cska32_and10_26(.a(a[10]), .b(b[26]), .out(u_csamul_cska32_and10_26));
  fa fa_u_csamul_cska32_fa10_26_out(.a(u_csamul_cska32_and10_26[0]), .b(u_csamul_cska32_fa11_25_xor1[0]), .cin(u_csamul_cska32_fa10_25_or0[0]), .fa_xor1(u_csamul_cska32_fa10_26_xor1), .fa_or0(u_csamul_cska32_fa10_26_or0));
  and_gate and_gate_u_csamul_cska32_and11_26(.a(a[11]), .b(b[26]), .out(u_csamul_cska32_and11_26));
  fa fa_u_csamul_cska32_fa11_26_out(.a(u_csamul_cska32_and11_26[0]), .b(u_csamul_cska32_fa12_25_xor1[0]), .cin(u_csamul_cska32_fa11_25_or0[0]), .fa_xor1(u_csamul_cska32_fa11_26_xor1), .fa_or0(u_csamul_cska32_fa11_26_or0));
  and_gate and_gate_u_csamul_cska32_and12_26(.a(a[12]), .b(b[26]), .out(u_csamul_cska32_and12_26));
  fa fa_u_csamul_cska32_fa12_26_out(.a(u_csamul_cska32_and12_26[0]), .b(u_csamul_cska32_fa13_25_xor1[0]), .cin(u_csamul_cska32_fa12_25_or0[0]), .fa_xor1(u_csamul_cska32_fa12_26_xor1), .fa_or0(u_csamul_cska32_fa12_26_or0));
  and_gate and_gate_u_csamul_cska32_and13_26(.a(a[13]), .b(b[26]), .out(u_csamul_cska32_and13_26));
  fa fa_u_csamul_cska32_fa13_26_out(.a(u_csamul_cska32_and13_26[0]), .b(u_csamul_cska32_fa14_25_xor1[0]), .cin(u_csamul_cska32_fa13_25_or0[0]), .fa_xor1(u_csamul_cska32_fa13_26_xor1), .fa_or0(u_csamul_cska32_fa13_26_or0));
  and_gate and_gate_u_csamul_cska32_and14_26(.a(a[14]), .b(b[26]), .out(u_csamul_cska32_and14_26));
  fa fa_u_csamul_cska32_fa14_26_out(.a(u_csamul_cska32_and14_26[0]), .b(u_csamul_cska32_fa15_25_xor1[0]), .cin(u_csamul_cska32_fa14_25_or0[0]), .fa_xor1(u_csamul_cska32_fa14_26_xor1), .fa_or0(u_csamul_cska32_fa14_26_or0));
  and_gate and_gate_u_csamul_cska32_and15_26(.a(a[15]), .b(b[26]), .out(u_csamul_cska32_and15_26));
  fa fa_u_csamul_cska32_fa15_26_out(.a(u_csamul_cska32_and15_26[0]), .b(u_csamul_cska32_fa16_25_xor1[0]), .cin(u_csamul_cska32_fa15_25_or0[0]), .fa_xor1(u_csamul_cska32_fa15_26_xor1), .fa_or0(u_csamul_cska32_fa15_26_or0));
  and_gate and_gate_u_csamul_cska32_and16_26(.a(a[16]), .b(b[26]), .out(u_csamul_cska32_and16_26));
  fa fa_u_csamul_cska32_fa16_26_out(.a(u_csamul_cska32_and16_26[0]), .b(u_csamul_cska32_fa17_25_xor1[0]), .cin(u_csamul_cska32_fa16_25_or0[0]), .fa_xor1(u_csamul_cska32_fa16_26_xor1), .fa_or0(u_csamul_cska32_fa16_26_or0));
  and_gate and_gate_u_csamul_cska32_and17_26(.a(a[17]), .b(b[26]), .out(u_csamul_cska32_and17_26));
  fa fa_u_csamul_cska32_fa17_26_out(.a(u_csamul_cska32_and17_26[0]), .b(u_csamul_cska32_fa18_25_xor1[0]), .cin(u_csamul_cska32_fa17_25_or0[0]), .fa_xor1(u_csamul_cska32_fa17_26_xor1), .fa_or0(u_csamul_cska32_fa17_26_or0));
  and_gate and_gate_u_csamul_cska32_and18_26(.a(a[18]), .b(b[26]), .out(u_csamul_cska32_and18_26));
  fa fa_u_csamul_cska32_fa18_26_out(.a(u_csamul_cska32_and18_26[0]), .b(u_csamul_cska32_fa19_25_xor1[0]), .cin(u_csamul_cska32_fa18_25_or0[0]), .fa_xor1(u_csamul_cska32_fa18_26_xor1), .fa_or0(u_csamul_cska32_fa18_26_or0));
  and_gate and_gate_u_csamul_cska32_and19_26(.a(a[19]), .b(b[26]), .out(u_csamul_cska32_and19_26));
  fa fa_u_csamul_cska32_fa19_26_out(.a(u_csamul_cska32_and19_26[0]), .b(u_csamul_cska32_fa20_25_xor1[0]), .cin(u_csamul_cska32_fa19_25_or0[0]), .fa_xor1(u_csamul_cska32_fa19_26_xor1), .fa_or0(u_csamul_cska32_fa19_26_or0));
  and_gate and_gate_u_csamul_cska32_and20_26(.a(a[20]), .b(b[26]), .out(u_csamul_cska32_and20_26));
  fa fa_u_csamul_cska32_fa20_26_out(.a(u_csamul_cska32_and20_26[0]), .b(u_csamul_cska32_fa21_25_xor1[0]), .cin(u_csamul_cska32_fa20_25_or0[0]), .fa_xor1(u_csamul_cska32_fa20_26_xor1), .fa_or0(u_csamul_cska32_fa20_26_or0));
  and_gate and_gate_u_csamul_cska32_and21_26(.a(a[21]), .b(b[26]), .out(u_csamul_cska32_and21_26));
  fa fa_u_csamul_cska32_fa21_26_out(.a(u_csamul_cska32_and21_26[0]), .b(u_csamul_cska32_fa22_25_xor1[0]), .cin(u_csamul_cska32_fa21_25_or0[0]), .fa_xor1(u_csamul_cska32_fa21_26_xor1), .fa_or0(u_csamul_cska32_fa21_26_or0));
  and_gate and_gate_u_csamul_cska32_and22_26(.a(a[22]), .b(b[26]), .out(u_csamul_cska32_and22_26));
  fa fa_u_csamul_cska32_fa22_26_out(.a(u_csamul_cska32_and22_26[0]), .b(u_csamul_cska32_fa23_25_xor1[0]), .cin(u_csamul_cska32_fa22_25_or0[0]), .fa_xor1(u_csamul_cska32_fa22_26_xor1), .fa_or0(u_csamul_cska32_fa22_26_or0));
  and_gate and_gate_u_csamul_cska32_and23_26(.a(a[23]), .b(b[26]), .out(u_csamul_cska32_and23_26));
  fa fa_u_csamul_cska32_fa23_26_out(.a(u_csamul_cska32_and23_26[0]), .b(u_csamul_cska32_fa24_25_xor1[0]), .cin(u_csamul_cska32_fa23_25_or0[0]), .fa_xor1(u_csamul_cska32_fa23_26_xor1), .fa_or0(u_csamul_cska32_fa23_26_or0));
  and_gate and_gate_u_csamul_cska32_and24_26(.a(a[24]), .b(b[26]), .out(u_csamul_cska32_and24_26));
  fa fa_u_csamul_cska32_fa24_26_out(.a(u_csamul_cska32_and24_26[0]), .b(u_csamul_cska32_fa25_25_xor1[0]), .cin(u_csamul_cska32_fa24_25_or0[0]), .fa_xor1(u_csamul_cska32_fa24_26_xor1), .fa_or0(u_csamul_cska32_fa24_26_or0));
  and_gate and_gate_u_csamul_cska32_and25_26(.a(a[25]), .b(b[26]), .out(u_csamul_cska32_and25_26));
  fa fa_u_csamul_cska32_fa25_26_out(.a(u_csamul_cska32_and25_26[0]), .b(u_csamul_cska32_fa26_25_xor1[0]), .cin(u_csamul_cska32_fa25_25_or0[0]), .fa_xor1(u_csamul_cska32_fa25_26_xor1), .fa_or0(u_csamul_cska32_fa25_26_or0));
  and_gate and_gate_u_csamul_cska32_and26_26(.a(a[26]), .b(b[26]), .out(u_csamul_cska32_and26_26));
  fa fa_u_csamul_cska32_fa26_26_out(.a(u_csamul_cska32_and26_26[0]), .b(u_csamul_cska32_fa27_25_xor1[0]), .cin(u_csamul_cska32_fa26_25_or0[0]), .fa_xor1(u_csamul_cska32_fa26_26_xor1), .fa_or0(u_csamul_cska32_fa26_26_or0));
  and_gate and_gate_u_csamul_cska32_and27_26(.a(a[27]), .b(b[26]), .out(u_csamul_cska32_and27_26));
  fa fa_u_csamul_cska32_fa27_26_out(.a(u_csamul_cska32_and27_26[0]), .b(u_csamul_cska32_fa28_25_xor1[0]), .cin(u_csamul_cska32_fa27_25_or0[0]), .fa_xor1(u_csamul_cska32_fa27_26_xor1), .fa_or0(u_csamul_cska32_fa27_26_or0));
  and_gate and_gate_u_csamul_cska32_and28_26(.a(a[28]), .b(b[26]), .out(u_csamul_cska32_and28_26));
  fa fa_u_csamul_cska32_fa28_26_out(.a(u_csamul_cska32_and28_26[0]), .b(u_csamul_cska32_fa29_25_xor1[0]), .cin(u_csamul_cska32_fa28_25_or0[0]), .fa_xor1(u_csamul_cska32_fa28_26_xor1), .fa_or0(u_csamul_cska32_fa28_26_or0));
  and_gate and_gate_u_csamul_cska32_and29_26(.a(a[29]), .b(b[26]), .out(u_csamul_cska32_and29_26));
  fa fa_u_csamul_cska32_fa29_26_out(.a(u_csamul_cska32_and29_26[0]), .b(u_csamul_cska32_fa30_25_xor1[0]), .cin(u_csamul_cska32_fa29_25_or0[0]), .fa_xor1(u_csamul_cska32_fa29_26_xor1), .fa_or0(u_csamul_cska32_fa29_26_or0));
  and_gate and_gate_u_csamul_cska32_and30_26(.a(a[30]), .b(b[26]), .out(u_csamul_cska32_and30_26));
  fa fa_u_csamul_cska32_fa30_26_out(.a(u_csamul_cska32_and30_26[0]), .b(u_csamul_cska32_and31_25[0]), .cin(u_csamul_cska32_fa30_25_or0[0]), .fa_xor1(u_csamul_cska32_fa30_26_xor1), .fa_or0(u_csamul_cska32_fa30_26_or0));
  and_gate and_gate_u_csamul_cska32_and31_26(.a(a[31]), .b(b[26]), .out(u_csamul_cska32_and31_26));
  and_gate and_gate_u_csamul_cska32_and0_27(.a(a[0]), .b(b[27]), .out(u_csamul_cska32_and0_27));
  fa fa_u_csamul_cska32_fa0_27_out(.a(u_csamul_cska32_and0_27[0]), .b(u_csamul_cska32_fa1_26_xor1[0]), .cin(u_csamul_cska32_fa0_26_or0[0]), .fa_xor1(u_csamul_cska32_fa0_27_xor1), .fa_or0(u_csamul_cska32_fa0_27_or0));
  and_gate and_gate_u_csamul_cska32_and1_27(.a(a[1]), .b(b[27]), .out(u_csamul_cska32_and1_27));
  fa fa_u_csamul_cska32_fa1_27_out(.a(u_csamul_cska32_and1_27[0]), .b(u_csamul_cska32_fa2_26_xor1[0]), .cin(u_csamul_cska32_fa1_26_or0[0]), .fa_xor1(u_csamul_cska32_fa1_27_xor1), .fa_or0(u_csamul_cska32_fa1_27_or0));
  and_gate and_gate_u_csamul_cska32_and2_27(.a(a[2]), .b(b[27]), .out(u_csamul_cska32_and2_27));
  fa fa_u_csamul_cska32_fa2_27_out(.a(u_csamul_cska32_and2_27[0]), .b(u_csamul_cska32_fa3_26_xor1[0]), .cin(u_csamul_cska32_fa2_26_or0[0]), .fa_xor1(u_csamul_cska32_fa2_27_xor1), .fa_or0(u_csamul_cska32_fa2_27_or0));
  and_gate and_gate_u_csamul_cska32_and3_27(.a(a[3]), .b(b[27]), .out(u_csamul_cska32_and3_27));
  fa fa_u_csamul_cska32_fa3_27_out(.a(u_csamul_cska32_and3_27[0]), .b(u_csamul_cska32_fa4_26_xor1[0]), .cin(u_csamul_cska32_fa3_26_or0[0]), .fa_xor1(u_csamul_cska32_fa3_27_xor1), .fa_or0(u_csamul_cska32_fa3_27_or0));
  and_gate and_gate_u_csamul_cska32_and4_27(.a(a[4]), .b(b[27]), .out(u_csamul_cska32_and4_27));
  fa fa_u_csamul_cska32_fa4_27_out(.a(u_csamul_cska32_and4_27[0]), .b(u_csamul_cska32_fa5_26_xor1[0]), .cin(u_csamul_cska32_fa4_26_or0[0]), .fa_xor1(u_csamul_cska32_fa4_27_xor1), .fa_or0(u_csamul_cska32_fa4_27_or0));
  and_gate and_gate_u_csamul_cska32_and5_27(.a(a[5]), .b(b[27]), .out(u_csamul_cska32_and5_27));
  fa fa_u_csamul_cska32_fa5_27_out(.a(u_csamul_cska32_and5_27[0]), .b(u_csamul_cska32_fa6_26_xor1[0]), .cin(u_csamul_cska32_fa5_26_or0[0]), .fa_xor1(u_csamul_cska32_fa5_27_xor1), .fa_or0(u_csamul_cska32_fa5_27_or0));
  and_gate and_gate_u_csamul_cska32_and6_27(.a(a[6]), .b(b[27]), .out(u_csamul_cska32_and6_27));
  fa fa_u_csamul_cska32_fa6_27_out(.a(u_csamul_cska32_and6_27[0]), .b(u_csamul_cska32_fa7_26_xor1[0]), .cin(u_csamul_cska32_fa6_26_or0[0]), .fa_xor1(u_csamul_cska32_fa6_27_xor1), .fa_or0(u_csamul_cska32_fa6_27_or0));
  and_gate and_gate_u_csamul_cska32_and7_27(.a(a[7]), .b(b[27]), .out(u_csamul_cska32_and7_27));
  fa fa_u_csamul_cska32_fa7_27_out(.a(u_csamul_cska32_and7_27[0]), .b(u_csamul_cska32_fa8_26_xor1[0]), .cin(u_csamul_cska32_fa7_26_or0[0]), .fa_xor1(u_csamul_cska32_fa7_27_xor1), .fa_or0(u_csamul_cska32_fa7_27_or0));
  and_gate and_gate_u_csamul_cska32_and8_27(.a(a[8]), .b(b[27]), .out(u_csamul_cska32_and8_27));
  fa fa_u_csamul_cska32_fa8_27_out(.a(u_csamul_cska32_and8_27[0]), .b(u_csamul_cska32_fa9_26_xor1[0]), .cin(u_csamul_cska32_fa8_26_or0[0]), .fa_xor1(u_csamul_cska32_fa8_27_xor1), .fa_or0(u_csamul_cska32_fa8_27_or0));
  and_gate and_gate_u_csamul_cska32_and9_27(.a(a[9]), .b(b[27]), .out(u_csamul_cska32_and9_27));
  fa fa_u_csamul_cska32_fa9_27_out(.a(u_csamul_cska32_and9_27[0]), .b(u_csamul_cska32_fa10_26_xor1[0]), .cin(u_csamul_cska32_fa9_26_or0[0]), .fa_xor1(u_csamul_cska32_fa9_27_xor1), .fa_or0(u_csamul_cska32_fa9_27_or0));
  and_gate and_gate_u_csamul_cska32_and10_27(.a(a[10]), .b(b[27]), .out(u_csamul_cska32_and10_27));
  fa fa_u_csamul_cska32_fa10_27_out(.a(u_csamul_cska32_and10_27[0]), .b(u_csamul_cska32_fa11_26_xor1[0]), .cin(u_csamul_cska32_fa10_26_or0[0]), .fa_xor1(u_csamul_cska32_fa10_27_xor1), .fa_or0(u_csamul_cska32_fa10_27_or0));
  and_gate and_gate_u_csamul_cska32_and11_27(.a(a[11]), .b(b[27]), .out(u_csamul_cska32_and11_27));
  fa fa_u_csamul_cska32_fa11_27_out(.a(u_csamul_cska32_and11_27[0]), .b(u_csamul_cska32_fa12_26_xor1[0]), .cin(u_csamul_cska32_fa11_26_or0[0]), .fa_xor1(u_csamul_cska32_fa11_27_xor1), .fa_or0(u_csamul_cska32_fa11_27_or0));
  and_gate and_gate_u_csamul_cska32_and12_27(.a(a[12]), .b(b[27]), .out(u_csamul_cska32_and12_27));
  fa fa_u_csamul_cska32_fa12_27_out(.a(u_csamul_cska32_and12_27[0]), .b(u_csamul_cska32_fa13_26_xor1[0]), .cin(u_csamul_cska32_fa12_26_or0[0]), .fa_xor1(u_csamul_cska32_fa12_27_xor1), .fa_or0(u_csamul_cska32_fa12_27_or0));
  and_gate and_gate_u_csamul_cska32_and13_27(.a(a[13]), .b(b[27]), .out(u_csamul_cska32_and13_27));
  fa fa_u_csamul_cska32_fa13_27_out(.a(u_csamul_cska32_and13_27[0]), .b(u_csamul_cska32_fa14_26_xor1[0]), .cin(u_csamul_cska32_fa13_26_or0[0]), .fa_xor1(u_csamul_cska32_fa13_27_xor1), .fa_or0(u_csamul_cska32_fa13_27_or0));
  and_gate and_gate_u_csamul_cska32_and14_27(.a(a[14]), .b(b[27]), .out(u_csamul_cska32_and14_27));
  fa fa_u_csamul_cska32_fa14_27_out(.a(u_csamul_cska32_and14_27[0]), .b(u_csamul_cska32_fa15_26_xor1[0]), .cin(u_csamul_cska32_fa14_26_or0[0]), .fa_xor1(u_csamul_cska32_fa14_27_xor1), .fa_or0(u_csamul_cska32_fa14_27_or0));
  and_gate and_gate_u_csamul_cska32_and15_27(.a(a[15]), .b(b[27]), .out(u_csamul_cska32_and15_27));
  fa fa_u_csamul_cska32_fa15_27_out(.a(u_csamul_cska32_and15_27[0]), .b(u_csamul_cska32_fa16_26_xor1[0]), .cin(u_csamul_cska32_fa15_26_or0[0]), .fa_xor1(u_csamul_cska32_fa15_27_xor1), .fa_or0(u_csamul_cska32_fa15_27_or0));
  and_gate and_gate_u_csamul_cska32_and16_27(.a(a[16]), .b(b[27]), .out(u_csamul_cska32_and16_27));
  fa fa_u_csamul_cska32_fa16_27_out(.a(u_csamul_cska32_and16_27[0]), .b(u_csamul_cska32_fa17_26_xor1[0]), .cin(u_csamul_cska32_fa16_26_or0[0]), .fa_xor1(u_csamul_cska32_fa16_27_xor1), .fa_or0(u_csamul_cska32_fa16_27_or0));
  and_gate and_gate_u_csamul_cska32_and17_27(.a(a[17]), .b(b[27]), .out(u_csamul_cska32_and17_27));
  fa fa_u_csamul_cska32_fa17_27_out(.a(u_csamul_cska32_and17_27[0]), .b(u_csamul_cska32_fa18_26_xor1[0]), .cin(u_csamul_cska32_fa17_26_or0[0]), .fa_xor1(u_csamul_cska32_fa17_27_xor1), .fa_or0(u_csamul_cska32_fa17_27_or0));
  and_gate and_gate_u_csamul_cska32_and18_27(.a(a[18]), .b(b[27]), .out(u_csamul_cska32_and18_27));
  fa fa_u_csamul_cska32_fa18_27_out(.a(u_csamul_cska32_and18_27[0]), .b(u_csamul_cska32_fa19_26_xor1[0]), .cin(u_csamul_cska32_fa18_26_or0[0]), .fa_xor1(u_csamul_cska32_fa18_27_xor1), .fa_or0(u_csamul_cska32_fa18_27_or0));
  and_gate and_gate_u_csamul_cska32_and19_27(.a(a[19]), .b(b[27]), .out(u_csamul_cska32_and19_27));
  fa fa_u_csamul_cska32_fa19_27_out(.a(u_csamul_cska32_and19_27[0]), .b(u_csamul_cska32_fa20_26_xor1[0]), .cin(u_csamul_cska32_fa19_26_or0[0]), .fa_xor1(u_csamul_cska32_fa19_27_xor1), .fa_or0(u_csamul_cska32_fa19_27_or0));
  and_gate and_gate_u_csamul_cska32_and20_27(.a(a[20]), .b(b[27]), .out(u_csamul_cska32_and20_27));
  fa fa_u_csamul_cska32_fa20_27_out(.a(u_csamul_cska32_and20_27[0]), .b(u_csamul_cska32_fa21_26_xor1[0]), .cin(u_csamul_cska32_fa20_26_or0[0]), .fa_xor1(u_csamul_cska32_fa20_27_xor1), .fa_or0(u_csamul_cska32_fa20_27_or0));
  and_gate and_gate_u_csamul_cska32_and21_27(.a(a[21]), .b(b[27]), .out(u_csamul_cska32_and21_27));
  fa fa_u_csamul_cska32_fa21_27_out(.a(u_csamul_cska32_and21_27[0]), .b(u_csamul_cska32_fa22_26_xor1[0]), .cin(u_csamul_cska32_fa21_26_or0[0]), .fa_xor1(u_csamul_cska32_fa21_27_xor1), .fa_or0(u_csamul_cska32_fa21_27_or0));
  and_gate and_gate_u_csamul_cska32_and22_27(.a(a[22]), .b(b[27]), .out(u_csamul_cska32_and22_27));
  fa fa_u_csamul_cska32_fa22_27_out(.a(u_csamul_cska32_and22_27[0]), .b(u_csamul_cska32_fa23_26_xor1[0]), .cin(u_csamul_cska32_fa22_26_or0[0]), .fa_xor1(u_csamul_cska32_fa22_27_xor1), .fa_or0(u_csamul_cska32_fa22_27_or0));
  and_gate and_gate_u_csamul_cska32_and23_27(.a(a[23]), .b(b[27]), .out(u_csamul_cska32_and23_27));
  fa fa_u_csamul_cska32_fa23_27_out(.a(u_csamul_cska32_and23_27[0]), .b(u_csamul_cska32_fa24_26_xor1[0]), .cin(u_csamul_cska32_fa23_26_or0[0]), .fa_xor1(u_csamul_cska32_fa23_27_xor1), .fa_or0(u_csamul_cska32_fa23_27_or0));
  and_gate and_gate_u_csamul_cska32_and24_27(.a(a[24]), .b(b[27]), .out(u_csamul_cska32_and24_27));
  fa fa_u_csamul_cska32_fa24_27_out(.a(u_csamul_cska32_and24_27[0]), .b(u_csamul_cska32_fa25_26_xor1[0]), .cin(u_csamul_cska32_fa24_26_or0[0]), .fa_xor1(u_csamul_cska32_fa24_27_xor1), .fa_or0(u_csamul_cska32_fa24_27_or0));
  and_gate and_gate_u_csamul_cska32_and25_27(.a(a[25]), .b(b[27]), .out(u_csamul_cska32_and25_27));
  fa fa_u_csamul_cska32_fa25_27_out(.a(u_csamul_cska32_and25_27[0]), .b(u_csamul_cska32_fa26_26_xor1[0]), .cin(u_csamul_cska32_fa25_26_or0[0]), .fa_xor1(u_csamul_cska32_fa25_27_xor1), .fa_or0(u_csamul_cska32_fa25_27_or0));
  and_gate and_gate_u_csamul_cska32_and26_27(.a(a[26]), .b(b[27]), .out(u_csamul_cska32_and26_27));
  fa fa_u_csamul_cska32_fa26_27_out(.a(u_csamul_cska32_and26_27[0]), .b(u_csamul_cska32_fa27_26_xor1[0]), .cin(u_csamul_cska32_fa26_26_or0[0]), .fa_xor1(u_csamul_cska32_fa26_27_xor1), .fa_or0(u_csamul_cska32_fa26_27_or0));
  and_gate and_gate_u_csamul_cska32_and27_27(.a(a[27]), .b(b[27]), .out(u_csamul_cska32_and27_27));
  fa fa_u_csamul_cska32_fa27_27_out(.a(u_csamul_cska32_and27_27[0]), .b(u_csamul_cska32_fa28_26_xor1[0]), .cin(u_csamul_cska32_fa27_26_or0[0]), .fa_xor1(u_csamul_cska32_fa27_27_xor1), .fa_or0(u_csamul_cska32_fa27_27_or0));
  and_gate and_gate_u_csamul_cska32_and28_27(.a(a[28]), .b(b[27]), .out(u_csamul_cska32_and28_27));
  fa fa_u_csamul_cska32_fa28_27_out(.a(u_csamul_cska32_and28_27[0]), .b(u_csamul_cska32_fa29_26_xor1[0]), .cin(u_csamul_cska32_fa28_26_or0[0]), .fa_xor1(u_csamul_cska32_fa28_27_xor1), .fa_or0(u_csamul_cska32_fa28_27_or0));
  and_gate and_gate_u_csamul_cska32_and29_27(.a(a[29]), .b(b[27]), .out(u_csamul_cska32_and29_27));
  fa fa_u_csamul_cska32_fa29_27_out(.a(u_csamul_cska32_and29_27[0]), .b(u_csamul_cska32_fa30_26_xor1[0]), .cin(u_csamul_cska32_fa29_26_or0[0]), .fa_xor1(u_csamul_cska32_fa29_27_xor1), .fa_or0(u_csamul_cska32_fa29_27_or0));
  and_gate and_gate_u_csamul_cska32_and30_27(.a(a[30]), .b(b[27]), .out(u_csamul_cska32_and30_27));
  fa fa_u_csamul_cska32_fa30_27_out(.a(u_csamul_cska32_and30_27[0]), .b(u_csamul_cska32_and31_26[0]), .cin(u_csamul_cska32_fa30_26_or0[0]), .fa_xor1(u_csamul_cska32_fa30_27_xor1), .fa_or0(u_csamul_cska32_fa30_27_or0));
  and_gate and_gate_u_csamul_cska32_and31_27(.a(a[31]), .b(b[27]), .out(u_csamul_cska32_and31_27));
  and_gate and_gate_u_csamul_cska32_and0_28(.a(a[0]), .b(b[28]), .out(u_csamul_cska32_and0_28));
  fa fa_u_csamul_cska32_fa0_28_out(.a(u_csamul_cska32_and0_28[0]), .b(u_csamul_cska32_fa1_27_xor1[0]), .cin(u_csamul_cska32_fa0_27_or0[0]), .fa_xor1(u_csamul_cska32_fa0_28_xor1), .fa_or0(u_csamul_cska32_fa0_28_or0));
  and_gate and_gate_u_csamul_cska32_and1_28(.a(a[1]), .b(b[28]), .out(u_csamul_cska32_and1_28));
  fa fa_u_csamul_cska32_fa1_28_out(.a(u_csamul_cska32_and1_28[0]), .b(u_csamul_cska32_fa2_27_xor1[0]), .cin(u_csamul_cska32_fa1_27_or0[0]), .fa_xor1(u_csamul_cska32_fa1_28_xor1), .fa_or0(u_csamul_cska32_fa1_28_or0));
  and_gate and_gate_u_csamul_cska32_and2_28(.a(a[2]), .b(b[28]), .out(u_csamul_cska32_and2_28));
  fa fa_u_csamul_cska32_fa2_28_out(.a(u_csamul_cska32_and2_28[0]), .b(u_csamul_cska32_fa3_27_xor1[0]), .cin(u_csamul_cska32_fa2_27_or0[0]), .fa_xor1(u_csamul_cska32_fa2_28_xor1), .fa_or0(u_csamul_cska32_fa2_28_or0));
  and_gate and_gate_u_csamul_cska32_and3_28(.a(a[3]), .b(b[28]), .out(u_csamul_cska32_and3_28));
  fa fa_u_csamul_cska32_fa3_28_out(.a(u_csamul_cska32_and3_28[0]), .b(u_csamul_cska32_fa4_27_xor1[0]), .cin(u_csamul_cska32_fa3_27_or0[0]), .fa_xor1(u_csamul_cska32_fa3_28_xor1), .fa_or0(u_csamul_cska32_fa3_28_or0));
  and_gate and_gate_u_csamul_cska32_and4_28(.a(a[4]), .b(b[28]), .out(u_csamul_cska32_and4_28));
  fa fa_u_csamul_cska32_fa4_28_out(.a(u_csamul_cska32_and4_28[0]), .b(u_csamul_cska32_fa5_27_xor1[0]), .cin(u_csamul_cska32_fa4_27_or0[0]), .fa_xor1(u_csamul_cska32_fa4_28_xor1), .fa_or0(u_csamul_cska32_fa4_28_or0));
  and_gate and_gate_u_csamul_cska32_and5_28(.a(a[5]), .b(b[28]), .out(u_csamul_cska32_and5_28));
  fa fa_u_csamul_cska32_fa5_28_out(.a(u_csamul_cska32_and5_28[0]), .b(u_csamul_cska32_fa6_27_xor1[0]), .cin(u_csamul_cska32_fa5_27_or0[0]), .fa_xor1(u_csamul_cska32_fa5_28_xor1), .fa_or0(u_csamul_cska32_fa5_28_or0));
  and_gate and_gate_u_csamul_cska32_and6_28(.a(a[6]), .b(b[28]), .out(u_csamul_cska32_and6_28));
  fa fa_u_csamul_cska32_fa6_28_out(.a(u_csamul_cska32_and6_28[0]), .b(u_csamul_cska32_fa7_27_xor1[0]), .cin(u_csamul_cska32_fa6_27_or0[0]), .fa_xor1(u_csamul_cska32_fa6_28_xor1), .fa_or0(u_csamul_cska32_fa6_28_or0));
  and_gate and_gate_u_csamul_cska32_and7_28(.a(a[7]), .b(b[28]), .out(u_csamul_cska32_and7_28));
  fa fa_u_csamul_cska32_fa7_28_out(.a(u_csamul_cska32_and7_28[0]), .b(u_csamul_cska32_fa8_27_xor1[0]), .cin(u_csamul_cska32_fa7_27_or0[0]), .fa_xor1(u_csamul_cska32_fa7_28_xor1), .fa_or0(u_csamul_cska32_fa7_28_or0));
  and_gate and_gate_u_csamul_cska32_and8_28(.a(a[8]), .b(b[28]), .out(u_csamul_cska32_and8_28));
  fa fa_u_csamul_cska32_fa8_28_out(.a(u_csamul_cska32_and8_28[0]), .b(u_csamul_cska32_fa9_27_xor1[0]), .cin(u_csamul_cska32_fa8_27_or0[0]), .fa_xor1(u_csamul_cska32_fa8_28_xor1), .fa_or0(u_csamul_cska32_fa8_28_or0));
  and_gate and_gate_u_csamul_cska32_and9_28(.a(a[9]), .b(b[28]), .out(u_csamul_cska32_and9_28));
  fa fa_u_csamul_cska32_fa9_28_out(.a(u_csamul_cska32_and9_28[0]), .b(u_csamul_cska32_fa10_27_xor1[0]), .cin(u_csamul_cska32_fa9_27_or0[0]), .fa_xor1(u_csamul_cska32_fa9_28_xor1), .fa_or0(u_csamul_cska32_fa9_28_or0));
  and_gate and_gate_u_csamul_cska32_and10_28(.a(a[10]), .b(b[28]), .out(u_csamul_cska32_and10_28));
  fa fa_u_csamul_cska32_fa10_28_out(.a(u_csamul_cska32_and10_28[0]), .b(u_csamul_cska32_fa11_27_xor1[0]), .cin(u_csamul_cska32_fa10_27_or0[0]), .fa_xor1(u_csamul_cska32_fa10_28_xor1), .fa_or0(u_csamul_cska32_fa10_28_or0));
  and_gate and_gate_u_csamul_cska32_and11_28(.a(a[11]), .b(b[28]), .out(u_csamul_cska32_and11_28));
  fa fa_u_csamul_cska32_fa11_28_out(.a(u_csamul_cska32_and11_28[0]), .b(u_csamul_cska32_fa12_27_xor1[0]), .cin(u_csamul_cska32_fa11_27_or0[0]), .fa_xor1(u_csamul_cska32_fa11_28_xor1), .fa_or0(u_csamul_cska32_fa11_28_or0));
  and_gate and_gate_u_csamul_cska32_and12_28(.a(a[12]), .b(b[28]), .out(u_csamul_cska32_and12_28));
  fa fa_u_csamul_cska32_fa12_28_out(.a(u_csamul_cska32_and12_28[0]), .b(u_csamul_cska32_fa13_27_xor1[0]), .cin(u_csamul_cska32_fa12_27_or0[0]), .fa_xor1(u_csamul_cska32_fa12_28_xor1), .fa_or0(u_csamul_cska32_fa12_28_or0));
  and_gate and_gate_u_csamul_cska32_and13_28(.a(a[13]), .b(b[28]), .out(u_csamul_cska32_and13_28));
  fa fa_u_csamul_cska32_fa13_28_out(.a(u_csamul_cska32_and13_28[0]), .b(u_csamul_cska32_fa14_27_xor1[0]), .cin(u_csamul_cska32_fa13_27_or0[0]), .fa_xor1(u_csamul_cska32_fa13_28_xor1), .fa_or0(u_csamul_cska32_fa13_28_or0));
  and_gate and_gate_u_csamul_cska32_and14_28(.a(a[14]), .b(b[28]), .out(u_csamul_cska32_and14_28));
  fa fa_u_csamul_cska32_fa14_28_out(.a(u_csamul_cska32_and14_28[0]), .b(u_csamul_cska32_fa15_27_xor1[0]), .cin(u_csamul_cska32_fa14_27_or0[0]), .fa_xor1(u_csamul_cska32_fa14_28_xor1), .fa_or0(u_csamul_cska32_fa14_28_or0));
  and_gate and_gate_u_csamul_cska32_and15_28(.a(a[15]), .b(b[28]), .out(u_csamul_cska32_and15_28));
  fa fa_u_csamul_cska32_fa15_28_out(.a(u_csamul_cska32_and15_28[0]), .b(u_csamul_cska32_fa16_27_xor1[0]), .cin(u_csamul_cska32_fa15_27_or0[0]), .fa_xor1(u_csamul_cska32_fa15_28_xor1), .fa_or0(u_csamul_cska32_fa15_28_or0));
  and_gate and_gate_u_csamul_cska32_and16_28(.a(a[16]), .b(b[28]), .out(u_csamul_cska32_and16_28));
  fa fa_u_csamul_cska32_fa16_28_out(.a(u_csamul_cska32_and16_28[0]), .b(u_csamul_cska32_fa17_27_xor1[0]), .cin(u_csamul_cska32_fa16_27_or0[0]), .fa_xor1(u_csamul_cska32_fa16_28_xor1), .fa_or0(u_csamul_cska32_fa16_28_or0));
  and_gate and_gate_u_csamul_cska32_and17_28(.a(a[17]), .b(b[28]), .out(u_csamul_cska32_and17_28));
  fa fa_u_csamul_cska32_fa17_28_out(.a(u_csamul_cska32_and17_28[0]), .b(u_csamul_cska32_fa18_27_xor1[0]), .cin(u_csamul_cska32_fa17_27_or0[0]), .fa_xor1(u_csamul_cska32_fa17_28_xor1), .fa_or0(u_csamul_cska32_fa17_28_or0));
  and_gate and_gate_u_csamul_cska32_and18_28(.a(a[18]), .b(b[28]), .out(u_csamul_cska32_and18_28));
  fa fa_u_csamul_cska32_fa18_28_out(.a(u_csamul_cska32_and18_28[0]), .b(u_csamul_cska32_fa19_27_xor1[0]), .cin(u_csamul_cska32_fa18_27_or0[0]), .fa_xor1(u_csamul_cska32_fa18_28_xor1), .fa_or0(u_csamul_cska32_fa18_28_or0));
  and_gate and_gate_u_csamul_cska32_and19_28(.a(a[19]), .b(b[28]), .out(u_csamul_cska32_and19_28));
  fa fa_u_csamul_cska32_fa19_28_out(.a(u_csamul_cska32_and19_28[0]), .b(u_csamul_cska32_fa20_27_xor1[0]), .cin(u_csamul_cska32_fa19_27_or0[0]), .fa_xor1(u_csamul_cska32_fa19_28_xor1), .fa_or0(u_csamul_cska32_fa19_28_or0));
  and_gate and_gate_u_csamul_cska32_and20_28(.a(a[20]), .b(b[28]), .out(u_csamul_cska32_and20_28));
  fa fa_u_csamul_cska32_fa20_28_out(.a(u_csamul_cska32_and20_28[0]), .b(u_csamul_cska32_fa21_27_xor1[0]), .cin(u_csamul_cska32_fa20_27_or0[0]), .fa_xor1(u_csamul_cska32_fa20_28_xor1), .fa_or0(u_csamul_cska32_fa20_28_or0));
  and_gate and_gate_u_csamul_cska32_and21_28(.a(a[21]), .b(b[28]), .out(u_csamul_cska32_and21_28));
  fa fa_u_csamul_cska32_fa21_28_out(.a(u_csamul_cska32_and21_28[0]), .b(u_csamul_cska32_fa22_27_xor1[0]), .cin(u_csamul_cska32_fa21_27_or0[0]), .fa_xor1(u_csamul_cska32_fa21_28_xor1), .fa_or0(u_csamul_cska32_fa21_28_or0));
  and_gate and_gate_u_csamul_cska32_and22_28(.a(a[22]), .b(b[28]), .out(u_csamul_cska32_and22_28));
  fa fa_u_csamul_cska32_fa22_28_out(.a(u_csamul_cska32_and22_28[0]), .b(u_csamul_cska32_fa23_27_xor1[0]), .cin(u_csamul_cska32_fa22_27_or0[0]), .fa_xor1(u_csamul_cska32_fa22_28_xor1), .fa_or0(u_csamul_cska32_fa22_28_or0));
  and_gate and_gate_u_csamul_cska32_and23_28(.a(a[23]), .b(b[28]), .out(u_csamul_cska32_and23_28));
  fa fa_u_csamul_cska32_fa23_28_out(.a(u_csamul_cska32_and23_28[0]), .b(u_csamul_cska32_fa24_27_xor1[0]), .cin(u_csamul_cska32_fa23_27_or0[0]), .fa_xor1(u_csamul_cska32_fa23_28_xor1), .fa_or0(u_csamul_cska32_fa23_28_or0));
  and_gate and_gate_u_csamul_cska32_and24_28(.a(a[24]), .b(b[28]), .out(u_csamul_cska32_and24_28));
  fa fa_u_csamul_cska32_fa24_28_out(.a(u_csamul_cska32_and24_28[0]), .b(u_csamul_cska32_fa25_27_xor1[0]), .cin(u_csamul_cska32_fa24_27_or0[0]), .fa_xor1(u_csamul_cska32_fa24_28_xor1), .fa_or0(u_csamul_cska32_fa24_28_or0));
  and_gate and_gate_u_csamul_cska32_and25_28(.a(a[25]), .b(b[28]), .out(u_csamul_cska32_and25_28));
  fa fa_u_csamul_cska32_fa25_28_out(.a(u_csamul_cska32_and25_28[0]), .b(u_csamul_cska32_fa26_27_xor1[0]), .cin(u_csamul_cska32_fa25_27_or0[0]), .fa_xor1(u_csamul_cska32_fa25_28_xor1), .fa_or0(u_csamul_cska32_fa25_28_or0));
  and_gate and_gate_u_csamul_cska32_and26_28(.a(a[26]), .b(b[28]), .out(u_csamul_cska32_and26_28));
  fa fa_u_csamul_cska32_fa26_28_out(.a(u_csamul_cska32_and26_28[0]), .b(u_csamul_cska32_fa27_27_xor1[0]), .cin(u_csamul_cska32_fa26_27_or0[0]), .fa_xor1(u_csamul_cska32_fa26_28_xor1), .fa_or0(u_csamul_cska32_fa26_28_or0));
  and_gate and_gate_u_csamul_cska32_and27_28(.a(a[27]), .b(b[28]), .out(u_csamul_cska32_and27_28));
  fa fa_u_csamul_cska32_fa27_28_out(.a(u_csamul_cska32_and27_28[0]), .b(u_csamul_cska32_fa28_27_xor1[0]), .cin(u_csamul_cska32_fa27_27_or0[0]), .fa_xor1(u_csamul_cska32_fa27_28_xor1), .fa_or0(u_csamul_cska32_fa27_28_or0));
  and_gate and_gate_u_csamul_cska32_and28_28(.a(a[28]), .b(b[28]), .out(u_csamul_cska32_and28_28));
  fa fa_u_csamul_cska32_fa28_28_out(.a(u_csamul_cska32_and28_28[0]), .b(u_csamul_cska32_fa29_27_xor1[0]), .cin(u_csamul_cska32_fa28_27_or0[0]), .fa_xor1(u_csamul_cska32_fa28_28_xor1), .fa_or0(u_csamul_cska32_fa28_28_or0));
  and_gate and_gate_u_csamul_cska32_and29_28(.a(a[29]), .b(b[28]), .out(u_csamul_cska32_and29_28));
  fa fa_u_csamul_cska32_fa29_28_out(.a(u_csamul_cska32_and29_28[0]), .b(u_csamul_cska32_fa30_27_xor1[0]), .cin(u_csamul_cska32_fa29_27_or0[0]), .fa_xor1(u_csamul_cska32_fa29_28_xor1), .fa_or0(u_csamul_cska32_fa29_28_or0));
  and_gate and_gate_u_csamul_cska32_and30_28(.a(a[30]), .b(b[28]), .out(u_csamul_cska32_and30_28));
  fa fa_u_csamul_cska32_fa30_28_out(.a(u_csamul_cska32_and30_28[0]), .b(u_csamul_cska32_and31_27[0]), .cin(u_csamul_cska32_fa30_27_or0[0]), .fa_xor1(u_csamul_cska32_fa30_28_xor1), .fa_or0(u_csamul_cska32_fa30_28_or0));
  and_gate and_gate_u_csamul_cska32_and31_28(.a(a[31]), .b(b[28]), .out(u_csamul_cska32_and31_28));
  and_gate and_gate_u_csamul_cska32_and0_29(.a(a[0]), .b(b[29]), .out(u_csamul_cska32_and0_29));
  fa fa_u_csamul_cska32_fa0_29_out(.a(u_csamul_cska32_and0_29[0]), .b(u_csamul_cska32_fa1_28_xor1[0]), .cin(u_csamul_cska32_fa0_28_or0[0]), .fa_xor1(u_csamul_cska32_fa0_29_xor1), .fa_or0(u_csamul_cska32_fa0_29_or0));
  and_gate and_gate_u_csamul_cska32_and1_29(.a(a[1]), .b(b[29]), .out(u_csamul_cska32_and1_29));
  fa fa_u_csamul_cska32_fa1_29_out(.a(u_csamul_cska32_and1_29[0]), .b(u_csamul_cska32_fa2_28_xor1[0]), .cin(u_csamul_cska32_fa1_28_or0[0]), .fa_xor1(u_csamul_cska32_fa1_29_xor1), .fa_or0(u_csamul_cska32_fa1_29_or0));
  and_gate and_gate_u_csamul_cska32_and2_29(.a(a[2]), .b(b[29]), .out(u_csamul_cska32_and2_29));
  fa fa_u_csamul_cska32_fa2_29_out(.a(u_csamul_cska32_and2_29[0]), .b(u_csamul_cska32_fa3_28_xor1[0]), .cin(u_csamul_cska32_fa2_28_or0[0]), .fa_xor1(u_csamul_cska32_fa2_29_xor1), .fa_or0(u_csamul_cska32_fa2_29_or0));
  and_gate and_gate_u_csamul_cska32_and3_29(.a(a[3]), .b(b[29]), .out(u_csamul_cska32_and3_29));
  fa fa_u_csamul_cska32_fa3_29_out(.a(u_csamul_cska32_and3_29[0]), .b(u_csamul_cska32_fa4_28_xor1[0]), .cin(u_csamul_cska32_fa3_28_or0[0]), .fa_xor1(u_csamul_cska32_fa3_29_xor1), .fa_or0(u_csamul_cska32_fa3_29_or0));
  and_gate and_gate_u_csamul_cska32_and4_29(.a(a[4]), .b(b[29]), .out(u_csamul_cska32_and4_29));
  fa fa_u_csamul_cska32_fa4_29_out(.a(u_csamul_cska32_and4_29[0]), .b(u_csamul_cska32_fa5_28_xor1[0]), .cin(u_csamul_cska32_fa4_28_or0[0]), .fa_xor1(u_csamul_cska32_fa4_29_xor1), .fa_or0(u_csamul_cska32_fa4_29_or0));
  and_gate and_gate_u_csamul_cska32_and5_29(.a(a[5]), .b(b[29]), .out(u_csamul_cska32_and5_29));
  fa fa_u_csamul_cska32_fa5_29_out(.a(u_csamul_cska32_and5_29[0]), .b(u_csamul_cska32_fa6_28_xor1[0]), .cin(u_csamul_cska32_fa5_28_or0[0]), .fa_xor1(u_csamul_cska32_fa5_29_xor1), .fa_or0(u_csamul_cska32_fa5_29_or0));
  and_gate and_gate_u_csamul_cska32_and6_29(.a(a[6]), .b(b[29]), .out(u_csamul_cska32_and6_29));
  fa fa_u_csamul_cska32_fa6_29_out(.a(u_csamul_cska32_and6_29[0]), .b(u_csamul_cska32_fa7_28_xor1[0]), .cin(u_csamul_cska32_fa6_28_or0[0]), .fa_xor1(u_csamul_cska32_fa6_29_xor1), .fa_or0(u_csamul_cska32_fa6_29_or0));
  and_gate and_gate_u_csamul_cska32_and7_29(.a(a[7]), .b(b[29]), .out(u_csamul_cska32_and7_29));
  fa fa_u_csamul_cska32_fa7_29_out(.a(u_csamul_cska32_and7_29[0]), .b(u_csamul_cska32_fa8_28_xor1[0]), .cin(u_csamul_cska32_fa7_28_or0[0]), .fa_xor1(u_csamul_cska32_fa7_29_xor1), .fa_or0(u_csamul_cska32_fa7_29_or0));
  and_gate and_gate_u_csamul_cska32_and8_29(.a(a[8]), .b(b[29]), .out(u_csamul_cska32_and8_29));
  fa fa_u_csamul_cska32_fa8_29_out(.a(u_csamul_cska32_and8_29[0]), .b(u_csamul_cska32_fa9_28_xor1[0]), .cin(u_csamul_cska32_fa8_28_or0[0]), .fa_xor1(u_csamul_cska32_fa8_29_xor1), .fa_or0(u_csamul_cska32_fa8_29_or0));
  and_gate and_gate_u_csamul_cska32_and9_29(.a(a[9]), .b(b[29]), .out(u_csamul_cska32_and9_29));
  fa fa_u_csamul_cska32_fa9_29_out(.a(u_csamul_cska32_and9_29[0]), .b(u_csamul_cska32_fa10_28_xor1[0]), .cin(u_csamul_cska32_fa9_28_or0[0]), .fa_xor1(u_csamul_cska32_fa9_29_xor1), .fa_or0(u_csamul_cska32_fa9_29_or0));
  and_gate and_gate_u_csamul_cska32_and10_29(.a(a[10]), .b(b[29]), .out(u_csamul_cska32_and10_29));
  fa fa_u_csamul_cska32_fa10_29_out(.a(u_csamul_cska32_and10_29[0]), .b(u_csamul_cska32_fa11_28_xor1[0]), .cin(u_csamul_cska32_fa10_28_or0[0]), .fa_xor1(u_csamul_cska32_fa10_29_xor1), .fa_or0(u_csamul_cska32_fa10_29_or0));
  and_gate and_gate_u_csamul_cska32_and11_29(.a(a[11]), .b(b[29]), .out(u_csamul_cska32_and11_29));
  fa fa_u_csamul_cska32_fa11_29_out(.a(u_csamul_cska32_and11_29[0]), .b(u_csamul_cska32_fa12_28_xor1[0]), .cin(u_csamul_cska32_fa11_28_or0[0]), .fa_xor1(u_csamul_cska32_fa11_29_xor1), .fa_or0(u_csamul_cska32_fa11_29_or0));
  and_gate and_gate_u_csamul_cska32_and12_29(.a(a[12]), .b(b[29]), .out(u_csamul_cska32_and12_29));
  fa fa_u_csamul_cska32_fa12_29_out(.a(u_csamul_cska32_and12_29[0]), .b(u_csamul_cska32_fa13_28_xor1[0]), .cin(u_csamul_cska32_fa12_28_or0[0]), .fa_xor1(u_csamul_cska32_fa12_29_xor1), .fa_or0(u_csamul_cska32_fa12_29_or0));
  and_gate and_gate_u_csamul_cska32_and13_29(.a(a[13]), .b(b[29]), .out(u_csamul_cska32_and13_29));
  fa fa_u_csamul_cska32_fa13_29_out(.a(u_csamul_cska32_and13_29[0]), .b(u_csamul_cska32_fa14_28_xor1[0]), .cin(u_csamul_cska32_fa13_28_or0[0]), .fa_xor1(u_csamul_cska32_fa13_29_xor1), .fa_or0(u_csamul_cska32_fa13_29_or0));
  and_gate and_gate_u_csamul_cska32_and14_29(.a(a[14]), .b(b[29]), .out(u_csamul_cska32_and14_29));
  fa fa_u_csamul_cska32_fa14_29_out(.a(u_csamul_cska32_and14_29[0]), .b(u_csamul_cska32_fa15_28_xor1[0]), .cin(u_csamul_cska32_fa14_28_or0[0]), .fa_xor1(u_csamul_cska32_fa14_29_xor1), .fa_or0(u_csamul_cska32_fa14_29_or0));
  and_gate and_gate_u_csamul_cska32_and15_29(.a(a[15]), .b(b[29]), .out(u_csamul_cska32_and15_29));
  fa fa_u_csamul_cska32_fa15_29_out(.a(u_csamul_cska32_and15_29[0]), .b(u_csamul_cska32_fa16_28_xor1[0]), .cin(u_csamul_cska32_fa15_28_or0[0]), .fa_xor1(u_csamul_cska32_fa15_29_xor1), .fa_or0(u_csamul_cska32_fa15_29_or0));
  and_gate and_gate_u_csamul_cska32_and16_29(.a(a[16]), .b(b[29]), .out(u_csamul_cska32_and16_29));
  fa fa_u_csamul_cska32_fa16_29_out(.a(u_csamul_cska32_and16_29[0]), .b(u_csamul_cska32_fa17_28_xor1[0]), .cin(u_csamul_cska32_fa16_28_or0[0]), .fa_xor1(u_csamul_cska32_fa16_29_xor1), .fa_or0(u_csamul_cska32_fa16_29_or0));
  and_gate and_gate_u_csamul_cska32_and17_29(.a(a[17]), .b(b[29]), .out(u_csamul_cska32_and17_29));
  fa fa_u_csamul_cska32_fa17_29_out(.a(u_csamul_cska32_and17_29[0]), .b(u_csamul_cska32_fa18_28_xor1[0]), .cin(u_csamul_cska32_fa17_28_or0[0]), .fa_xor1(u_csamul_cska32_fa17_29_xor1), .fa_or0(u_csamul_cska32_fa17_29_or0));
  and_gate and_gate_u_csamul_cska32_and18_29(.a(a[18]), .b(b[29]), .out(u_csamul_cska32_and18_29));
  fa fa_u_csamul_cska32_fa18_29_out(.a(u_csamul_cska32_and18_29[0]), .b(u_csamul_cska32_fa19_28_xor1[0]), .cin(u_csamul_cska32_fa18_28_or0[0]), .fa_xor1(u_csamul_cska32_fa18_29_xor1), .fa_or0(u_csamul_cska32_fa18_29_or0));
  and_gate and_gate_u_csamul_cska32_and19_29(.a(a[19]), .b(b[29]), .out(u_csamul_cska32_and19_29));
  fa fa_u_csamul_cska32_fa19_29_out(.a(u_csamul_cska32_and19_29[0]), .b(u_csamul_cska32_fa20_28_xor1[0]), .cin(u_csamul_cska32_fa19_28_or0[0]), .fa_xor1(u_csamul_cska32_fa19_29_xor1), .fa_or0(u_csamul_cska32_fa19_29_or0));
  and_gate and_gate_u_csamul_cska32_and20_29(.a(a[20]), .b(b[29]), .out(u_csamul_cska32_and20_29));
  fa fa_u_csamul_cska32_fa20_29_out(.a(u_csamul_cska32_and20_29[0]), .b(u_csamul_cska32_fa21_28_xor1[0]), .cin(u_csamul_cska32_fa20_28_or0[0]), .fa_xor1(u_csamul_cska32_fa20_29_xor1), .fa_or0(u_csamul_cska32_fa20_29_or0));
  and_gate and_gate_u_csamul_cska32_and21_29(.a(a[21]), .b(b[29]), .out(u_csamul_cska32_and21_29));
  fa fa_u_csamul_cska32_fa21_29_out(.a(u_csamul_cska32_and21_29[0]), .b(u_csamul_cska32_fa22_28_xor1[0]), .cin(u_csamul_cska32_fa21_28_or0[0]), .fa_xor1(u_csamul_cska32_fa21_29_xor1), .fa_or0(u_csamul_cska32_fa21_29_or0));
  and_gate and_gate_u_csamul_cska32_and22_29(.a(a[22]), .b(b[29]), .out(u_csamul_cska32_and22_29));
  fa fa_u_csamul_cska32_fa22_29_out(.a(u_csamul_cska32_and22_29[0]), .b(u_csamul_cska32_fa23_28_xor1[0]), .cin(u_csamul_cska32_fa22_28_or0[0]), .fa_xor1(u_csamul_cska32_fa22_29_xor1), .fa_or0(u_csamul_cska32_fa22_29_or0));
  and_gate and_gate_u_csamul_cska32_and23_29(.a(a[23]), .b(b[29]), .out(u_csamul_cska32_and23_29));
  fa fa_u_csamul_cska32_fa23_29_out(.a(u_csamul_cska32_and23_29[0]), .b(u_csamul_cska32_fa24_28_xor1[0]), .cin(u_csamul_cska32_fa23_28_or0[0]), .fa_xor1(u_csamul_cska32_fa23_29_xor1), .fa_or0(u_csamul_cska32_fa23_29_or0));
  and_gate and_gate_u_csamul_cska32_and24_29(.a(a[24]), .b(b[29]), .out(u_csamul_cska32_and24_29));
  fa fa_u_csamul_cska32_fa24_29_out(.a(u_csamul_cska32_and24_29[0]), .b(u_csamul_cska32_fa25_28_xor1[0]), .cin(u_csamul_cska32_fa24_28_or0[0]), .fa_xor1(u_csamul_cska32_fa24_29_xor1), .fa_or0(u_csamul_cska32_fa24_29_or0));
  and_gate and_gate_u_csamul_cska32_and25_29(.a(a[25]), .b(b[29]), .out(u_csamul_cska32_and25_29));
  fa fa_u_csamul_cska32_fa25_29_out(.a(u_csamul_cska32_and25_29[0]), .b(u_csamul_cska32_fa26_28_xor1[0]), .cin(u_csamul_cska32_fa25_28_or0[0]), .fa_xor1(u_csamul_cska32_fa25_29_xor1), .fa_or0(u_csamul_cska32_fa25_29_or0));
  and_gate and_gate_u_csamul_cska32_and26_29(.a(a[26]), .b(b[29]), .out(u_csamul_cska32_and26_29));
  fa fa_u_csamul_cska32_fa26_29_out(.a(u_csamul_cska32_and26_29[0]), .b(u_csamul_cska32_fa27_28_xor1[0]), .cin(u_csamul_cska32_fa26_28_or0[0]), .fa_xor1(u_csamul_cska32_fa26_29_xor1), .fa_or0(u_csamul_cska32_fa26_29_or0));
  and_gate and_gate_u_csamul_cska32_and27_29(.a(a[27]), .b(b[29]), .out(u_csamul_cska32_and27_29));
  fa fa_u_csamul_cska32_fa27_29_out(.a(u_csamul_cska32_and27_29[0]), .b(u_csamul_cska32_fa28_28_xor1[0]), .cin(u_csamul_cska32_fa27_28_or0[0]), .fa_xor1(u_csamul_cska32_fa27_29_xor1), .fa_or0(u_csamul_cska32_fa27_29_or0));
  and_gate and_gate_u_csamul_cska32_and28_29(.a(a[28]), .b(b[29]), .out(u_csamul_cska32_and28_29));
  fa fa_u_csamul_cska32_fa28_29_out(.a(u_csamul_cska32_and28_29[0]), .b(u_csamul_cska32_fa29_28_xor1[0]), .cin(u_csamul_cska32_fa28_28_or0[0]), .fa_xor1(u_csamul_cska32_fa28_29_xor1), .fa_or0(u_csamul_cska32_fa28_29_or0));
  and_gate and_gate_u_csamul_cska32_and29_29(.a(a[29]), .b(b[29]), .out(u_csamul_cska32_and29_29));
  fa fa_u_csamul_cska32_fa29_29_out(.a(u_csamul_cska32_and29_29[0]), .b(u_csamul_cska32_fa30_28_xor1[0]), .cin(u_csamul_cska32_fa29_28_or0[0]), .fa_xor1(u_csamul_cska32_fa29_29_xor1), .fa_or0(u_csamul_cska32_fa29_29_or0));
  and_gate and_gate_u_csamul_cska32_and30_29(.a(a[30]), .b(b[29]), .out(u_csamul_cska32_and30_29));
  fa fa_u_csamul_cska32_fa30_29_out(.a(u_csamul_cska32_and30_29[0]), .b(u_csamul_cska32_and31_28[0]), .cin(u_csamul_cska32_fa30_28_or0[0]), .fa_xor1(u_csamul_cska32_fa30_29_xor1), .fa_or0(u_csamul_cska32_fa30_29_or0));
  and_gate and_gate_u_csamul_cska32_and31_29(.a(a[31]), .b(b[29]), .out(u_csamul_cska32_and31_29));
  and_gate and_gate_u_csamul_cska32_and0_30(.a(a[0]), .b(b[30]), .out(u_csamul_cska32_and0_30));
  fa fa_u_csamul_cska32_fa0_30_out(.a(u_csamul_cska32_and0_30[0]), .b(u_csamul_cska32_fa1_29_xor1[0]), .cin(u_csamul_cska32_fa0_29_or0[0]), .fa_xor1(u_csamul_cska32_fa0_30_xor1), .fa_or0(u_csamul_cska32_fa0_30_or0));
  and_gate and_gate_u_csamul_cska32_and1_30(.a(a[1]), .b(b[30]), .out(u_csamul_cska32_and1_30));
  fa fa_u_csamul_cska32_fa1_30_out(.a(u_csamul_cska32_and1_30[0]), .b(u_csamul_cska32_fa2_29_xor1[0]), .cin(u_csamul_cska32_fa1_29_or0[0]), .fa_xor1(u_csamul_cska32_fa1_30_xor1), .fa_or0(u_csamul_cska32_fa1_30_or0));
  and_gate and_gate_u_csamul_cska32_and2_30(.a(a[2]), .b(b[30]), .out(u_csamul_cska32_and2_30));
  fa fa_u_csamul_cska32_fa2_30_out(.a(u_csamul_cska32_and2_30[0]), .b(u_csamul_cska32_fa3_29_xor1[0]), .cin(u_csamul_cska32_fa2_29_or0[0]), .fa_xor1(u_csamul_cska32_fa2_30_xor1), .fa_or0(u_csamul_cska32_fa2_30_or0));
  and_gate and_gate_u_csamul_cska32_and3_30(.a(a[3]), .b(b[30]), .out(u_csamul_cska32_and3_30));
  fa fa_u_csamul_cska32_fa3_30_out(.a(u_csamul_cska32_and3_30[0]), .b(u_csamul_cska32_fa4_29_xor1[0]), .cin(u_csamul_cska32_fa3_29_or0[0]), .fa_xor1(u_csamul_cska32_fa3_30_xor1), .fa_or0(u_csamul_cska32_fa3_30_or0));
  and_gate and_gate_u_csamul_cska32_and4_30(.a(a[4]), .b(b[30]), .out(u_csamul_cska32_and4_30));
  fa fa_u_csamul_cska32_fa4_30_out(.a(u_csamul_cska32_and4_30[0]), .b(u_csamul_cska32_fa5_29_xor1[0]), .cin(u_csamul_cska32_fa4_29_or0[0]), .fa_xor1(u_csamul_cska32_fa4_30_xor1), .fa_or0(u_csamul_cska32_fa4_30_or0));
  and_gate and_gate_u_csamul_cska32_and5_30(.a(a[5]), .b(b[30]), .out(u_csamul_cska32_and5_30));
  fa fa_u_csamul_cska32_fa5_30_out(.a(u_csamul_cska32_and5_30[0]), .b(u_csamul_cska32_fa6_29_xor1[0]), .cin(u_csamul_cska32_fa5_29_or0[0]), .fa_xor1(u_csamul_cska32_fa5_30_xor1), .fa_or0(u_csamul_cska32_fa5_30_or0));
  and_gate and_gate_u_csamul_cska32_and6_30(.a(a[6]), .b(b[30]), .out(u_csamul_cska32_and6_30));
  fa fa_u_csamul_cska32_fa6_30_out(.a(u_csamul_cska32_and6_30[0]), .b(u_csamul_cska32_fa7_29_xor1[0]), .cin(u_csamul_cska32_fa6_29_or0[0]), .fa_xor1(u_csamul_cska32_fa6_30_xor1), .fa_or0(u_csamul_cska32_fa6_30_or0));
  and_gate and_gate_u_csamul_cska32_and7_30(.a(a[7]), .b(b[30]), .out(u_csamul_cska32_and7_30));
  fa fa_u_csamul_cska32_fa7_30_out(.a(u_csamul_cska32_and7_30[0]), .b(u_csamul_cska32_fa8_29_xor1[0]), .cin(u_csamul_cska32_fa7_29_or0[0]), .fa_xor1(u_csamul_cska32_fa7_30_xor1), .fa_or0(u_csamul_cska32_fa7_30_or0));
  and_gate and_gate_u_csamul_cska32_and8_30(.a(a[8]), .b(b[30]), .out(u_csamul_cska32_and8_30));
  fa fa_u_csamul_cska32_fa8_30_out(.a(u_csamul_cska32_and8_30[0]), .b(u_csamul_cska32_fa9_29_xor1[0]), .cin(u_csamul_cska32_fa8_29_or0[0]), .fa_xor1(u_csamul_cska32_fa8_30_xor1), .fa_or0(u_csamul_cska32_fa8_30_or0));
  and_gate and_gate_u_csamul_cska32_and9_30(.a(a[9]), .b(b[30]), .out(u_csamul_cska32_and9_30));
  fa fa_u_csamul_cska32_fa9_30_out(.a(u_csamul_cska32_and9_30[0]), .b(u_csamul_cska32_fa10_29_xor1[0]), .cin(u_csamul_cska32_fa9_29_or0[0]), .fa_xor1(u_csamul_cska32_fa9_30_xor1), .fa_or0(u_csamul_cska32_fa9_30_or0));
  and_gate and_gate_u_csamul_cska32_and10_30(.a(a[10]), .b(b[30]), .out(u_csamul_cska32_and10_30));
  fa fa_u_csamul_cska32_fa10_30_out(.a(u_csamul_cska32_and10_30[0]), .b(u_csamul_cska32_fa11_29_xor1[0]), .cin(u_csamul_cska32_fa10_29_or0[0]), .fa_xor1(u_csamul_cska32_fa10_30_xor1), .fa_or0(u_csamul_cska32_fa10_30_or0));
  and_gate and_gate_u_csamul_cska32_and11_30(.a(a[11]), .b(b[30]), .out(u_csamul_cska32_and11_30));
  fa fa_u_csamul_cska32_fa11_30_out(.a(u_csamul_cska32_and11_30[0]), .b(u_csamul_cska32_fa12_29_xor1[0]), .cin(u_csamul_cska32_fa11_29_or0[0]), .fa_xor1(u_csamul_cska32_fa11_30_xor1), .fa_or0(u_csamul_cska32_fa11_30_or0));
  and_gate and_gate_u_csamul_cska32_and12_30(.a(a[12]), .b(b[30]), .out(u_csamul_cska32_and12_30));
  fa fa_u_csamul_cska32_fa12_30_out(.a(u_csamul_cska32_and12_30[0]), .b(u_csamul_cska32_fa13_29_xor1[0]), .cin(u_csamul_cska32_fa12_29_or0[0]), .fa_xor1(u_csamul_cska32_fa12_30_xor1), .fa_or0(u_csamul_cska32_fa12_30_or0));
  and_gate and_gate_u_csamul_cska32_and13_30(.a(a[13]), .b(b[30]), .out(u_csamul_cska32_and13_30));
  fa fa_u_csamul_cska32_fa13_30_out(.a(u_csamul_cska32_and13_30[0]), .b(u_csamul_cska32_fa14_29_xor1[0]), .cin(u_csamul_cska32_fa13_29_or0[0]), .fa_xor1(u_csamul_cska32_fa13_30_xor1), .fa_or0(u_csamul_cska32_fa13_30_or0));
  and_gate and_gate_u_csamul_cska32_and14_30(.a(a[14]), .b(b[30]), .out(u_csamul_cska32_and14_30));
  fa fa_u_csamul_cska32_fa14_30_out(.a(u_csamul_cska32_and14_30[0]), .b(u_csamul_cska32_fa15_29_xor1[0]), .cin(u_csamul_cska32_fa14_29_or0[0]), .fa_xor1(u_csamul_cska32_fa14_30_xor1), .fa_or0(u_csamul_cska32_fa14_30_or0));
  and_gate and_gate_u_csamul_cska32_and15_30(.a(a[15]), .b(b[30]), .out(u_csamul_cska32_and15_30));
  fa fa_u_csamul_cska32_fa15_30_out(.a(u_csamul_cska32_and15_30[0]), .b(u_csamul_cska32_fa16_29_xor1[0]), .cin(u_csamul_cska32_fa15_29_or0[0]), .fa_xor1(u_csamul_cska32_fa15_30_xor1), .fa_or0(u_csamul_cska32_fa15_30_or0));
  and_gate and_gate_u_csamul_cska32_and16_30(.a(a[16]), .b(b[30]), .out(u_csamul_cska32_and16_30));
  fa fa_u_csamul_cska32_fa16_30_out(.a(u_csamul_cska32_and16_30[0]), .b(u_csamul_cska32_fa17_29_xor1[0]), .cin(u_csamul_cska32_fa16_29_or0[0]), .fa_xor1(u_csamul_cska32_fa16_30_xor1), .fa_or0(u_csamul_cska32_fa16_30_or0));
  and_gate and_gate_u_csamul_cska32_and17_30(.a(a[17]), .b(b[30]), .out(u_csamul_cska32_and17_30));
  fa fa_u_csamul_cska32_fa17_30_out(.a(u_csamul_cska32_and17_30[0]), .b(u_csamul_cska32_fa18_29_xor1[0]), .cin(u_csamul_cska32_fa17_29_or0[0]), .fa_xor1(u_csamul_cska32_fa17_30_xor1), .fa_or0(u_csamul_cska32_fa17_30_or0));
  and_gate and_gate_u_csamul_cska32_and18_30(.a(a[18]), .b(b[30]), .out(u_csamul_cska32_and18_30));
  fa fa_u_csamul_cska32_fa18_30_out(.a(u_csamul_cska32_and18_30[0]), .b(u_csamul_cska32_fa19_29_xor1[0]), .cin(u_csamul_cska32_fa18_29_or0[0]), .fa_xor1(u_csamul_cska32_fa18_30_xor1), .fa_or0(u_csamul_cska32_fa18_30_or0));
  and_gate and_gate_u_csamul_cska32_and19_30(.a(a[19]), .b(b[30]), .out(u_csamul_cska32_and19_30));
  fa fa_u_csamul_cska32_fa19_30_out(.a(u_csamul_cska32_and19_30[0]), .b(u_csamul_cska32_fa20_29_xor1[0]), .cin(u_csamul_cska32_fa19_29_or0[0]), .fa_xor1(u_csamul_cska32_fa19_30_xor1), .fa_or0(u_csamul_cska32_fa19_30_or0));
  and_gate and_gate_u_csamul_cska32_and20_30(.a(a[20]), .b(b[30]), .out(u_csamul_cska32_and20_30));
  fa fa_u_csamul_cska32_fa20_30_out(.a(u_csamul_cska32_and20_30[0]), .b(u_csamul_cska32_fa21_29_xor1[0]), .cin(u_csamul_cska32_fa20_29_or0[0]), .fa_xor1(u_csamul_cska32_fa20_30_xor1), .fa_or0(u_csamul_cska32_fa20_30_or0));
  and_gate and_gate_u_csamul_cska32_and21_30(.a(a[21]), .b(b[30]), .out(u_csamul_cska32_and21_30));
  fa fa_u_csamul_cska32_fa21_30_out(.a(u_csamul_cska32_and21_30[0]), .b(u_csamul_cska32_fa22_29_xor1[0]), .cin(u_csamul_cska32_fa21_29_or0[0]), .fa_xor1(u_csamul_cska32_fa21_30_xor1), .fa_or0(u_csamul_cska32_fa21_30_or0));
  and_gate and_gate_u_csamul_cska32_and22_30(.a(a[22]), .b(b[30]), .out(u_csamul_cska32_and22_30));
  fa fa_u_csamul_cska32_fa22_30_out(.a(u_csamul_cska32_and22_30[0]), .b(u_csamul_cska32_fa23_29_xor1[0]), .cin(u_csamul_cska32_fa22_29_or0[0]), .fa_xor1(u_csamul_cska32_fa22_30_xor1), .fa_or0(u_csamul_cska32_fa22_30_or0));
  and_gate and_gate_u_csamul_cska32_and23_30(.a(a[23]), .b(b[30]), .out(u_csamul_cska32_and23_30));
  fa fa_u_csamul_cska32_fa23_30_out(.a(u_csamul_cska32_and23_30[0]), .b(u_csamul_cska32_fa24_29_xor1[0]), .cin(u_csamul_cska32_fa23_29_or0[0]), .fa_xor1(u_csamul_cska32_fa23_30_xor1), .fa_or0(u_csamul_cska32_fa23_30_or0));
  and_gate and_gate_u_csamul_cska32_and24_30(.a(a[24]), .b(b[30]), .out(u_csamul_cska32_and24_30));
  fa fa_u_csamul_cska32_fa24_30_out(.a(u_csamul_cska32_and24_30[0]), .b(u_csamul_cska32_fa25_29_xor1[0]), .cin(u_csamul_cska32_fa24_29_or0[0]), .fa_xor1(u_csamul_cska32_fa24_30_xor1), .fa_or0(u_csamul_cska32_fa24_30_or0));
  and_gate and_gate_u_csamul_cska32_and25_30(.a(a[25]), .b(b[30]), .out(u_csamul_cska32_and25_30));
  fa fa_u_csamul_cska32_fa25_30_out(.a(u_csamul_cska32_and25_30[0]), .b(u_csamul_cska32_fa26_29_xor1[0]), .cin(u_csamul_cska32_fa25_29_or0[0]), .fa_xor1(u_csamul_cska32_fa25_30_xor1), .fa_or0(u_csamul_cska32_fa25_30_or0));
  and_gate and_gate_u_csamul_cska32_and26_30(.a(a[26]), .b(b[30]), .out(u_csamul_cska32_and26_30));
  fa fa_u_csamul_cska32_fa26_30_out(.a(u_csamul_cska32_and26_30[0]), .b(u_csamul_cska32_fa27_29_xor1[0]), .cin(u_csamul_cska32_fa26_29_or0[0]), .fa_xor1(u_csamul_cska32_fa26_30_xor1), .fa_or0(u_csamul_cska32_fa26_30_or0));
  and_gate and_gate_u_csamul_cska32_and27_30(.a(a[27]), .b(b[30]), .out(u_csamul_cska32_and27_30));
  fa fa_u_csamul_cska32_fa27_30_out(.a(u_csamul_cska32_and27_30[0]), .b(u_csamul_cska32_fa28_29_xor1[0]), .cin(u_csamul_cska32_fa27_29_or0[0]), .fa_xor1(u_csamul_cska32_fa27_30_xor1), .fa_or0(u_csamul_cska32_fa27_30_or0));
  and_gate and_gate_u_csamul_cska32_and28_30(.a(a[28]), .b(b[30]), .out(u_csamul_cska32_and28_30));
  fa fa_u_csamul_cska32_fa28_30_out(.a(u_csamul_cska32_and28_30[0]), .b(u_csamul_cska32_fa29_29_xor1[0]), .cin(u_csamul_cska32_fa28_29_or0[0]), .fa_xor1(u_csamul_cska32_fa28_30_xor1), .fa_or0(u_csamul_cska32_fa28_30_or0));
  and_gate and_gate_u_csamul_cska32_and29_30(.a(a[29]), .b(b[30]), .out(u_csamul_cska32_and29_30));
  fa fa_u_csamul_cska32_fa29_30_out(.a(u_csamul_cska32_and29_30[0]), .b(u_csamul_cska32_fa30_29_xor1[0]), .cin(u_csamul_cska32_fa29_29_or0[0]), .fa_xor1(u_csamul_cska32_fa29_30_xor1), .fa_or0(u_csamul_cska32_fa29_30_or0));
  and_gate and_gate_u_csamul_cska32_and30_30(.a(a[30]), .b(b[30]), .out(u_csamul_cska32_and30_30));
  fa fa_u_csamul_cska32_fa30_30_out(.a(u_csamul_cska32_and30_30[0]), .b(u_csamul_cska32_and31_29[0]), .cin(u_csamul_cska32_fa30_29_or0[0]), .fa_xor1(u_csamul_cska32_fa30_30_xor1), .fa_or0(u_csamul_cska32_fa30_30_or0));
  and_gate and_gate_u_csamul_cska32_and31_30(.a(a[31]), .b(b[30]), .out(u_csamul_cska32_and31_30));
  and_gate and_gate_u_csamul_cska32_and0_31(.a(a[0]), .b(b[31]), .out(u_csamul_cska32_and0_31));
  fa fa_u_csamul_cska32_fa0_31_out(.a(u_csamul_cska32_and0_31[0]), .b(u_csamul_cska32_fa1_30_xor1[0]), .cin(u_csamul_cska32_fa0_30_or0[0]), .fa_xor1(u_csamul_cska32_fa0_31_xor1), .fa_or0(u_csamul_cska32_fa0_31_or0));
  and_gate and_gate_u_csamul_cska32_and1_31(.a(a[1]), .b(b[31]), .out(u_csamul_cska32_and1_31));
  fa fa_u_csamul_cska32_fa1_31_out(.a(u_csamul_cska32_and1_31[0]), .b(u_csamul_cska32_fa2_30_xor1[0]), .cin(u_csamul_cska32_fa1_30_or0[0]), .fa_xor1(u_csamul_cska32_fa1_31_xor1), .fa_or0(u_csamul_cska32_fa1_31_or0));
  and_gate and_gate_u_csamul_cska32_and2_31(.a(a[2]), .b(b[31]), .out(u_csamul_cska32_and2_31));
  fa fa_u_csamul_cska32_fa2_31_out(.a(u_csamul_cska32_and2_31[0]), .b(u_csamul_cska32_fa3_30_xor1[0]), .cin(u_csamul_cska32_fa2_30_or0[0]), .fa_xor1(u_csamul_cska32_fa2_31_xor1), .fa_or0(u_csamul_cska32_fa2_31_or0));
  and_gate and_gate_u_csamul_cska32_and3_31(.a(a[3]), .b(b[31]), .out(u_csamul_cska32_and3_31));
  fa fa_u_csamul_cska32_fa3_31_out(.a(u_csamul_cska32_and3_31[0]), .b(u_csamul_cska32_fa4_30_xor1[0]), .cin(u_csamul_cska32_fa3_30_or0[0]), .fa_xor1(u_csamul_cska32_fa3_31_xor1), .fa_or0(u_csamul_cska32_fa3_31_or0));
  and_gate and_gate_u_csamul_cska32_and4_31(.a(a[4]), .b(b[31]), .out(u_csamul_cska32_and4_31));
  fa fa_u_csamul_cska32_fa4_31_out(.a(u_csamul_cska32_and4_31[0]), .b(u_csamul_cska32_fa5_30_xor1[0]), .cin(u_csamul_cska32_fa4_30_or0[0]), .fa_xor1(u_csamul_cska32_fa4_31_xor1), .fa_or0(u_csamul_cska32_fa4_31_or0));
  and_gate and_gate_u_csamul_cska32_and5_31(.a(a[5]), .b(b[31]), .out(u_csamul_cska32_and5_31));
  fa fa_u_csamul_cska32_fa5_31_out(.a(u_csamul_cska32_and5_31[0]), .b(u_csamul_cska32_fa6_30_xor1[0]), .cin(u_csamul_cska32_fa5_30_or0[0]), .fa_xor1(u_csamul_cska32_fa5_31_xor1), .fa_or0(u_csamul_cska32_fa5_31_or0));
  and_gate and_gate_u_csamul_cska32_and6_31(.a(a[6]), .b(b[31]), .out(u_csamul_cska32_and6_31));
  fa fa_u_csamul_cska32_fa6_31_out(.a(u_csamul_cska32_and6_31[0]), .b(u_csamul_cska32_fa7_30_xor1[0]), .cin(u_csamul_cska32_fa6_30_or0[0]), .fa_xor1(u_csamul_cska32_fa6_31_xor1), .fa_or0(u_csamul_cska32_fa6_31_or0));
  and_gate and_gate_u_csamul_cska32_and7_31(.a(a[7]), .b(b[31]), .out(u_csamul_cska32_and7_31));
  fa fa_u_csamul_cska32_fa7_31_out(.a(u_csamul_cska32_and7_31[0]), .b(u_csamul_cska32_fa8_30_xor1[0]), .cin(u_csamul_cska32_fa7_30_or0[0]), .fa_xor1(u_csamul_cska32_fa7_31_xor1), .fa_or0(u_csamul_cska32_fa7_31_or0));
  and_gate and_gate_u_csamul_cska32_and8_31(.a(a[8]), .b(b[31]), .out(u_csamul_cska32_and8_31));
  fa fa_u_csamul_cska32_fa8_31_out(.a(u_csamul_cska32_and8_31[0]), .b(u_csamul_cska32_fa9_30_xor1[0]), .cin(u_csamul_cska32_fa8_30_or0[0]), .fa_xor1(u_csamul_cska32_fa8_31_xor1), .fa_or0(u_csamul_cska32_fa8_31_or0));
  and_gate and_gate_u_csamul_cska32_and9_31(.a(a[9]), .b(b[31]), .out(u_csamul_cska32_and9_31));
  fa fa_u_csamul_cska32_fa9_31_out(.a(u_csamul_cska32_and9_31[0]), .b(u_csamul_cska32_fa10_30_xor1[0]), .cin(u_csamul_cska32_fa9_30_or0[0]), .fa_xor1(u_csamul_cska32_fa9_31_xor1), .fa_or0(u_csamul_cska32_fa9_31_or0));
  and_gate and_gate_u_csamul_cska32_and10_31(.a(a[10]), .b(b[31]), .out(u_csamul_cska32_and10_31));
  fa fa_u_csamul_cska32_fa10_31_out(.a(u_csamul_cska32_and10_31[0]), .b(u_csamul_cska32_fa11_30_xor1[0]), .cin(u_csamul_cska32_fa10_30_or0[0]), .fa_xor1(u_csamul_cska32_fa10_31_xor1), .fa_or0(u_csamul_cska32_fa10_31_or0));
  and_gate and_gate_u_csamul_cska32_and11_31(.a(a[11]), .b(b[31]), .out(u_csamul_cska32_and11_31));
  fa fa_u_csamul_cska32_fa11_31_out(.a(u_csamul_cska32_and11_31[0]), .b(u_csamul_cska32_fa12_30_xor1[0]), .cin(u_csamul_cska32_fa11_30_or0[0]), .fa_xor1(u_csamul_cska32_fa11_31_xor1), .fa_or0(u_csamul_cska32_fa11_31_or0));
  and_gate and_gate_u_csamul_cska32_and12_31(.a(a[12]), .b(b[31]), .out(u_csamul_cska32_and12_31));
  fa fa_u_csamul_cska32_fa12_31_out(.a(u_csamul_cska32_and12_31[0]), .b(u_csamul_cska32_fa13_30_xor1[0]), .cin(u_csamul_cska32_fa12_30_or0[0]), .fa_xor1(u_csamul_cska32_fa12_31_xor1), .fa_or0(u_csamul_cska32_fa12_31_or0));
  and_gate and_gate_u_csamul_cska32_and13_31(.a(a[13]), .b(b[31]), .out(u_csamul_cska32_and13_31));
  fa fa_u_csamul_cska32_fa13_31_out(.a(u_csamul_cska32_and13_31[0]), .b(u_csamul_cska32_fa14_30_xor1[0]), .cin(u_csamul_cska32_fa13_30_or0[0]), .fa_xor1(u_csamul_cska32_fa13_31_xor1), .fa_or0(u_csamul_cska32_fa13_31_or0));
  and_gate and_gate_u_csamul_cska32_and14_31(.a(a[14]), .b(b[31]), .out(u_csamul_cska32_and14_31));
  fa fa_u_csamul_cska32_fa14_31_out(.a(u_csamul_cska32_and14_31[0]), .b(u_csamul_cska32_fa15_30_xor1[0]), .cin(u_csamul_cska32_fa14_30_or0[0]), .fa_xor1(u_csamul_cska32_fa14_31_xor1), .fa_or0(u_csamul_cska32_fa14_31_or0));
  and_gate and_gate_u_csamul_cska32_and15_31(.a(a[15]), .b(b[31]), .out(u_csamul_cska32_and15_31));
  fa fa_u_csamul_cska32_fa15_31_out(.a(u_csamul_cska32_and15_31[0]), .b(u_csamul_cska32_fa16_30_xor1[0]), .cin(u_csamul_cska32_fa15_30_or0[0]), .fa_xor1(u_csamul_cska32_fa15_31_xor1), .fa_or0(u_csamul_cska32_fa15_31_or0));
  and_gate and_gate_u_csamul_cska32_and16_31(.a(a[16]), .b(b[31]), .out(u_csamul_cska32_and16_31));
  fa fa_u_csamul_cska32_fa16_31_out(.a(u_csamul_cska32_and16_31[0]), .b(u_csamul_cska32_fa17_30_xor1[0]), .cin(u_csamul_cska32_fa16_30_or0[0]), .fa_xor1(u_csamul_cska32_fa16_31_xor1), .fa_or0(u_csamul_cska32_fa16_31_or0));
  and_gate and_gate_u_csamul_cska32_and17_31(.a(a[17]), .b(b[31]), .out(u_csamul_cska32_and17_31));
  fa fa_u_csamul_cska32_fa17_31_out(.a(u_csamul_cska32_and17_31[0]), .b(u_csamul_cska32_fa18_30_xor1[0]), .cin(u_csamul_cska32_fa17_30_or0[0]), .fa_xor1(u_csamul_cska32_fa17_31_xor1), .fa_or0(u_csamul_cska32_fa17_31_or0));
  and_gate and_gate_u_csamul_cska32_and18_31(.a(a[18]), .b(b[31]), .out(u_csamul_cska32_and18_31));
  fa fa_u_csamul_cska32_fa18_31_out(.a(u_csamul_cska32_and18_31[0]), .b(u_csamul_cska32_fa19_30_xor1[0]), .cin(u_csamul_cska32_fa18_30_or0[0]), .fa_xor1(u_csamul_cska32_fa18_31_xor1), .fa_or0(u_csamul_cska32_fa18_31_or0));
  and_gate and_gate_u_csamul_cska32_and19_31(.a(a[19]), .b(b[31]), .out(u_csamul_cska32_and19_31));
  fa fa_u_csamul_cska32_fa19_31_out(.a(u_csamul_cska32_and19_31[0]), .b(u_csamul_cska32_fa20_30_xor1[0]), .cin(u_csamul_cska32_fa19_30_or0[0]), .fa_xor1(u_csamul_cska32_fa19_31_xor1), .fa_or0(u_csamul_cska32_fa19_31_or0));
  and_gate and_gate_u_csamul_cska32_and20_31(.a(a[20]), .b(b[31]), .out(u_csamul_cska32_and20_31));
  fa fa_u_csamul_cska32_fa20_31_out(.a(u_csamul_cska32_and20_31[0]), .b(u_csamul_cska32_fa21_30_xor1[0]), .cin(u_csamul_cska32_fa20_30_or0[0]), .fa_xor1(u_csamul_cska32_fa20_31_xor1), .fa_or0(u_csamul_cska32_fa20_31_or0));
  and_gate and_gate_u_csamul_cska32_and21_31(.a(a[21]), .b(b[31]), .out(u_csamul_cska32_and21_31));
  fa fa_u_csamul_cska32_fa21_31_out(.a(u_csamul_cska32_and21_31[0]), .b(u_csamul_cska32_fa22_30_xor1[0]), .cin(u_csamul_cska32_fa21_30_or0[0]), .fa_xor1(u_csamul_cska32_fa21_31_xor1), .fa_or0(u_csamul_cska32_fa21_31_or0));
  and_gate and_gate_u_csamul_cska32_and22_31(.a(a[22]), .b(b[31]), .out(u_csamul_cska32_and22_31));
  fa fa_u_csamul_cska32_fa22_31_out(.a(u_csamul_cska32_and22_31[0]), .b(u_csamul_cska32_fa23_30_xor1[0]), .cin(u_csamul_cska32_fa22_30_or0[0]), .fa_xor1(u_csamul_cska32_fa22_31_xor1), .fa_or0(u_csamul_cska32_fa22_31_or0));
  and_gate and_gate_u_csamul_cska32_and23_31(.a(a[23]), .b(b[31]), .out(u_csamul_cska32_and23_31));
  fa fa_u_csamul_cska32_fa23_31_out(.a(u_csamul_cska32_and23_31[0]), .b(u_csamul_cska32_fa24_30_xor1[0]), .cin(u_csamul_cska32_fa23_30_or0[0]), .fa_xor1(u_csamul_cska32_fa23_31_xor1), .fa_or0(u_csamul_cska32_fa23_31_or0));
  and_gate and_gate_u_csamul_cska32_and24_31(.a(a[24]), .b(b[31]), .out(u_csamul_cska32_and24_31));
  fa fa_u_csamul_cska32_fa24_31_out(.a(u_csamul_cska32_and24_31[0]), .b(u_csamul_cska32_fa25_30_xor1[0]), .cin(u_csamul_cska32_fa24_30_or0[0]), .fa_xor1(u_csamul_cska32_fa24_31_xor1), .fa_or0(u_csamul_cska32_fa24_31_or0));
  and_gate and_gate_u_csamul_cska32_and25_31(.a(a[25]), .b(b[31]), .out(u_csamul_cska32_and25_31));
  fa fa_u_csamul_cska32_fa25_31_out(.a(u_csamul_cska32_and25_31[0]), .b(u_csamul_cska32_fa26_30_xor1[0]), .cin(u_csamul_cska32_fa25_30_or0[0]), .fa_xor1(u_csamul_cska32_fa25_31_xor1), .fa_or0(u_csamul_cska32_fa25_31_or0));
  and_gate and_gate_u_csamul_cska32_and26_31(.a(a[26]), .b(b[31]), .out(u_csamul_cska32_and26_31));
  fa fa_u_csamul_cska32_fa26_31_out(.a(u_csamul_cska32_and26_31[0]), .b(u_csamul_cska32_fa27_30_xor1[0]), .cin(u_csamul_cska32_fa26_30_or0[0]), .fa_xor1(u_csamul_cska32_fa26_31_xor1), .fa_or0(u_csamul_cska32_fa26_31_or0));
  and_gate and_gate_u_csamul_cska32_and27_31(.a(a[27]), .b(b[31]), .out(u_csamul_cska32_and27_31));
  fa fa_u_csamul_cska32_fa27_31_out(.a(u_csamul_cska32_and27_31[0]), .b(u_csamul_cska32_fa28_30_xor1[0]), .cin(u_csamul_cska32_fa27_30_or0[0]), .fa_xor1(u_csamul_cska32_fa27_31_xor1), .fa_or0(u_csamul_cska32_fa27_31_or0));
  and_gate and_gate_u_csamul_cska32_and28_31(.a(a[28]), .b(b[31]), .out(u_csamul_cska32_and28_31));
  fa fa_u_csamul_cska32_fa28_31_out(.a(u_csamul_cska32_and28_31[0]), .b(u_csamul_cska32_fa29_30_xor1[0]), .cin(u_csamul_cska32_fa28_30_or0[0]), .fa_xor1(u_csamul_cska32_fa28_31_xor1), .fa_or0(u_csamul_cska32_fa28_31_or0));
  and_gate and_gate_u_csamul_cska32_and29_31(.a(a[29]), .b(b[31]), .out(u_csamul_cska32_and29_31));
  fa fa_u_csamul_cska32_fa29_31_out(.a(u_csamul_cska32_and29_31[0]), .b(u_csamul_cska32_fa30_30_xor1[0]), .cin(u_csamul_cska32_fa29_30_or0[0]), .fa_xor1(u_csamul_cska32_fa29_31_xor1), .fa_or0(u_csamul_cska32_fa29_31_or0));
  and_gate and_gate_u_csamul_cska32_and30_31(.a(a[30]), .b(b[31]), .out(u_csamul_cska32_and30_31));
  fa fa_u_csamul_cska32_fa30_31_out(.a(u_csamul_cska32_and30_31[0]), .b(u_csamul_cska32_and31_30[0]), .cin(u_csamul_cska32_fa30_30_or0[0]), .fa_xor1(u_csamul_cska32_fa30_31_xor1), .fa_or0(u_csamul_cska32_fa30_31_or0));
  and_gate and_gate_u_csamul_cska32_and31_31(.a(a[31]), .b(b[31]), .out(u_csamul_cska32_and31_31));
  assign u_csamul_cska32_u_cska32_a[0] = u_csamul_cska32_fa1_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[1] = u_csamul_cska32_fa2_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[2] = u_csamul_cska32_fa3_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[3] = u_csamul_cska32_fa4_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[4] = u_csamul_cska32_fa5_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[5] = u_csamul_cska32_fa6_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[6] = u_csamul_cska32_fa7_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[7] = u_csamul_cska32_fa8_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[8] = u_csamul_cska32_fa9_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[9] = u_csamul_cska32_fa10_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[10] = u_csamul_cska32_fa11_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[11] = u_csamul_cska32_fa12_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[12] = u_csamul_cska32_fa13_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[13] = u_csamul_cska32_fa14_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[14] = u_csamul_cska32_fa15_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[15] = u_csamul_cska32_fa16_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[16] = u_csamul_cska32_fa17_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[17] = u_csamul_cska32_fa18_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[18] = u_csamul_cska32_fa19_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[19] = u_csamul_cska32_fa20_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[20] = u_csamul_cska32_fa21_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[21] = u_csamul_cska32_fa22_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[22] = u_csamul_cska32_fa23_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[23] = u_csamul_cska32_fa24_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[24] = u_csamul_cska32_fa25_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[25] = u_csamul_cska32_fa26_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[26] = u_csamul_cska32_fa27_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[27] = u_csamul_cska32_fa28_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[28] = u_csamul_cska32_fa29_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[29] = u_csamul_cska32_fa30_31_xor1[0];
  assign u_csamul_cska32_u_cska32_a[30] = u_csamul_cska32_and31_31[0];
  assign u_csamul_cska32_u_cska32_a[31] = 1'b0;
  assign u_csamul_cska32_u_cska32_b[0] = u_csamul_cska32_fa0_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[1] = u_csamul_cska32_fa1_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[2] = u_csamul_cska32_fa2_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[3] = u_csamul_cska32_fa3_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[4] = u_csamul_cska32_fa4_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[5] = u_csamul_cska32_fa5_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[6] = u_csamul_cska32_fa6_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[7] = u_csamul_cska32_fa7_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[8] = u_csamul_cska32_fa8_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[9] = u_csamul_cska32_fa9_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[10] = u_csamul_cska32_fa10_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[11] = u_csamul_cska32_fa11_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[12] = u_csamul_cska32_fa12_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[13] = u_csamul_cska32_fa13_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[14] = u_csamul_cska32_fa14_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[15] = u_csamul_cska32_fa15_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[16] = u_csamul_cska32_fa16_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[17] = u_csamul_cska32_fa17_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[18] = u_csamul_cska32_fa18_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[19] = u_csamul_cska32_fa19_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[20] = u_csamul_cska32_fa20_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[21] = u_csamul_cska32_fa21_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[22] = u_csamul_cska32_fa22_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[23] = u_csamul_cska32_fa23_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[24] = u_csamul_cska32_fa24_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[25] = u_csamul_cska32_fa25_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[26] = u_csamul_cska32_fa26_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[27] = u_csamul_cska32_fa27_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[28] = u_csamul_cska32_fa28_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[29] = u_csamul_cska32_fa29_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[30] = u_csamul_cska32_fa30_31_or0[0];
  assign u_csamul_cska32_u_cska32_b[31] = 1'b0;
  u_cska32 u_cska32_u_csamul_cska32_u_cska32_out(.a(u_csamul_cska32_u_cska32_a), .b(u_csamul_cska32_u_cska32_b), .u_cska32_out(u_csamul_cska32_u_cska32_out));

  assign u_csamul_cska32_out[0] = u_csamul_cska32_and0_0[0];
  assign u_csamul_cska32_out[1] = u_csamul_cska32_ha0_1_xor0[0];
  assign u_csamul_cska32_out[2] = u_csamul_cska32_fa0_2_xor1[0];
  assign u_csamul_cska32_out[3] = u_csamul_cska32_fa0_3_xor1[0];
  assign u_csamul_cska32_out[4] = u_csamul_cska32_fa0_4_xor1[0];
  assign u_csamul_cska32_out[5] = u_csamul_cska32_fa0_5_xor1[0];
  assign u_csamul_cska32_out[6] = u_csamul_cska32_fa0_6_xor1[0];
  assign u_csamul_cska32_out[7] = u_csamul_cska32_fa0_7_xor1[0];
  assign u_csamul_cska32_out[8] = u_csamul_cska32_fa0_8_xor1[0];
  assign u_csamul_cska32_out[9] = u_csamul_cska32_fa0_9_xor1[0];
  assign u_csamul_cska32_out[10] = u_csamul_cska32_fa0_10_xor1[0];
  assign u_csamul_cska32_out[11] = u_csamul_cska32_fa0_11_xor1[0];
  assign u_csamul_cska32_out[12] = u_csamul_cska32_fa0_12_xor1[0];
  assign u_csamul_cska32_out[13] = u_csamul_cska32_fa0_13_xor1[0];
  assign u_csamul_cska32_out[14] = u_csamul_cska32_fa0_14_xor1[0];
  assign u_csamul_cska32_out[15] = u_csamul_cska32_fa0_15_xor1[0];
  assign u_csamul_cska32_out[16] = u_csamul_cska32_fa0_16_xor1[0];
  assign u_csamul_cska32_out[17] = u_csamul_cska32_fa0_17_xor1[0];
  assign u_csamul_cska32_out[18] = u_csamul_cska32_fa0_18_xor1[0];
  assign u_csamul_cska32_out[19] = u_csamul_cska32_fa0_19_xor1[0];
  assign u_csamul_cska32_out[20] = u_csamul_cska32_fa0_20_xor1[0];
  assign u_csamul_cska32_out[21] = u_csamul_cska32_fa0_21_xor1[0];
  assign u_csamul_cska32_out[22] = u_csamul_cska32_fa0_22_xor1[0];
  assign u_csamul_cska32_out[23] = u_csamul_cska32_fa0_23_xor1[0];
  assign u_csamul_cska32_out[24] = u_csamul_cska32_fa0_24_xor1[0];
  assign u_csamul_cska32_out[25] = u_csamul_cska32_fa0_25_xor1[0];
  assign u_csamul_cska32_out[26] = u_csamul_cska32_fa0_26_xor1[0];
  assign u_csamul_cska32_out[27] = u_csamul_cska32_fa0_27_xor1[0];
  assign u_csamul_cska32_out[28] = u_csamul_cska32_fa0_28_xor1[0];
  assign u_csamul_cska32_out[29] = u_csamul_cska32_fa0_29_xor1[0];
  assign u_csamul_cska32_out[30] = u_csamul_cska32_fa0_30_xor1[0];
  assign u_csamul_cska32_out[31] = u_csamul_cska32_fa0_31_xor1[0];
  assign u_csamul_cska32_out[32] = u_csamul_cska32_u_cska32_out[0];
  assign u_csamul_cska32_out[33] = u_csamul_cska32_u_cska32_out[1];
  assign u_csamul_cska32_out[34] = u_csamul_cska32_u_cska32_out[2];
  assign u_csamul_cska32_out[35] = u_csamul_cska32_u_cska32_out[3];
  assign u_csamul_cska32_out[36] = u_csamul_cska32_u_cska32_out[4];
  assign u_csamul_cska32_out[37] = u_csamul_cska32_u_cska32_out[5];
  assign u_csamul_cska32_out[38] = u_csamul_cska32_u_cska32_out[6];
  assign u_csamul_cska32_out[39] = u_csamul_cska32_u_cska32_out[7];
  assign u_csamul_cska32_out[40] = u_csamul_cska32_u_cska32_out[8];
  assign u_csamul_cska32_out[41] = u_csamul_cska32_u_cska32_out[9];
  assign u_csamul_cska32_out[42] = u_csamul_cska32_u_cska32_out[10];
  assign u_csamul_cska32_out[43] = u_csamul_cska32_u_cska32_out[11];
  assign u_csamul_cska32_out[44] = u_csamul_cska32_u_cska32_out[12];
  assign u_csamul_cska32_out[45] = u_csamul_cska32_u_cska32_out[13];
  assign u_csamul_cska32_out[46] = u_csamul_cska32_u_cska32_out[14];
  assign u_csamul_cska32_out[47] = u_csamul_cska32_u_cska32_out[15];
  assign u_csamul_cska32_out[48] = u_csamul_cska32_u_cska32_out[16];
  assign u_csamul_cska32_out[49] = u_csamul_cska32_u_cska32_out[17];
  assign u_csamul_cska32_out[50] = u_csamul_cska32_u_cska32_out[18];
  assign u_csamul_cska32_out[51] = u_csamul_cska32_u_cska32_out[19];
  assign u_csamul_cska32_out[52] = u_csamul_cska32_u_cska32_out[20];
  assign u_csamul_cska32_out[53] = u_csamul_cska32_u_cska32_out[21];
  assign u_csamul_cska32_out[54] = u_csamul_cska32_u_cska32_out[22];
  assign u_csamul_cska32_out[55] = u_csamul_cska32_u_cska32_out[23];
  assign u_csamul_cska32_out[56] = u_csamul_cska32_u_cska32_out[24];
  assign u_csamul_cska32_out[57] = u_csamul_cska32_u_cska32_out[25];
  assign u_csamul_cska32_out[58] = u_csamul_cska32_u_cska32_out[26];
  assign u_csamul_cska32_out[59] = u_csamul_cska32_u_cska32_out[27];
  assign u_csamul_cska32_out[60] = u_csamul_cska32_u_cska32_out[28];
  assign u_csamul_cska32_out[61] = u_csamul_cska32_u_cska32_out[29];
  assign u_csamul_cska32_out[62] = u_csamul_cska32_u_cska32_out[30];
  assign u_csamul_cska32_out[63] = u_csamul_cska32_u_cska32_out[31];
endmodule