module u_CSAwallace_pg_rca12(input [11:0] a, input [11:0] b, output [23:0] u_CSAwallace_pg_rca12_out);
  wire u_CSAwallace_pg_rca12_and_0_0;
  wire u_CSAwallace_pg_rca12_and_1_0;
  wire u_CSAwallace_pg_rca12_and_2_0;
  wire u_CSAwallace_pg_rca12_and_3_0;
  wire u_CSAwallace_pg_rca12_and_4_0;
  wire u_CSAwallace_pg_rca12_and_5_0;
  wire u_CSAwallace_pg_rca12_and_6_0;
  wire u_CSAwallace_pg_rca12_and_7_0;
  wire u_CSAwallace_pg_rca12_and_8_0;
  wire u_CSAwallace_pg_rca12_and_9_0;
  wire u_CSAwallace_pg_rca12_and_10_0;
  wire u_CSAwallace_pg_rca12_and_11_0;
  wire u_CSAwallace_pg_rca12_and_0_1;
  wire u_CSAwallace_pg_rca12_and_1_1;
  wire u_CSAwallace_pg_rca12_and_2_1;
  wire u_CSAwallace_pg_rca12_and_3_1;
  wire u_CSAwallace_pg_rca12_and_4_1;
  wire u_CSAwallace_pg_rca12_and_5_1;
  wire u_CSAwallace_pg_rca12_and_6_1;
  wire u_CSAwallace_pg_rca12_and_7_1;
  wire u_CSAwallace_pg_rca12_and_8_1;
  wire u_CSAwallace_pg_rca12_and_9_1;
  wire u_CSAwallace_pg_rca12_and_10_1;
  wire u_CSAwallace_pg_rca12_and_11_1;
  wire u_CSAwallace_pg_rca12_and_0_2;
  wire u_CSAwallace_pg_rca12_and_1_2;
  wire u_CSAwallace_pg_rca12_and_2_2;
  wire u_CSAwallace_pg_rca12_and_3_2;
  wire u_CSAwallace_pg_rca12_and_4_2;
  wire u_CSAwallace_pg_rca12_and_5_2;
  wire u_CSAwallace_pg_rca12_and_6_2;
  wire u_CSAwallace_pg_rca12_and_7_2;
  wire u_CSAwallace_pg_rca12_and_8_2;
  wire u_CSAwallace_pg_rca12_and_9_2;
  wire u_CSAwallace_pg_rca12_and_10_2;
  wire u_CSAwallace_pg_rca12_and_11_2;
  wire u_CSAwallace_pg_rca12_and_0_3;
  wire u_CSAwallace_pg_rca12_and_1_3;
  wire u_CSAwallace_pg_rca12_and_2_3;
  wire u_CSAwallace_pg_rca12_and_3_3;
  wire u_CSAwallace_pg_rca12_and_4_3;
  wire u_CSAwallace_pg_rca12_and_5_3;
  wire u_CSAwallace_pg_rca12_and_6_3;
  wire u_CSAwallace_pg_rca12_and_7_3;
  wire u_CSAwallace_pg_rca12_and_8_3;
  wire u_CSAwallace_pg_rca12_and_9_3;
  wire u_CSAwallace_pg_rca12_and_10_3;
  wire u_CSAwallace_pg_rca12_and_11_3;
  wire u_CSAwallace_pg_rca12_and_0_4;
  wire u_CSAwallace_pg_rca12_and_1_4;
  wire u_CSAwallace_pg_rca12_and_2_4;
  wire u_CSAwallace_pg_rca12_and_3_4;
  wire u_CSAwallace_pg_rca12_and_4_4;
  wire u_CSAwallace_pg_rca12_and_5_4;
  wire u_CSAwallace_pg_rca12_and_6_4;
  wire u_CSAwallace_pg_rca12_and_7_4;
  wire u_CSAwallace_pg_rca12_and_8_4;
  wire u_CSAwallace_pg_rca12_and_9_4;
  wire u_CSAwallace_pg_rca12_and_10_4;
  wire u_CSAwallace_pg_rca12_and_11_4;
  wire u_CSAwallace_pg_rca12_and_0_5;
  wire u_CSAwallace_pg_rca12_and_1_5;
  wire u_CSAwallace_pg_rca12_and_2_5;
  wire u_CSAwallace_pg_rca12_and_3_5;
  wire u_CSAwallace_pg_rca12_and_4_5;
  wire u_CSAwallace_pg_rca12_and_5_5;
  wire u_CSAwallace_pg_rca12_and_6_5;
  wire u_CSAwallace_pg_rca12_and_7_5;
  wire u_CSAwallace_pg_rca12_and_8_5;
  wire u_CSAwallace_pg_rca12_and_9_5;
  wire u_CSAwallace_pg_rca12_and_10_5;
  wire u_CSAwallace_pg_rca12_and_11_5;
  wire u_CSAwallace_pg_rca12_and_0_6;
  wire u_CSAwallace_pg_rca12_and_1_6;
  wire u_CSAwallace_pg_rca12_and_2_6;
  wire u_CSAwallace_pg_rca12_and_3_6;
  wire u_CSAwallace_pg_rca12_and_4_6;
  wire u_CSAwallace_pg_rca12_and_5_6;
  wire u_CSAwallace_pg_rca12_and_6_6;
  wire u_CSAwallace_pg_rca12_and_7_6;
  wire u_CSAwallace_pg_rca12_and_8_6;
  wire u_CSAwallace_pg_rca12_and_9_6;
  wire u_CSAwallace_pg_rca12_and_10_6;
  wire u_CSAwallace_pg_rca12_and_11_6;
  wire u_CSAwallace_pg_rca12_and_0_7;
  wire u_CSAwallace_pg_rca12_and_1_7;
  wire u_CSAwallace_pg_rca12_and_2_7;
  wire u_CSAwallace_pg_rca12_and_3_7;
  wire u_CSAwallace_pg_rca12_and_4_7;
  wire u_CSAwallace_pg_rca12_and_5_7;
  wire u_CSAwallace_pg_rca12_and_6_7;
  wire u_CSAwallace_pg_rca12_and_7_7;
  wire u_CSAwallace_pg_rca12_and_8_7;
  wire u_CSAwallace_pg_rca12_and_9_7;
  wire u_CSAwallace_pg_rca12_and_10_7;
  wire u_CSAwallace_pg_rca12_and_11_7;
  wire u_CSAwallace_pg_rca12_and_0_8;
  wire u_CSAwallace_pg_rca12_and_1_8;
  wire u_CSAwallace_pg_rca12_and_2_8;
  wire u_CSAwallace_pg_rca12_and_3_8;
  wire u_CSAwallace_pg_rca12_and_4_8;
  wire u_CSAwallace_pg_rca12_and_5_8;
  wire u_CSAwallace_pg_rca12_and_6_8;
  wire u_CSAwallace_pg_rca12_and_7_8;
  wire u_CSAwallace_pg_rca12_and_8_8;
  wire u_CSAwallace_pg_rca12_and_9_8;
  wire u_CSAwallace_pg_rca12_and_10_8;
  wire u_CSAwallace_pg_rca12_and_11_8;
  wire u_CSAwallace_pg_rca12_and_0_9;
  wire u_CSAwallace_pg_rca12_and_1_9;
  wire u_CSAwallace_pg_rca12_and_2_9;
  wire u_CSAwallace_pg_rca12_and_3_9;
  wire u_CSAwallace_pg_rca12_and_4_9;
  wire u_CSAwallace_pg_rca12_and_5_9;
  wire u_CSAwallace_pg_rca12_and_6_9;
  wire u_CSAwallace_pg_rca12_and_7_9;
  wire u_CSAwallace_pg_rca12_and_8_9;
  wire u_CSAwallace_pg_rca12_and_9_9;
  wire u_CSAwallace_pg_rca12_and_10_9;
  wire u_CSAwallace_pg_rca12_and_11_9;
  wire u_CSAwallace_pg_rca12_and_0_10;
  wire u_CSAwallace_pg_rca12_and_1_10;
  wire u_CSAwallace_pg_rca12_and_2_10;
  wire u_CSAwallace_pg_rca12_and_3_10;
  wire u_CSAwallace_pg_rca12_and_4_10;
  wire u_CSAwallace_pg_rca12_and_5_10;
  wire u_CSAwallace_pg_rca12_and_6_10;
  wire u_CSAwallace_pg_rca12_and_7_10;
  wire u_CSAwallace_pg_rca12_and_8_10;
  wire u_CSAwallace_pg_rca12_and_9_10;
  wire u_CSAwallace_pg_rca12_and_10_10;
  wire u_CSAwallace_pg_rca12_and_11_10;
  wire u_CSAwallace_pg_rca12_and_0_11;
  wire u_CSAwallace_pg_rca12_and_1_11;
  wire u_CSAwallace_pg_rca12_and_2_11;
  wire u_CSAwallace_pg_rca12_and_3_11;
  wire u_CSAwallace_pg_rca12_and_4_11;
  wire u_CSAwallace_pg_rca12_and_5_11;
  wire u_CSAwallace_pg_rca12_and_6_11;
  wire u_CSAwallace_pg_rca12_and_7_11;
  wire u_CSAwallace_pg_rca12_and_8_11;
  wire u_CSAwallace_pg_rca12_and_9_11;
  wire u_CSAwallace_pg_rca12_and_10_11;
  wire u_CSAwallace_pg_rca12_and_11_11;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa1_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa1_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa2_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa2_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa2_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa2_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa2_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa3_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa3_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa3_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa3_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa3_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa4_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa4_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa4_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa4_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa4_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa5_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa5_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa5_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa5_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa5_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa6_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa6_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa6_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa6_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa6_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa7_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa7_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa7_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa7_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa7_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa8_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa8_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa8_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa8_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa8_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa9_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa9_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa9_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa9_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa9_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa10_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa10_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa10_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa0_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa4_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa4_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa5_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa5_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa5_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa5_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa5_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa6_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa6_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa6_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa6_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa6_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa7_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa7_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa7_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa7_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa7_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa8_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa8_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa8_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa8_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa8_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa9_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa9_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa9_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa9_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa9_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa10_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa10_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa10_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa12_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa12_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa12_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa13_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa13_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa13_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa13_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa13_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa14_xor0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa14_and0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa14_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa14_and1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa14_or0;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa15_xor1;
  wire u_CSAwallace_pg_rca12_csa1_csa_component_fa15_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa7_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa7_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa8_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa8_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa8_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa8_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa8_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa9_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa9_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa9_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa9_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa9_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa10_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa10_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa10_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa12_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa12_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa12_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa13_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa13_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa13_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa13_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa13_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa14_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa14_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa14_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa14_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa14_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa15_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa15_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa15_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa15_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa15_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa16_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa16_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa16_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa16_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa16_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa17_xor0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa17_and0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa17_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa17_and1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa17_or0;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa18_xor1;
  wire u_CSAwallace_pg_rca12_csa2_csa_component_fa18_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa12_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa12_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa12_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa13_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa13_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa13_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa13_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa13_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa14_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa14_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa14_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa14_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa14_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa15_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa15_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa15_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa15_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa15_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa16_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa16_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa16_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa16_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa16_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa17_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa17_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa17_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa17_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa17_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa18_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa18_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa18_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa18_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa18_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa19_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa19_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa19_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa19_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa19_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa20_xor0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa20_and0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa20_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa20_and1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa20_or0;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa21_xor1;
  wire u_CSAwallace_pg_rca12_csa3_csa_component_fa21_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa2_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa2_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa3_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa3_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa3_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa3_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa3_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa4_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa4_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa4_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa4_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa4_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa5_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa5_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa5_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa5_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa5_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa6_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa6_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa6_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa6_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa6_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa7_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa7_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa7_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa7_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa7_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa8_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa8_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa8_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa8_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa8_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa9_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa9_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa9_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa9_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa9_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa10_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa10_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa10_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa12_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa12_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa12_or0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa13_xor0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa13_and0;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa13_xor1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa13_and1;
  wire u_CSAwallace_pg_rca12_csa4_csa_component_fa13_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa6_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa6_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa7_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa7_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa8_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa8_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa8_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa8_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa8_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa9_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa9_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa9_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa9_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa9_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa10_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa10_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa10_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa12_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa12_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa12_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa13_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa13_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa13_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa13_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa13_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa14_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa14_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa14_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa14_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa14_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa15_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa15_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa15_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa15_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa15_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa16_xor0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa16_and0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa16_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa16_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa16_or0;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa17_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa17_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa18_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa18_and1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa19_xor1;
  wire u_CSAwallace_pg_rca12_csa5_csa_component_fa19_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa3_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa3_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa4_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa4_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa5_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa5_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa5_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa5_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa5_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa6_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa6_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa6_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa6_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa6_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa7_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa7_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa7_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa7_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa7_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa8_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa8_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa8_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa8_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa8_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa9_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa9_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa9_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa9_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa9_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa10_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa10_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa10_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa12_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa12_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa12_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa13_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa13_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa13_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa13_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa13_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa14_xor0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa14_and0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa14_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa14_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa14_or0;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa15_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa15_and1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa16_xor1;
  wire u_CSAwallace_pg_rca12_csa6_csa_component_fa16_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa9_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa9_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa12_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa12_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa12_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa13_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa13_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa13_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa13_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa13_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa14_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa14_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa14_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa14_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa14_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa15_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa15_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa15_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa15_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa15_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa16_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa16_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa16_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa16_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa16_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa17_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa17_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa17_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa17_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa17_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa18_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa18_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa18_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa18_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa18_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa19_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa19_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa19_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa19_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa19_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa20_xor0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa20_and0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa20_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa20_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa20_or0;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa21_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa21_and1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa22_xor1;
  wire u_CSAwallace_pg_rca12_csa7_csa_component_fa22_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa4_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa4_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa5_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa5_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa6_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa6_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa7_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa7_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa7_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa7_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa7_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa8_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa8_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa8_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa8_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa8_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa9_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa9_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa9_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa9_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa9_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa10_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa10_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa10_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa12_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa12_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa12_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa13_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa13_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa13_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa13_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa13_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa14_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa14_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa14_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa14_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa14_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa15_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa15_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa15_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa15_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa15_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa16_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa16_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa16_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa16_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa16_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa17_xor0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa17_and0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa17_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa17_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa17_or0;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa18_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa18_and1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa19_xor1;
  wire u_CSAwallace_pg_rca12_csa8_csa_component_fa19_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa5_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa5_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa6_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa6_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa7_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa7_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa8_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa8_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa9_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa9_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa10_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa10_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa10_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa10_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa10_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa11_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa11_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa11_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa11_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa11_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa12_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa12_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa12_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa12_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa12_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa13_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa13_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa13_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa13_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa13_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa14_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa14_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa14_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa14_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa14_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa15_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa15_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa15_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa15_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa15_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa16_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa16_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa16_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa16_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa16_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa17_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa17_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa17_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa17_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa17_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa18_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa18_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa18_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa18_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa18_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa19_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa19_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa19_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa19_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa19_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa20_xor0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa20_and0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa20_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa20_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa20_or0;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa21_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa21_and1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa22_xor1;
  wire u_CSAwallace_pg_rca12_csa9_csa_component_fa22_and1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa6_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa6_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and7;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or7;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and8;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or8;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and9;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or9;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and10;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or10;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and11;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or11;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and12;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or12;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and13;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or13;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and14;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or14;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and15;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or15;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and16;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or16;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and17;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or17;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and18;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or18;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and19;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or19;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and20;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or20;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and21;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or21;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and22;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or22;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_xor0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_and0;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_xor1;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_and23;
  wire u_CSAwallace_pg_rca12_u_pg_rca24_or23;

  assign u_CSAwallace_pg_rca12_and_0_0 = a[0] & b[0];
  assign u_CSAwallace_pg_rca12_and_1_0 = a[1] & b[0];
  assign u_CSAwallace_pg_rca12_and_2_0 = a[2] & b[0];
  assign u_CSAwallace_pg_rca12_and_3_0 = a[3] & b[0];
  assign u_CSAwallace_pg_rca12_and_4_0 = a[4] & b[0];
  assign u_CSAwallace_pg_rca12_and_5_0 = a[5] & b[0];
  assign u_CSAwallace_pg_rca12_and_6_0 = a[6] & b[0];
  assign u_CSAwallace_pg_rca12_and_7_0 = a[7] & b[0];
  assign u_CSAwallace_pg_rca12_and_8_0 = a[8] & b[0];
  assign u_CSAwallace_pg_rca12_and_9_0 = a[9] & b[0];
  assign u_CSAwallace_pg_rca12_and_10_0 = a[10] & b[0];
  assign u_CSAwallace_pg_rca12_and_11_0 = a[11] & b[0];
  assign u_CSAwallace_pg_rca12_and_0_1 = a[0] & b[1];
  assign u_CSAwallace_pg_rca12_and_1_1 = a[1] & b[1];
  assign u_CSAwallace_pg_rca12_and_2_1 = a[2] & b[1];
  assign u_CSAwallace_pg_rca12_and_3_1 = a[3] & b[1];
  assign u_CSAwallace_pg_rca12_and_4_1 = a[4] & b[1];
  assign u_CSAwallace_pg_rca12_and_5_1 = a[5] & b[1];
  assign u_CSAwallace_pg_rca12_and_6_1 = a[6] & b[1];
  assign u_CSAwallace_pg_rca12_and_7_1 = a[7] & b[1];
  assign u_CSAwallace_pg_rca12_and_8_1 = a[8] & b[1];
  assign u_CSAwallace_pg_rca12_and_9_1 = a[9] & b[1];
  assign u_CSAwallace_pg_rca12_and_10_1 = a[10] & b[1];
  assign u_CSAwallace_pg_rca12_and_11_1 = a[11] & b[1];
  assign u_CSAwallace_pg_rca12_and_0_2 = a[0] & b[2];
  assign u_CSAwallace_pg_rca12_and_1_2 = a[1] & b[2];
  assign u_CSAwallace_pg_rca12_and_2_2 = a[2] & b[2];
  assign u_CSAwallace_pg_rca12_and_3_2 = a[3] & b[2];
  assign u_CSAwallace_pg_rca12_and_4_2 = a[4] & b[2];
  assign u_CSAwallace_pg_rca12_and_5_2 = a[5] & b[2];
  assign u_CSAwallace_pg_rca12_and_6_2 = a[6] & b[2];
  assign u_CSAwallace_pg_rca12_and_7_2 = a[7] & b[2];
  assign u_CSAwallace_pg_rca12_and_8_2 = a[8] & b[2];
  assign u_CSAwallace_pg_rca12_and_9_2 = a[9] & b[2];
  assign u_CSAwallace_pg_rca12_and_10_2 = a[10] & b[2];
  assign u_CSAwallace_pg_rca12_and_11_2 = a[11] & b[2];
  assign u_CSAwallace_pg_rca12_and_0_3 = a[0] & b[3];
  assign u_CSAwallace_pg_rca12_and_1_3 = a[1] & b[3];
  assign u_CSAwallace_pg_rca12_and_2_3 = a[2] & b[3];
  assign u_CSAwallace_pg_rca12_and_3_3 = a[3] & b[3];
  assign u_CSAwallace_pg_rca12_and_4_3 = a[4] & b[3];
  assign u_CSAwallace_pg_rca12_and_5_3 = a[5] & b[3];
  assign u_CSAwallace_pg_rca12_and_6_3 = a[6] & b[3];
  assign u_CSAwallace_pg_rca12_and_7_3 = a[7] & b[3];
  assign u_CSAwallace_pg_rca12_and_8_3 = a[8] & b[3];
  assign u_CSAwallace_pg_rca12_and_9_3 = a[9] & b[3];
  assign u_CSAwallace_pg_rca12_and_10_3 = a[10] & b[3];
  assign u_CSAwallace_pg_rca12_and_11_3 = a[11] & b[3];
  assign u_CSAwallace_pg_rca12_and_0_4 = a[0] & b[4];
  assign u_CSAwallace_pg_rca12_and_1_4 = a[1] & b[4];
  assign u_CSAwallace_pg_rca12_and_2_4 = a[2] & b[4];
  assign u_CSAwallace_pg_rca12_and_3_4 = a[3] & b[4];
  assign u_CSAwallace_pg_rca12_and_4_4 = a[4] & b[4];
  assign u_CSAwallace_pg_rca12_and_5_4 = a[5] & b[4];
  assign u_CSAwallace_pg_rca12_and_6_4 = a[6] & b[4];
  assign u_CSAwallace_pg_rca12_and_7_4 = a[7] & b[4];
  assign u_CSAwallace_pg_rca12_and_8_4 = a[8] & b[4];
  assign u_CSAwallace_pg_rca12_and_9_4 = a[9] & b[4];
  assign u_CSAwallace_pg_rca12_and_10_4 = a[10] & b[4];
  assign u_CSAwallace_pg_rca12_and_11_4 = a[11] & b[4];
  assign u_CSAwallace_pg_rca12_and_0_5 = a[0] & b[5];
  assign u_CSAwallace_pg_rca12_and_1_5 = a[1] & b[5];
  assign u_CSAwallace_pg_rca12_and_2_5 = a[2] & b[5];
  assign u_CSAwallace_pg_rca12_and_3_5 = a[3] & b[5];
  assign u_CSAwallace_pg_rca12_and_4_5 = a[4] & b[5];
  assign u_CSAwallace_pg_rca12_and_5_5 = a[5] & b[5];
  assign u_CSAwallace_pg_rca12_and_6_5 = a[6] & b[5];
  assign u_CSAwallace_pg_rca12_and_7_5 = a[7] & b[5];
  assign u_CSAwallace_pg_rca12_and_8_5 = a[8] & b[5];
  assign u_CSAwallace_pg_rca12_and_9_5 = a[9] & b[5];
  assign u_CSAwallace_pg_rca12_and_10_5 = a[10] & b[5];
  assign u_CSAwallace_pg_rca12_and_11_5 = a[11] & b[5];
  assign u_CSAwallace_pg_rca12_and_0_6 = a[0] & b[6];
  assign u_CSAwallace_pg_rca12_and_1_6 = a[1] & b[6];
  assign u_CSAwallace_pg_rca12_and_2_6 = a[2] & b[6];
  assign u_CSAwallace_pg_rca12_and_3_6 = a[3] & b[6];
  assign u_CSAwallace_pg_rca12_and_4_6 = a[4] & b[6];
  assign u_CSAwallace_pg_rca12_and_5_6 = a[5] & b[6];
  assign u_CSAwallace_pg_rca12_and_6_6 = a[6] & b[6];
  assign u_CSAwallace_pg_rca12_and_7_6 = a[7] & b[6];
  assign u_CSAwallace_pg_rca12_and_8_6 = a[8] & b[6];
  assign u_CSAwallace_pg_rca12_and_9_6 = a[9] & b[6];
  assign u_CSAwallace_pg_rca12_and_10_6 = a[10] & b[6];
  assign u_CSAwallace_pg_rca12_and_11_6 = a[11] & b[6];
  assign u_CSAwallace_pg_rca12_and_0_7 = a[0] & b[7];
  assign u_CSAwallace_pg_rca12_and_1_7 = a[1] & b[7];
  assign u_CSAwallace_pg_rca12_and_2_7 = a[2] & b[7];
  assign u_CSAwallace_pg_rca12_and_3_7 = a[3] & b[7];
  assign u_CSAwallace_pg_rca12_and_4_7 = a[4] & b[7];
  assign u_CSAwallace_pg_rca12_and_5_7 = a[5] & b[7];
  assign u_CSAwallace_pg_rca12_and_6_7 = a[6] & b[7];
  assign u_CSAwallace_pg_rca12_and_7_7 = a[7] & b[7];
  assign u_CSAwallace_pg_rca12_and_8_7 = a[8] & b[7];
  assign u_CSAwallace_pg_rca12_and_9_7 = a[9] & b[7];
  assign u_CSAwallace_pg_rca12_and_10_7 = a[10] & b[7];
  assign u_CSAwallace_pg_rca12_and_11_7 = a[11] & b[7];
  assign u_CSAwallace_pg_rca12_and_0_8 = a[0] & b[8];
  assign u_CSAwallace_pg_rca12_and_1_8 = a[1] & b[8];
  assign u_CSAwallace_pg_rca12_and_2_8 = a[2] & b[8];
  assign u_CSAwallace_pg_rca12_and_3_8 = a[3] & b[8];
  assign u_CSAwallace_pg_rca12_and_4_8 = a[4] & b[8];
  assign u_CSAwallace_pg_rca12_and_5_8 = a[5] & b[8];
  assign u_CSAwallace_pg_rca12_and_6_8 = a[6] & b[8];
  assign u_CSAwallace_pg_rca12_and_7_8 = a[7] & b[8];
  assign u_CSAwallace_pg_rca12_and_8_8 = a[8] & b[8];
  assign u_CSAwallace_pg_rca12_and_9_8 = a[9] & b[8];
  assign u_CSAwallace_pg_rca12_and_10_8 = a[10] & b[8];
  assign u_CSAwallace_pg_rca12_and_11_8 = a[11] & b[8];
  assign u_CSAwallace_pg_rca12_and_0_9 = a[0] & b[9];
  assign u_CSAwallace_pg_rca12_and_1_9 = a[1] & b[9];
  assign u_CSAwallace_pg_rca12_and_2_9 = a[2] & b[9];
  assign u_CSAwallace_pg_rca12_and_3_9 = a[3] & b[9];
  assign u_CSAwallace_pg_rca12_and_4_9 = a[4] & b[9];
  assign u_CSAwallace_pg_rca12_and_5_9 = a[5] & b[9];
  assign u_CSAwallace_pg_rca12_and_6_9 = a[6] & b[9];
  assign u_CSAwallace_pg_rca12_and_7_9 = a[7] & b[9];
  assign u_CSAwallace_pg_rca12_and_8_9 = a[8] & b[9];
  assign u_CSAwallace_pg_rca12_and_9_9 = a[9] & b[9];
  assign u_CSAwallace_pg_rca12_and_10_9 = a[10] & b[9];
  assign u_CSAwallace_pg_rca12_and_11_9 = a[11] & b[9];
  assign u_CSAwallace_pg_rca12_and_0_10 = a[0] & b[10];
  assign u_CSAwallace_pg_rca12_and_1_10 = a[1] & b[10];
  assign u_CSAwallace_pg_rca12_and_2_10 = a[2] & b[10];
  assign u_CSAwallace_pg_rca12_and_3_10 = a[3] & b[10];
  assign u_CSAwallace_pg_rca12_and_4_10 = a[4] & b[10];
  assign u_CSAwallace_pg_rca12_and_5_10 = a[5] & b[10];
  assign u_CSAwallace_pg_rca12_and_6_10 = a[6] & b[10];
  assign u_CSAwallace_pg_rca12_and_7_10 = a[7] & b[10];
  assign u_CSAwallace_pg_rca12_and_8_10 = a[8] & b[10];
  assign u_CSAwallace_pg_rca12_and_9_10 = a[9] & b[10];
  assign u_CSAwallace_pg_rca12_and_10_10 = a[10] & b[10];
  assign u_CSAwallace_pg_rca12_and_11_10 = a[11] & b[10];
  assign u_CSAwallace_pg_rca12_and_0_11 = a[0] & b[11];
  assign u_CSAwallace_pg_rca12_and_1_11 = a[1] & b[11];
  assign u_CSAwallace_pg_rca12_and_2_11 = a[2] & b[11];
  assign u_CSAwallace_pg_rca12_and_3_11 = a[3] & b[11];
  assign u_CSAwallace_pg_rca12_and_4_11 = a[4] & b[11];
  assign u_CSAwallace_pg_rca12_and_5_11 = a[5] & b[11];
  assign u_CSAwallace_pg_rca12_and_6_11 = a[6] & b[11];
  assign u_CSAwallace_pg_rca12_and_7_11 = a[7] & b[11];
  assign u_CSAwallace_pg_rca12_and_8_11 = a[8] & b[11];
  assign u_CSAwallace_pg_rca12_and_9_11 = a[9] & b[11];
  assign u_CSAwallace_pg_rca12_and_10_11 = a[10] & b[11];
  assign u_CSAwallace_pg_rca12_and_11_11 = a[11] & b[11];
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa1_xor0 = u_CSAwallace_pg_rca12_and_1_0 ^ u_CSAwallace_pg_rca12_and_0_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa1_and0 = u_CSAwallace_pg_rca12_and_1_0 & u_CSAwallace_pg_rca12_and_0_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa2_xor0 = u_CSAwallace_pg_rca12_and_2_0 ^ u_CSAwallace_pg_rca12_and_1_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa2_and0 = u_CSAwallace_pg_rca12_and_2_0 & u_CSAwallace_pg_rca12_and_1_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa2_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa2_xor0 ^ u_CSAwallace_pg_rca12_and_0_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa2_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa2_xor0 & u_CSAwallace_pg_rca12_and_0_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa2_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa2_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa2_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa3_xor0 = u_CSAwallace_pg_rca12_and_3_0 ^ u_CSAwallace_pg_rca12_and_2_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa3_and0 = u_CSAwallace_pg_rca12_and_3_0 & u_CSAwallace_pg_rca12_and_2_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa3_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa3_xor0 ^ u_CSAwallace_pg_rca12_and_1_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa3_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa3_xor0 & u_CSAwallace_pg_rca12_and_1_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa3_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa3_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa3_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa4_xor0 = u_CSAwallace_pg_rca12_and_4_0 ^ u_CSAwallace_pg_rca12_and_3_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa4_and0 = u_CSAwallace_pg_rca12_and_4_0 & u_CSAwallace_pg_rca12_and_3_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa4_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa4_xor0 ^ u_CSAwallace_pg_rca12_and_2_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa4_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa4_xor0 & u_CSAwallace_pg_rca12_and_2_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa4_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa4_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa4_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa5_xor0 = u_CSAwallace_pg_rca12_and_5_0 ^ u_CSAwallace_pg_rca12_and_4_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa5_and0 = u_CSAwallace_pg_rca12_and_5_0 & u_CSAwallace_pg_rca12_and_4_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa5_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa5_xor0 ^ u_CSAwallace_pg_rca12_and_3_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa5_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa5_xor0 & u_CSAwallace_pg_rca12_and_3_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa5_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa5_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa5_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa6_xor0 = u_CSAwallace_pg_rca12_and_6_0 ^ u_CSAwallace_pg_rca12_and_5_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa6_and0 = u_CSAwallace_pg_rca12_and_6_0 & u_CSAwallace_pg_rca12_and_5_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa6_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa6_xor0 ^ u_CSAwallace_pg_rca12_and_4_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa6_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa6_xor0 & u_CSAwallace_pg_rca12_and_4_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa6_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa6_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa6_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa7_xor0 = u_CSAwallace_pg_rca12_and_7_0 ^ u_CSAwallace_pg_rca12_and_6_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa7_and0 = u_CSAwallace_pg_rca12_and_7_0 & u_CSAwallace_pg_rca12_and_6_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa7_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa7_xor0 ^ u_CSAwallace_pg_rca12_and_5_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa7_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa7_xor0 & u_CSAwallace_pg_rca12_and_5_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa7_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa7_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa7_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa8_xor0 = u_CSAwallace_pg_rca12_and_8_0 ^ u_CSAwallace_pg_rca12_and_7_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa8_and0 = u_CSAwallace_pg_rca12_and_8_0 & u_CSAwallace_pg_rca12_and_7_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa8_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa8_xor0 ^ u_CSAwallace_pg_rca12_and_6_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa8_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa8_xor0 & u_CSAwallace_pg_rca12_and_6_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa8_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa8_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa8_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa9_xor0 = u_CSAwallace_pg_rca12_and_9_0 ^ u_CSAwallace_pg_rca12_and_8_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa9_and0 = u_CSAwallace_pg_rca12_and_9_0 & u_CSAwallace_pg_rca12_and_8_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa9_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa9_xor0 ^ u_CSAwallace_pg_rca12_and_7_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa9_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa9_xor0 & u_CSAwallace_pg_rca12_and_7_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa9_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa9_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa9_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_and_10_0 ^ u_CSAwallace_pg_rca12_and_9_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_and_10_0 & u_CSAwallace_pg_rca12_and_9_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa10_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa10_xor0 ^ u_CSAwallace_pg_rca12_and_8_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa10_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa10_xor0 & u_CSAwallace_pg_rca12_and_8_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa10_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa10_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa10_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_and_11_0 ^ u_CSAwallace_pg_rca12_and_10_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_and_11_0 & u_CSAwallace_pg_rca12_and_10_1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_and_9_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa0_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_and_9_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa0_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_and_11_1 ^ u_CSAwallace_pg_rca12_and_10_2;
  assign u_CSAwallace_pg_rca12_csa0_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_and_11_1 & u_CSAwallace_pg_rca12_and_10_2;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa4_xor0 = u_CSAwallace_pg_rca12_and_1_3 ^ u_CSAwallace_pg_rca12_and_0_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa4_and0 = u_CSAwallace_pg_rca12_and_1_3 & u_CSAwallace_pg_rca12_and_0_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa5_xor0 = u_CSAwallace_pg_rca12_and_2_3 ^ u_CSAwallace_pg_rca12_and_1_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa5_and0 = u_CSAwallace_pg_rca12_and_2_3 & u_CSAwallace_pg_rca12_and_1_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa5_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa5_xor0 ^ u_CSAwallace_pg_rca12_and_0_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa5_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa5_xor0 & u_CSAwallace_pg_rca12_and_0_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa5_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa5_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa5_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa6_xor0 = u_CSAwallace_pg_rca12_and_3_3 ^ u_CSAwallace_pg_rca12_and_2_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa6_and0 = u_CSAwallace_pg_rca12_and_3_3 & u_CSAwallace_pg_rca12_and_2_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa6_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa6_xor0 ^ u_CSAwallace_pg_rca12_and_1_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa6_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa6_xor0 & u_CSAwallace_pg_rca12_and_1_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa6_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa6_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa6_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa7_xor0 = u_CSAwallace_pg_rca12_and_4_3 ^ u_CSAwallace_pg_rca12_and_3_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa7_and0 = u_CSAwallace_pg_rca12_and_4_3 & u_CSAwallace_pg_rca12_and_3_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa7_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa7_xor0 ^ u_CSAwallace_pg_rca12_and_2_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa7_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa7_xor0 & u_CSAwallace_pg_rca12_and_2_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa7_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa7_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa7_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa8_xor0 = u_CSAwallace_pg_rca12_and_5_3 ^ u_CSAwallace_pg_rca12_and_4_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa8_and0 = u_CSAwallace_pg_rca12_and_5_3 & u_CSAwallace_pg_rca12_and_4_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa8_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa8_xor0 ^ u_CSAwallace_pg_rca12_and_3_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa8_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa8_xor0 & u_CSAwallace_pg_rca12_and_3_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa8_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa8_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa8_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa9_xor0 = u_CSAwallace_pg_rca12_and_6_3 ^ u_CSAwallace_pg_rca12_and_5_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa9_and0 = u_CSAwallace_pg_rca12_and_6_3 & u_CSAwallace_pg_rca12_and_5_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa9_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa9_xor0 ^ u_CSAwallace_pg_rca12_and_4_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa9_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa9_xor0 & u_CSAwallace_pg_rca12_and_4_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa9_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa9_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa9_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_and_7_3 ^ u_CSAwallace_pg_rca12_and_6_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_and_7_3 & u_CSAwallace_pg_rca12_and_6_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa10_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa10_xor0 ^ u_CSAwallace_pg_rca12_and_5_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa10_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa10_xor0 & u_CSAwallace_pg_rca12_and_5_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa10_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa10_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa10_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_and_8_3 ^ u_CSAwallace_pg_rca12_and_7_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_and_8_3 & u_CSAwallace_pg_rca12_and_7_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_and_6_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_and_6_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa12_xor0 = u_CSAwallace_pg_rca12_and_9_3 ^ u_CSAwallace_pg_rca12_and_8_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa12_and0 = u_CSAwallace_pg_rca12_and_9_3 & u_CSAwallace_pg_rca12_and_8_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa12_xor0 ^ u_CSAwallace_pg_rca12_and_7_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa12_xor0 & u_CSAwallace_pg_rca12_and_7_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa12_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa12_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa13_xor0 = u_CSAwallace_pg_rca12_and_10_3 ^ u_CSAwallace_pg_rca12_and_9_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa13_and0 = u_CSAwallace_pg_rca12_and_10_3 & u_CSAwallace_pg_rca12_and_9_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa13_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa13_xor0 ^ u_CSAwallace_pg_rca12_and_8_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa13_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa13_xor0 & u_CSAwallace_pg_rca12_and_8_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa13_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa13_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa13_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa14_xor0 = u_CSAwallace_pg_rca12_and_11_3 ^ u_CSAwallace_pg_rca12_and_10_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa14_and0 = u_CSAwallace_pg_rca12_and_11_3 & u_CSAwallace_pg_rca12_and_10_4;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa14_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa14_xor0 ^ u_CSAwallace_pg_rca12_and_9_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa14_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa14_xor0 & u_CSAwallace_pg_rca12_and_9_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa14_or0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa14_and0 | u_CSAwallace_pg_rca12_csa1_csa_component_fa14_and1;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa15_xor1 = u_CSAwallace_pg_rca12_and_11_4 ^ u_CSAwallace_pg_rca12_and_10_5;
  assign u_CSAwallace_pg_rca12_csa1_csa_component_fa15_and1 = u_CSAwallace_pg_rca12_and_11_4 & u_CSAwallace_pg_rca12_and_10_5;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa7_xor0 = u_CSAwallace_pg_rca12_and_1_6 ^ u_CSAwallace_pg_rca12_and_0_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa7_and0 = u_CSAwallace_pg_rca12_and_1_6 & u_CSAwallace_pg_rca12_and_0_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa8_xor0 = u_CSAwallace_pg_rca12_and_2_6 ^ u_CSAwallace_pg_rca12_and_1_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa8_and0 = u_CSAwallace_pg_rca12_and_2_6 & u_CSAwallace_pg_rca12_and_1_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa8_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa8_xor0 ^ u_CSAwallace_pg_rca12_and_0_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa8_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa8_xor0 & u_CSAwallace_pg_rca12_and_0_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa8_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa8_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa8_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa9_xor0 = u_CSAwallace_pg_rca12_and_3_6 ^ u_CSAwallace_pg_rca12_and_2_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa9_and0 = u_CSAwallace_pg_rca12_and_3_6 & u_CSAwallace_pg_rca12_and_2_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa9_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa9_xor0 ^ u_CSAwallace_pg_rca12_and_1_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa9_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa9_xor0 & u_CSAwallace_pg_rca12_and_1_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa9_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa9_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa9_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_and_4_6 ^ u_CSAwallace_pg_rca12_and_3_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_and_4_6 & u_CSAwallace_pg_rca12_and_3_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa10_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa10_xor0 ^ u_CSAwallace_pg_rca12_and_2_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa10_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa10_xor0 & u_CSAwallace_pg_rca12_and_2_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa10_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa10_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa10_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_and_5_6 ^ u_CSAwallace_pg_rca12_and_4_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_and_5_6 & u_CSAwallace_pg_rca12_and_4_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_and_3_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_and_3_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa12_xor0 = u_CSAwallace_pg_rca12_and_6_6 ^ u_CSAwallace_pg_rca12_and_5_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa12_and0 = u_CSAwallace_pg_rca12_and_6_6 & u_CSAwallace_pg_rca12_and_5_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa12_xor0 ^ u_CSAwallace_pg_rca12_and_4_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa12_xor0 & u_CSAwallace_pg_rca12_and_4_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa12_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa12_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa13_xor0 = u_CSAwallace_pg_rca12_and_7_6 ^ u_CSAwallace_pg_rca12_and_6_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa13_and0 = u_CSAwallace_pg_rca12_and_7_6 & u_CSAwallace_pg_rca12_and_6_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa13_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa13_xor0 ^ u_CSAwallace_pg_rca12_and_5_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa13_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa13_xor0 & u_CSAwallace_pg_rca12_and_5_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa13_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa13_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa13_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa14_xor0 = u_CSAwallace_pg_rca12_and_8_6 ^ u_CSAwallace_pg_rca12_and_7_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa14_and0 = u_CSAwallace_pg_rca12_and_8_6 & u_CSAwallace_pg_rca12_and_7_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa14_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa14_xor0 ^ u_CSAwallace_pg_rca12_and_6_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa14_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa14_xor0 & u_CSAwallace_pg_rca12_and_6_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa14_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa14_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa14_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa15_xor0 = u_CSAwallace_pg_rca12_and_9_6 ^ u_CSAwallace_pg_rca12_and_8_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa15_and0 = u_CSAwallace_pg_rca12_and_9_6 & u_CSAwallace_pg_rca12_and_8_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa15_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa15_xor0 ^ u_CSAwallace_pg_rca12_and_7_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa15_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa15_xor0 & u_CSAwallace_pg_rca12_and_7_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa15_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa15_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa15_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa16_xor0 = u_CSAwallace_pg_rca12_and_10_6 ^ u_CSAwallace_pg_rca12_and_9_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa16_and0 = u_CSAwallace_pg_rca12_and_10_6 & u_CSAwallace_pg_rca12_and_9_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa16_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa16_xor0 ^ u_CSAwallace_pg_rca12_and_8_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa16_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa16_xor0 & u_CSAwallace_pg_rca12_and_8_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa16_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa16_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa16_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa17_xor0 = u_CSAwallace_pg_rca12_and_11_6 ^ u_CSAwallace_pg_rca12_and_10_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa17_and0 = u_CSAwallace_pg_rca12_and_11_6 & u_CSAwallace_pg_rca12_and_10_7;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa17_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa17_xor0 ^ u_CSAwallace_pg_rca12_and_9_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa17_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa17_xor0 & u_CSAwallace_pg_rca12_and_9_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa17_or0 = u_CSAwallace_pg_rca12_csa2_csa_component_fa17_and0 | u_CSAwallace_pg_rca12_csa2_csa_component_fa17_and1;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa18_xor1 = u_CSAwallace_pg_rca12_and_11_7 ^ u_CSAwallace_pg_rca12_and_10_8;
  assign u_CSAwallace_pg_rca12_csa2_csa_component_fa18_and1 = u_CSAwallace_pg_rca12_and_11_7 & u_CSAwallace_pg_rca12_and_10_8;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_and_1_9 ^ u_CSAwallace_pg_rca12_and_0_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_and_1_9 & u_CSAwallace_pg_rca12_and_0_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_and_2_9 ^ u_CSAwallace_pg_rca12_and_1_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_and_2_9 & u_CSAwallace_pg_rca12_and_1_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_and_0_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_and_0_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa12_xor0 = u_CSAwallace_pg_rca12_and_3_9 ^ u_CSAwallace_pg_rca12_and_2_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa12_and0 = u_CSAwallace_pg_rca12_and_3_9 & u_CSAwallace_pg_rca12_and_2_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa12_xor0 ^ u_CSAwallace_pg_rca12_and_1_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa12_xor0 & u_CSAwallace_pg_rca12_and_1_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa12_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa12_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa13_xor0 = u_CSAwallace_pg_rca12_and_4_9 ^ u_CSAwallace_pg_rca12_and_3_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa13_and0 = u_CSAwallace_pg_rca12_and_4_9 & u_CSAwallace_pg_rca12_and_3_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa13_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa13_xor0 ^ u_CSAwallace_pg_rca12_and_2_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa13_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa13_xor0 & u_CSAwallace_pg_rca12_and_2_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa13_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa13_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa13_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa14_xor0 = u_CSAwallace_pg_rca12_and_5_9 ^ u_CSAwallace_pg_rca12_and_4_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa14_and0 = u_CSAwallace_pg_rca12_and_5_9 & u_CSAwallace_pg_rca12_and_4_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa14_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa14_xor0 ^ u_CSAwallace_pg_rca12_and_3_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa14_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa14_xor0 & u_CSAwallace_pg_rca12_and_3_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa14_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa14_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa14_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa15_xor0 = u_CSAwallace_pg_rca12_and_6_9 ^ u_CSAwallace_pg_rca12_and_5_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa15_and0 = u_CSAwallace_pg_rca12_and_6_9 & u_CSAwallace_pg_rca12_and_5_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa15_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa15_xor0 ^ u_CSAwallace_pg_rca12_and_4_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa15_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa15_xor0 & u_CSAwallace_pg_rca12_and_4_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa15_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa15_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa15_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa16_xor0 = u_CSAwallace_pg_rca12_and_7_9 ^ u_CSAwallace_pg_rca12_and_6_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa16_and0 = u_CSAwallace_pg_rca12_and_7_9 & u_CSAwallace_pg_rca12_and_6_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa16_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa16_xor0 ^ u_CSAwallace_pg_rca12_and_5_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa16_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa16_xor0 & u_CSAwallace_pg_rca12_and_5_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa16_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa16_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa16_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa17_xor0 = u_CSAwallace_pg_rca12_and_8_9 ^ u_CSAwallace_pg_rca12_and_7_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa17_and0 = u_CSAwallace_pg_rca12_and_8_9 & u_CSAwallace_pg_rca12_and_7_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa17_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa17_xor0 ^ u_CSAwallace_pg_rca12_and_6_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa17_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa17_xor0 & u_CSAwallace_pg_rca12_and_6_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa17_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa17_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa17_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa18_xor0 = u_CSAwallace_pg_rca12_and_9_9 ^ u_CSAwallace_pg_rca12_and_8_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa18_and0 = u_CSAwallace_pg_rca12_and_9_9 & u_CSAwallace_pg_rca12_and_8_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa18_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa18_xor0 ^ u_CSAwallace_pg_rca12_and_7_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa18_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa18_xor0 & u_CSAwallace_pg_rca12_and_7_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa18_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa18_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa18_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa19_xor0 = u_CSAwallace_pg_rca12_and_10_9 ^ u_CSAwallace_pg_rca12_and_9_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa19_and0 = u_CSAwallace_pg_rca12_and_10_9 & u_CSAwallace_pg_rca12_and_9_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa19_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa19_xor0 ^ u_CSAwallace_pg_rca12_and_8_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa19_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa19_xor0 & u_CSAwallace_pg_rca12_and_8_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa19_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa19_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa19_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa20_xor0 = u_CSAwallace_pg_rca12_and_11_9 ^ u_CSAwallace_pg_rca12_and_10_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa20_and0 = u_CSAwallace_pg_rca12_and_11_9 & u_CSAwallace_pg_rca12_and_10_10;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa20_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa20_xor0 ^ u_CSAwallace_pg_rca12_and_9_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa20_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa20_xor0 & u_CSAwallace_pg_rca12_and_9_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa20_or0 = u_CSAwallace_pg_rca12_csa3_csa_component_fa20_and0 | u_CSAwallace_pg_rca12_csa3_csa_component_fa20_and1;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa21_xor1 = u_CSAwallace_pg_rca12_and_11_10 ^ u_CSAwallace_pg_rca12_and_10_11;
  assign u_CSAwallace_pg_rca12_csa3_csa_component_fa21_and1 = u_CSAwallace_pg_rca12_and_11_10 & u_CSAwallace_pg_rca12_and_10_11;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa2_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa2_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa2_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa2_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa3_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa3_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa3_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa3_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa3_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa3_xor0 ^ u_CSAwallace_pg_rca12_and_0_3;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa3_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa3_xor0 & u_CSAwallace_pg_rca12_and_0_3;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa3_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa3_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa3_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa4_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa4_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa4_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa4_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa4_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa4_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa4_xor0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa4_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa4_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa4_xor0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa4_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa4_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa4_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa5_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa5_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa4_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa5_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa5_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa4_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa5_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa5_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa5_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa5_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa5_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa5_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa5_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa5_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa5_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa6_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa6_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa5_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa6_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa6_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa5_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa6_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa6_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa6_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa6_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa6_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa6_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa6_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa6_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa6_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa7_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa7_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa6_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa7_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa7_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa6_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa7_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa7_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa7_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa7_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa7_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa7_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa7_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa7_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa7_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa8_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa8_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa7_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa8_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa8_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa7_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa8_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa8_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa8_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa8_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa8_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa8_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa8_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa8_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa8_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa9_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa9_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa9_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa9_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa9_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa9_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa9_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa9_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa9_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa9_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa9_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa9_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa9_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa10_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa10_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa10_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa10_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa10_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa10_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa10_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa10_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa10_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa10_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa10_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa11_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa11_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa12_xor0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa12_xor1 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa12_and0 = u_CSAwallace_pg_rca12_csa0_csa_component_fa12_xor1 & u_CSAwallace_pg_rca12_csa0_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa12_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa12_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa12_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa12_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa13_xor0 = u_CSAwallace_pg_rca12_and_11_2 ^ u_CSAwallace_pg_rca12_csa0_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa13_and0 = u_CSAwallace_pg_rca12_and_11_2 & u_CSAwallace_pg_rca12_csa0_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa13_xor1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa13_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa13_and1 = u_CSAwallace_pg_rca12_csa4_csa_component_fa13_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa4_csa_component_fa13_or0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa13_and0 | u_CSAwallace_pg_rca12_csa4_csa_component_fa13_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa6_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa5_or0 ^ u_CSAwallace_pg_rca12_and_0_6;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa6_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa5_or0 & u_CSAwallace_pg_rca12_and_0_6;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa7_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa6_or0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa7_xor0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa7_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa6_or0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa7_xor0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa8_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa7_or0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa8_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa8_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa7_or0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa8_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa8_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa8_xor0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa7_and0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa8_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa8_xor0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa7_and0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa8_or0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa8_and0 | u_CSAwallace_pg_rca12_csa5_csa_component_fa8_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa9_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa8_or0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa9_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa9_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa8_or0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa9_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa9_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa9_xor0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa9_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa9_xor0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa9_or0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa9_and0 | u_CSAwallace_pg_rca12_csa5_csa_component_fa9_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa9_or0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa10_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa9_or0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa10_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa10_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa10_xor0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa10_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa10_xor0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa10_or0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa10_and0 | u_CSAwallace_pg_rca12_csa5_csa_component_fa10_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa10_or0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa10_or0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa5_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa12_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa11_or0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa12_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa11_or0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa12_xor0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa12_xor0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa12_or0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa12_and0 | u_CSAwallace_pg_rca12_csa5_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa13_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa12_or0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa13_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa12_or0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa13_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa13_xor0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa13_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa13_xor0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa13_or0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa13_and0 | u_CSAwallace_pg_rca12_csa5_csa_component_fa13_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa14_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa13_or0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa14_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa14_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa13_or0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa14_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa14_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa14_xor0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa14_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa14_xor0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa14_or0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa14_and0 | u_CSAwallace_pg_rca12_csa5_csa_component_fa14_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa15_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa14_or0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa15_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa15_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa14_or0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa15_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa15_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa15_xor0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa15_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa15_xor0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa15_or0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa15_and0 | u_CSAwallace_pg_rca12_csa5_csa_component_fa15_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa16_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa15_and1 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa16_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa16_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa15_and1 & u_CSAwallace_pg_rca12_csa2_csa_component_fa16_xor1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa16_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa16_xor0 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa16_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa16_xor0 & u_CSAwallace_pg_rca12_csa2_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa16_or0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa16_and0 | u_CSAwallace_pg_rca12_csa5_csa_component_fa16_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa17_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa17_xor1 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa17_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa17_xor1 & u_CSAwallace_pg_rca12_csa2_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa18_xor1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa18_xor1 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa18_and1 = u_CSAwallace_pg_rca12_csa2_csa_component_fa18_xor1 & u_CSAwallace_pg_rca12_csa2_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa19_xor1 = u_CSAwallace_pg_rca12_and_11_8 ^ u_CSAwallace_pg_rca12_csa2_csa_component_fa18_and1;
  assign u_CSAwallace_pg_rca12_csa5_csa_component_fa19_and1 = u_CSAwallace_pg_rca12_and_11_8 & u_CSAwallace_pg_rca12_csa2_csa_component_fa18_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa3_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa3_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa2_and0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa3_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa3_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa2_and0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa4_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa4_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa3_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa4_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa4_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa3_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa5_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa5_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa4_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa5_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa5_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa4_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa5_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa5_xor0 ^ u_CSAwallace_pg_rca12_csa1_csa_component_fa4_and0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa5_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa5_xor0 & u_CSAwallace_pg_rca12_csa1_csa_component_fa4_and0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa5_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa5_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa5_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa6_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa6_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa5_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa6_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa6_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa5_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa6_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa6_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa6_xor0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa6_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa6_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa6_xor0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa6_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa6_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa6_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa7_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa7_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa6_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa7_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa7_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa6_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa7_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa7_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa7_xor0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa7_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa7_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa7_xor0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa7_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa7_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa7_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa8_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa8_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa7_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa8_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa8_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa7_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa8_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa8_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa8_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa8_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa8_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa8_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa8_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa8_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa8_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa9_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa9_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa9_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa9_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa9_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa9_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa9_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa9_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa9_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa9_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa9_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa9_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa9_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa10_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa10_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa10_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa10_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa10_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa10_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa10_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa10_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa10_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa10_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa10_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa11_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa11_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa12_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa12_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa12_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa12_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa12_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa12_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa12_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa12_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa13_xor0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa13_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa13_and0 = u_CSAwallace_pg_rca12_csa4_csa_component_fa13_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa13_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa13_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa13_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa13_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa13_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa13_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa13_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa14_xor0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa14_xor1 ^ u_CSAwallace_pg_rca12_csa4_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa14_and0 = u_CSAwallace_pg_rca12_csa1_csa_component_fa14_xor1 & u_CSAwallace_pg_rca12_csa4_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa14_xor1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa14_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa14_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa14_and1 = u_CSAwallace_pg_rca12_csa6_csa_component_fa14_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa14_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa14_or0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa14_and0 | u_CSAwallace_pg_rca12_csa6_csa_component_fa14_and1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa15_xor1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa15_xor1 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa15_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa15_and1 = u_CSAwallace_pg_rca12_csa1_csa_component_fa15_xor1 & u_CSAwallace_pg_rca12_csa5_csa_component_fa15_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa16_xor1 = u_CSAwallace_pg_rca12_and_11_5 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa16_xor1;
  assign u_CSAwallace_pg_rca12_csa6_csa_component_fa16_and1 = u_CSAwallace_pg_rca12_and_11_5 & u_CSAwallace_pg_rca12_csa5_csa_component_fa16_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa9_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa8_or0 ^ u_CSAwallace_pg_rca12_and_0_9;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa9_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa8_or0 & u_CSAwallace_pg_rca12_and_0_9;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa9_or0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa10_xor0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa9_or0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa10_xor0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa10_or0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa10_or0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa10_and0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa10_and0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa12_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa11_or0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa12_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa11_or0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa12_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa12_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa12_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa12_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa13_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa12_or0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa13_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa12_or0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa13_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa13_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa13_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa13_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa13_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa13_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa13_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa14_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa13_or0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa14_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa14_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa13_or0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa14_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa14_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa14_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa14_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa14_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa14_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa14_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa14_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa15_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa14_or0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa15_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa15_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa14_or0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa15_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa15_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa15_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa15_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa15_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa15_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa15_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa15_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa16_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa15_or0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa16_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa16_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa15_or0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa16_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa16_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa16_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa16_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa16_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa16_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa16_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa16_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa17_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa16_or0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa17_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa17_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa16_or0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa17_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa17_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa17_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa17_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa17_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa17_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa17_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa17_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa18_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa17_and1 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa18_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa18_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa17_and1 & u_CSAwallace_pg_rca12_csa3_csa_component_fa18_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa18_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa18_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa18_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa18_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa18_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa18_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa18_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa19_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa18_and1 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa19_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa19_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa18_and1 & u_CSAwallace_pg_rca12_csa3_csa_component_fa19_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa19_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa19_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa18_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa19_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa19_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa18_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa19_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa19_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa19_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa20_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa19_and1 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa20_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa20_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa19_and1 & u_CSAwallace_pg_rca12_csa3_csa_component_fa20_xor1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa20_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa20_xor0 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa19_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa20_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa20_xor0 & u_CSAwallace_pg_rca12_csa3_csa_component_fa19_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa20_or0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa20_and0 | u_CSAwallace_pg_rca12_csa7_csa_component_fa20_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa21_xor1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa21_xor1 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa20_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa21_and1 = u_CSAwallace_pg_rca12_csa3_csa_component_fa21_xor1 & u_CSAwallace_pg_rca12_csa3_csa_component_fa20_or0;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa22_xor1 = u_CSAwallace_pg_rca12_and_11_11 ^ u_CSAwallace_pg_rca12_csa3_csa_component_fa21_and1;
  assign u_CSAwallace_pg_rca12_csa7_csa_component_fa22_and1 = u_CSAwallace_pg_rca12_and_11_11 & u_CSAwallace_pg_rca12_csa3_csa_component_fa21_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa4_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa4_xor0 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa3_and0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa4_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa4_xor0 & u_CSAwallace_pg_rca12_csa6_csa_component_fa3_and0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa5_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa5_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa4_and0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa5_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa5_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa4_and0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa6_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa6_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa5_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa6_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa6_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa5_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa7_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa7_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa6_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa7_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa7_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa6_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa7_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa7_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa6_and0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa7_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa7_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa6_and0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa7_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa7_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa7_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa8_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa8_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa7_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa8_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa8_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa7_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa8_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa8_xor0 ^ u_CSAwallace_pg_rca12_csa5_csa_component_fa7_and0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa8_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa8_xor0 & u_CSAwallace_pg_rca12_csa5_csa_component_fa7_and0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa8_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa8_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa8_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa9_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa9_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa9_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa9_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa9_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa9_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa9_xor0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa9_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa9_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa9_xor0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa9_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa9_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa9_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa10_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa10_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa10_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa10_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa10_xor0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa10_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa10_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa10_xor0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa10_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa10_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa10_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa11_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa11_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa11_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa12_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa12_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa12_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa12_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa12_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa12_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa12_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa12_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa12_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa13_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa13_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa13_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa13_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa13_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa13_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa13_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa13_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa13_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa13_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa13_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa13_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa14_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa14_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa14_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa14_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa14_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa14_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa14_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa14_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa14_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa14_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa14_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa14_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa14_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa15_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa15_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa15_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa15_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa15_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa15_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa15_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa15_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa15_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa15_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa15_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa15_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa15_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa16_xor0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa16_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa15_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa16_and0 = u_CSAwallace_pg_rca12_csa6_csa_component_fa16_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa15_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa16_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa16_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa16_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa16_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa16_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa16_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa16_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa16_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa16_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa17_xor0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa17_xor1 ^ u_CSAwallace_pg_rca12_csa6_csa_component_fa16_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa17_and0 = u_CSAwallace_pg_rca12_csa5_csa_component_fa17_xor1 & u_CSAwallace_pg_rca12_csa6_csa_component_fa16_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa17_xor1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa17_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa17_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa17_and1 = u_CSAwallace_pg_rca12_csa8_csa_component_fa17_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa17_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa17_or0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa17_and0 | u_CSAwallace_pg_rca12_csa8_csa_component_fa17_and1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa18_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa18_xor1 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa18_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa18_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa18_xor1 & u_CSAwallace_pg_rca12_csa7_csa_component_fa18_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa19_xor1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa19_xor1 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa19_xor1;
  assign u_CSAwallace_pg_rca12_csa8_csa_component_fa19_and1 = u_CSAwallace_pg_rca12_csa5_csa_component_fa19_xor1 & u_CSAwallace_pg_rca12_csa7_csa_component_fa19_xor1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa5_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa5_xor0 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa4_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa5_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa5_xor0 & u_CSAwallace_pg_rca12_csa8_csa_component_fa4_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa6_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa6_xor0 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa5_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa6_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa6_xor0 & u_CSAwallace_pg_rca12_csa8_csa_component_fa5_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa7_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa7_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa6_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa7_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa7_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa6_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa8_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa8_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa7_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa8_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa8_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa7_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa9_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa9_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa9_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa9_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa8_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa10_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa10_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa10_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa10_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa9_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa10_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa10_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa9_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa10_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa10_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa9_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa10_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa10_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa10_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa11_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa11_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa11_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa11_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa11_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa11_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa10_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa11_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa11_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa10_and0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa11_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa11_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa11_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa12_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa12_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa12_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa12_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa12_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa12_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa12_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa12_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa12_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa12_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa12_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa13_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa13_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa13_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa13_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa13_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa13_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa13_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa13_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa13_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa13_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa13_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa14_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa14_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa14_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa14_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa14_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa14_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa14_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa14_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa14_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa14_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa14_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa15_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa15_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa15_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa15_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa15_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa15_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa15_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa15_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa15_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa15_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa15_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa16_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa16_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa16_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa16_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa16_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa16_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa16_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa16_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa16_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa16_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa16_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa17_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa17_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa17_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa17_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa17_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa17_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa17_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa17_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa17_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa17_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa17_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa18_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa18_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa18_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa18_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa18_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa18_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa18_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa18_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa18_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa18_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa18_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa19_xor0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa19_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa18_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa19_and0 = u_CSAwallace_pg_rca12_csa8_csa_component_fa19_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa18_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa19_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa19_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa18_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa19_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa19_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa18_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa19_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa19_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa19_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa20_xor0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa20_xor1 ^ u_CSAwallace_pg_rca12_csa8_csa_component_fa19_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa20_and0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa20_xor1 & u_CSAwallace_pg_rca12_csa8_csa_component_fa19_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa20_xor1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa20_xor0 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa19_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa20_and1 = u_CSAwallace_pg_rca12_csa9_csa_component_fa20_xor0 & u_CSAwallace_pg_rca12_csa7_csa_component_fa19_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa20_or0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa20_and0 | u_CSAwallace_pg_rca12_csa9_csa_component_fa20_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa21_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa21_xor1 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa20_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa21_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa21_xor1 & u_CSAwallace_pg_rca12_csa7_csa_component_fa20_or0;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa22_xor1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa22_xor1 ^ u_CSAwallace_pg_rca12_csa7_csa_component_fa21_and1;
  assign u_CSAwallace_pg_rca12_csa9_csa_component_fa22_and1 = u_CSAwallace_pg_rca12_csa7_csa_component_fa22_xor1 & u_CSAwallace_pg_rca12_csa7_csa_component_fa21_and1;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa6_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa6_xor0 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa5_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa6_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa6_xor0 & u_CSAwallace_pg_rca12_csa9_csa_component_fa5_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa7_xor0 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa6_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa7_xor0 & u_CSAwallace_pg_rca12_csa9_csa_component_fa6_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa6_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and7 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa6_and0 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or7 = u_CSAwallace_pg_rca12_u_pg_rca24_and7 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa8_xor0 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa7_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa8_xor0 & u_CSAwallace_pg_rca12_csa9_csa_component_fa7_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or7;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and8 = u_CSAwallace_pg_rca12_u_pg_rca24_or7 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or8 = u_CSAwallace_pg_rca12_u_pg_rca24_and8 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa9_xor0 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa8_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa9_xor0 & u_CSAwallace_pg_rca12_csa9_csa_component_fa8_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or8;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and9 = u_CSAwallace_pg_rca12_u_pg_rca24_or8 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or9 = u_CSAwallace_pg_rca12_u_pg_rca24_and9 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa10_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa9_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa10_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa9_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or9;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and10 = u_CSAwallace_pg_rca12_u_pg_rca24_or9 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or10 = u_CSAwallace_pg_rca12_u_pg_rca24_and10 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa11_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa11_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa10_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or10;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and11 = u_CSAwallace_pg_rca12_u_pg_rca24_or10 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or11 = u_CSAwallace_pg_rca12_u_pg_rca24_and11 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa12_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa12_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa11_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or11;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and12 = u_CSAwallace_pg_rca12_u_pg_rca24_or11 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or12 = u_CSAwallace_pg_rca12_u_pg_rca24_and12 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa13_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa13_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa12_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or12;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and13 = u_CSAwallace_pg_rca12_u_pg_rca24_or12 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or13 = u_CSAwallace_pg_rca12_u_pg_rca24_and13 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa14_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa14_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa13_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or13;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and14 = u_CSAwallace_pg_rca12_u_pg_rca24_or13 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or14 = u_CSAwallace_pg_rca12_u_pg_rca24_and14 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa15_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa15_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa14_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or14;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and15 = u_CSAwallace_pg_rca12_u_pg_rca24_or14 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or15 = u_CSAwallace_pg_rca12_u_pg_rca24_and15 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa16_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa16_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa15_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or15;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and16 = u_CSAwallace_pg_rca12_u_pg_rca24_or15 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or16 = u_CSAwallace_pg_rca12_u_pg_rca24_and16 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa17_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa17_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa16_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or16;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and17 = u_CSAwallace_pg_rca12_u_pg_rca24_or16 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or17 = u_CSAwallace_pg_rca12_u_pg_rca24_and17 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa18_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa18_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa17_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or17;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and18 = u_CSAwallace_pg_rca12_u_pg_rca24_or17 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or18 = u_CSAwallace_pg_rca12_u_pg_rca24_and18 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa19_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa18_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa19_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa18_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or18;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and19 = u_CSAwallace_pg_rca12_u_pg_rca24_or18 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or19 = u_CSAwallace_pg_rca12_u_pg_rca24_and19 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa20_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa19_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa20_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa19_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or19;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and20 = u_CSAwallace_pg_rca12_u_pg_rca24_or19 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or20 = u_CSAwallace_pg_rca12_u_pg_rca24_and20 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa21_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa20_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa21_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa20_or0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or20;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and21 = u_CSAwallace_pg_rca12_u_pg_rca24_or20 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or21 = u_CSAwallace_pg_rca12_u_pg_rca24_and21 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_xor0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa22_xor1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa21_and1;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_and0 = u_CSAwallace_pg_rca12_csa9_csa_component_fa22_xor1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa21_and1;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or21;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and22 = u_CSAwallace_pg_rca12_u_pg_rca24_or21 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or22 = u_CSAwallace_pg_rca12_u_pg_rca24_and22 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_and0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_xor0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa22_and1 ^ u_CSAwallace_pg_rca12_csa9_csa_component_fa22_and1;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_and0 = u_CSAwallace_pg_rca12_csa7_csa_component_fa22_and1 & u_CSAwallace_pg_rca12_csa9_csa_component_fa22_and1;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_xor1 = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_xor0 ^ u_CSAwallace_pg_rca12_u_pg_rca24_or22;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_and23 = u_CSAwallace_pg_rca12_u_pg_rca24_or22 & u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_xor0;
  assign u_CSAwallace_pg_rca12_u_pg_rca24_or23 = u_CSAwallace_pg_rca12_u_pg_rca24_and23 | u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_and0;

  assign u_CSAwallace_pg_rca12_out[0] = u_CSAwallace_pg_rca12_and_0_0;
  assign u_CSAwallace_pg_rca12_out[1] = u_CSAwallace_pg_rca12_csa0_csa_component_fa1_xor0;
  assign u_CSAwallace_pg_rca12_out[2] = u_CSAwallace_pg_rca12_csa4_csa_component_fa2_xor0;
  assign u_CSAwallace_pg_rca12_out[3] = u_CSAwallace_pg_rca12_csa6_csa_component_fa3_xor0;
  assign u_CSAwallace_pg_rca12_out[4] = u_CSAwallace_pg_rca12_csa8_csa_component_fa4_xor0;
  assign u_CSAwallace_pg_rca12_out[5] = u_CSAwallace_pg_rca12_csa9_csa_component_fa5_xor0;
  assign u_CSAwallace_pg_rca12_out[6] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa6_xor0;
  assign u_CSAwallace_pg_rca12_out[7] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa7_xor1;
  assign u_CSAwallace_pg_rca12_out[8] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa8_xor1;
  assign u_CSAwallace_pg_rca12_out[9] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa9_xor1;
  assign u_CSAwallace_pg_rca12_out[10] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa10_xor1;
  assign u_CSAwallace_pg_rca12_out[11] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa11_xor1;
  assign u_CSAwallace_pg_rca12_out[12] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa12_xor1;
  assign u_CSAwallace_pg_rca12_out[13] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa13_xor1;
  assign u_CSAwallace_pg_rca12_out[14] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa14_xor1;
  assign u_CSAwallace_pg_rca12_out[15] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa15_xor1;
  assign u_CSAwallace_pg_rca12_out[16] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa16_xor1;
  assign u_CSAwallace_pg_rca12_out[17] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa17_xor1;
  assign u_CSAwallace_pg_rca12_out[18] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa18_xor1;
  assign u_CSAwallace_pg_rca12_out[19] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa19_xor1;
  assign u_CSAwallace_pg_rca12_out[20] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa20_xor1;
  assign u_CSAwallace_pg_rca12_out[21] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa21_xor1;
  assign u_CSAwallace_pg_rca12_out[22] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa22_xor1;
  assign u_CSAwallace_pg_rca12_out[23] = u_CSAwallace_pg_rca12_u_pg_rca24_pg_fa23_xor1;
endmodule