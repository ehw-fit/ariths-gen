module f_s_dadda_rca16(input [15:0] a, input [15:0] b, output [31:0] f_s_dadda_rca16_out);
  wire f_s_dadda_rca16_and_13_0;
  wire f_s_dadda_rca16_and_12_1;
  wire f_s_dadda_rca16_ha0_xor0;
  wire f_s_dadda_rca16_ha0_and0;
  wire f_s_dadda_rca16_and_14_0;
  wire f_s_dadda_rca16_and_13_1;
  wire f_s_dadda_rca16_fa0_xor0;
  wire f_s_dadda_rca16_fa0_and0;
  wire f_s_dadda_rca16_fa0_xor1;
  wire f_s_dadda_rca16_fa0_and1;
  wire f_s_dadda_rca16_fa0_or0;
  wire f_s_dadda_rca16_and_12_2;
  wire f_s_dadda_rca16_and_11_3;
  wire f_s_dadda_rca16_ha1_xor0;
  wire f_s_dadda_rca16_ha1_and0;
  wire f_s_dadda_rca16_nand_15_0;
  wire f_s_dadda_rca16_fa1_xor0;
  wire f_s_dadda_rca16_fa1_and0;
  wire f_s_dadda_rca16_fa1_xor1;
  wire f_s_dadda_rca16_fa1_and1;
  wire f_s_dadda_rca16_fa1_or0;
  wire f_s_dadda_rca16_and_14_1;
  wire f_s_dadda_rca16_and_13_2;
  wire f_s_dadda_rca16_and_12_3;
  wire f_s_dadda_rca16_fa2_xor0;
  wire f_s_dadda_rca16_fa2_and0;
  wire f_s_dadda_rca16_fa2_xor1;
  wire f_s_dadda_rca16_fa2_and1;
  wire f_s_dadda_rca16_fa2_or0;
  wire f_s_dadda_rca16_and_11_4;
  wire f_s_dadda_rca16_and_10_5;
  wire f_s_dadda_rca16_ha2_xor0;
  wire f_s_dadda_rca16_ha2_and0;
  wire f_s_dadda_rca16_fa3_xor0;
  wire f_s_dadda_rca16_fa3_and0;
  wire f_s_dadda_rca16_fa3_xor1;
  wire f_s_dadda_rca16_fa3_and1;
  wire f_s_dadda_rca16_fa3_or0;
  wire f_s_dadda_rca16_nand_15_1;
  wire f_s_dadda_rca16_and_14_2;
  wire f_s_dadda_rca16_fa4_xor0;
  wire f_s_dadda_rca16_fa4_xor1;
  wire f_s_dadda_rca16_fa4_and1;
  wire f_s_dadda_rca16_fa4_or0;
  wire f_s_dadda_rca16_and_13_3;
  wire f_s_dadda_rca16_and_12_4;
  wire f_s_dadda_rca16_and_11_5;
  wire f_s_dadda_rca16_fa5_xor0;
  wire f_s_dadda_rca16_fa5_and0;
  wire f_s_dadda_rca16_fa5_xor1;
  wire f_s_dadda_rca16_fa5_and1;
  wire f_s_dadda_rca16_fa5_or0;
  wire f_s_dadda_rca16_fa6_xor0;
  wire f_s_dadda_rca16_fa6_and0;
  wire f_s_dadda_rca16_fa6_xor1;
  wire f_s_dadda_rca16_fa6_and1;
  wire f_s_dadda_rca16_fa6_or0;
  wire f_s_dadda_rca16_nand_15_2;
  wire f_s_dadda_rca16_and_14_3;
  wire f_s_dadda_rca16_and_13_4;
  wire f_s_dadda_rca16_fa7_xor0;
  wire f_s_dadda_rca16_fa7_and0;
  wire f_s_dadda_rca16_fa7_xor1;
  wire f_s_dadda_rca16_fa7_and1;
  wire f_s_dadda_rca16_fa7_or0;
  wire f_s_dadda_rca16_nand_15_3;
  wire f_s_dadda_rca16_fa8_xor0;
  wire f_s_dadda_rca16_fa8_and0;
  wire f_s_dadda_rca16_fa8_xor1;
  wire f_s_dadda_rca16_fa8_and1;
  wire f_s_dadda_rca16_fa8_or0;
  wire f_s_dadda_rca16_and_4_0;
  wire f_s_dadda_rca16_and_3_1;
  wire f_s_dadda_rca16_ha3_xor0;
  wire f_s_dadda_rca16_ha3_and0;
  wire f_s_dadda_rca16_and_5_0;
  wire f_s_dadda_rca16_and_4_1;
  wire f_s_dadda_rca16_fa9_xor0;
  wire f_s_dadda_rca16_fa9_and0;
  wire f_s_dadda_rca16_fa9_xor1;
  wire f_s_dadda_rca16_fa9_and1;
  wire f_s_dadda_rca16_fa9_or0;
  wire f_s_dadda_rca16_and_3_2;
  wire f_s_dadda_rca16_and_2_3;
  wire f_s_dadda_rca16_ha4_xor0;
  wire f_s_dadda_rca16_ha4_and0;
  wire f_s_dadda_rca16_and_6_0;
  wire f_s_dadda_rca16_fa10_xor0;
  wire f_s_dadda_rca16_fa10_and0;
  wire f_s_dadda_rca16_fa10_xor1;
  wire f_s_dadda_rca16_fa10_and1;
  wire f_s_dadda_rca16_fa10_or0;
  wire f_s_dadda_rca16_and_5_1;
  wire f_s_dadda_rca16_and_4_2;
  wire f_s_dadda_rca16_and_3_3;
  wire f_s_dadda_rca16_fa11_xor0;
  wire f_s_dadda_rca16_fa11_and0;
  wire f_s_dadda_rca16_fa11_xor1;
  wire f_s_dadda_rca16_fa11_and1;
  wire f_s_dadda_rca16_fa11_or0;
  wire f_s_dadda_rca16_and_2_4;
  wire f_s_dadda_rca16_and_1_5;
  wire f_s_dadda_rca16_ha5_xor0;
  wire f_s_dadda_rca16_ha5_and0;
  wire f_s_dadda_rca16_fa12_xor0;
  wire f_s_dadda_rca16_fa12_and0;
  wire f_s_dadda_rca16_fa12_xor1;
  wire f_s_dadda_rca16_fa12_and1;
  wire f_s_dadda_rca16_fa12_or0;
  wire f_s_dadda_rca16_and_7_0;
  wire f_s_dadda_rca16_and_6_1;
  wire f_s_dadda_rca16_and_5_2;
  wire f_s_dadda_rca16_fa13_xor0;
  wire f_s_dadda_rca16_fa13_and0;
  wire f_s_dadda_rca16_fa13_xor1;
  wire f_s_dadda_rca16_fa13_and1;
  wire f_s_dadda_rca16_fa13_or0;
  wire f_s_dadda_rca16_and_4_3;
  wire f_s_dadda_rca16_and_3_4;
  wire f_s_dadda_rca16_and_2_5;
  wire f_s_dadda_rca16_fa14_xor0;
  wire f_s_dadda_rca16_fa14_and0;
  wire f_s_dadda_rca16_fa14_xor1;
  wire f_s_dadda_rca16_fa14_and1;
  wire f_s_dadda_rca16_fa14_or0;
  wire f_s_dadda_rca16_and_1_6;
  wire f_s_dadda_rca16_and_0_7;
  wire f_s_dadda_rca16_ha6_xor0;
  wire f_s_dadda_rca16_ha6_and0;
  wire f_s_dadda_rca16_fa15_xor0;
  wire f_s_dadda_rca16_fa15_and0;
  wire f_s_dadda_rca16_fa15_xor1;
  wire f_s_dadda_rca16_fa15_and1;
  wire f_s_dadda_rca16_fa15_or0;
  wire f_s_dadda_rca16_and_8_0;
  wire f_s_dadda_rca16_and_7_1;
  wire f_s_dadda_rca16_fa16_xor0;
  wire f_s_dadda_rca16_fa16_and0;
  wire f_s_dadda_rca16_fa16_xor1;
  wire f_s_dadda_rca16_fa16_and1;
  wire f_s_dadda_rca16_fa16_or0;
  wire f_s_dadda_rca16_and_6_2;
  wire f_s_dadda_rca16_and_5_3;
  wire f_s_dadda_rca16_and_4_4;
  wire f_s_dadda_rca16_fa17_xor0;
  wire f_s_dadda_rca16_fa17_and0;
  wire f_s_dadda_rca16_fa17_xor1;
  wire f_s_dadda_rca16_fa17_and1;
  wire f_s_dadda_rca16_fa17_or0;
  wire f_s_dadda_rca16_and_3_5;
  wire f_s_dadda_rca16_and_2_6;
  wire f_s_dadda_rca16_and_1_7;
  wire f_s_dadda_rca16_fa18_xor0;
  wire f_s_dadda_rca16_fa18_and0;
  wire f_s_dadda_rca16_fa18_xor1;
  wire f_s_dadda_rca16_fa18_and1;
  wire f_s_dadda_rca16_fa18_or0;
  wire f_s_dadda_rca16_and_0_8;
  wire f_s_dadda_rca16_ha7_xor0;
  wire f_s_dadda_rca16_ha7_and0;
  wire f_s_dadda_rca16_fa19_xor0;
  wire f_s_dadda_rca16_fa19_and0;
  wire f_s_dadda_rca16_fa19_xor1;
  wire f_s_dadda_rca16_fa19_and1;
  wire f_s_dadda_rca16_fa19_or0;
  wire f_s_dadda_rca16_and_9_0;
  wire f_s_dadda_rca16_fa20_xor0;
  wire f_s_dadda_rca16_fa20_and0;
  wire f_s_dadda_rca16_fa20_xor1;
  wire f_s_dadda_rca16_fa20_and1;
  wire f_s_dadda_rca16_fa20_or0;
  wire f_s_dadda_rca16_and_8_1;
  wire f_s_dadda_rca16_and_7_2;
  wire f_s_dadda_rca16_and_6_3;
  wire f_s_dadda_rca16_fa21_xor0;
  wire f_s_dadda_rca16_fa21_and0;
  wire f_s_dadda_rca16_fa21_xor1;
  wire f_s_dadda_rca16_fa21_and1;
  wire f_s_dadda_rca16_fa21_or0;
  wire f_s_dadda_rca16_and_5_4;
  wire f_s_dadda_rca16_and_4_5;
  wire f_s_dadda_rca16_and_3_6;
  wire f_s_dadda_rca16_fa22_xor0;
  wire f_s_dadda_rca16_fa22_and0;
  wire f_s_dadda_rca16_fa22_xor1;
  wire f_s_dadda_rca16_fa22_and1;
  wire f_s_dadda_rca16_fa22_or0;
  wire f_s_dadda_rca16_and_2_7;
  wire f_s_dadda_rca16_and_1_8;
  wire f_s_dadda_rca16_and_0_9;
  wire f_s_dadda_rca16_fa23_xor0;
  wire f_s_dadda_rca16_fa23_and0;
  wire f_s_dadda_rca16_fa23_xor1;
  wire f_s_dadda_rca16_fa23_and1;
  wire f_s_dadda_rca16_fa23_or0;
  wire f_s_dadda_rca16_ha8_xor0;
  wire f_s_dadda_rca16_ha8_and0;
  wire f_s_dadda_rca16_fa24_xor0;
  wire f_s_dadda_rca16_fa24_and0;
  wire f_s_dadda_rca16_fa24_xor1;
  wire f_s_dadda_rca16_fa24_and1;
  wire f_s_dadda_rca16_fa24_or0;
  wire f_s_dadda_rca16_fa25_xor0;
  wire f_s_dadda_rca16_fa25_and0;
  wire f_s_dadda_rca16_fa25_xor1;
  wire f_s_dadda_rca16_fa25_and1;
  wire f_s_dadda_rca16_fa25_or0;
  wire f_s_dadda_rca16_and_10_0;
  wire f_s_dadda_rca16_and_9_1;
  wire f_s_dadda_rca16_and_8_2;
  wire f_s_dadda_rca16_fa26_xor0;
  wire f_s_dadda_rca16_fa26_and0;
  wire f_s_dadda_rca16_fa26_xor1;
  wire f_s_dadda_rca16_fa26_and1;
  wire f_s_dadda_rca16_fa26_or0;
  wire f_s_dadda_rca16_and_7_3;
  wire f_s_dadda_rca16_and_6_4;
  wire f_s_dadda_rca16_and_5_5;
  wire f_s_dadda_rca16_fa27_xor0;
  wire f_s_dadda_rca16_fa27_and0;
  wire f_s_dadda_rca16_fa27_xor1;
  wire f_s_dadda_rca16_fa27_and1;
  wire f_s_dadda_rca16_fa27_or0;
  wire f_s_dadda_rca16_and_4_6;
  wire f_s_dadda_rca16_and_3_7;
  wire f_s_dadda_rca16_and_2_8;
  wire f_s_dadda_rca16_fa28_xor0;
  wire f_s_dadda_rca16_fa28_and0;
  wire f_s_dadda_rca16_fa28_xor1;
  wire f_s_dadda_rca16_fa28_and1;
  wire f_s_dadda_rca16_fa28_or0;
  wire f_s_dadda_rca16_and_1_9;
  wire f_s_dadda_rca16_and_0_10;
  wire f_s_dadda_rca16_fa29_xor0;
  wire f_s_dadda_rca16_fa29_and0;
  wire f_s_dadda_rca16_fa29_xor1;
  wire f_s_dadda_rca16_fa29_and1;
  wire f_s_dadda_rca16_fa29_or0;
  wire f_s_dadda_rca16_ha9_xor0;
  wire f_s_dadda_rca16_ha9_and0;
  wire f_s_dadda_rca16_fa30_xor0;
  wire f_s_dadda_rca16_fa30_and0;
  wire f_s_dadda_rca16_fa30_xor1;
  wire f_s_dadda_rca16_fa30_and1;
  wire f_s_dadda_rca16_fa30_or0;
  wire f_s_dadda_rca16_fa31_xor0;
  wire f_s_dadda_rca16_fa31_and0;
  wire f_s_dadda_rca16_fa31_xor1;
  wire f_s_dadda_rca16_fa31_and1;
  wire f_s_dadda_rca16_fa31_or0;
  wire f_s_dadda_rca16_and_11_0;
  wire f_s_dadda_rca16_and_10_1;
  wire f_s_dadda_rca16_fa32_xor0;
  wire f_s_dadda_rca16_fa32_and0;
  wire f_s_dadda_rca16_fa32_xor1;
  wire f_s_dadda_rca16_fa32_and1;
  wire f_s_dadda_rca16_fa32_or0;
  wire f_s_dadda_rca16_and_9_2;
  wire f_s_dadda_rca16_and_8_3;
  wire f_s_dadda_rca16_and_7_4;
  wire f_s_dadda_rca16_fa33_xor0;
  wire f_s_dadda_rca16_fa33_and0;
  wire f_s_dadda_rca16_fa33_xor1;
  wire f_s_dadda_rca16_fa33_and1;
  wire f_s_dadda_rca16_fa33_or0;
  wire f_s_dadda_rca16_and_6_5;
  wire f_s_dadda_rca16_and_5_6;
  wire f_s_dadda_rca16_and_4_7;
  wire f_s_dadda_rca16_fa34_xor0;
  wire f_s_dadda_rca16_fa34_and0;
  wire f_s_dadda_rca16_fa34_xor1;
  wire f_s_dadda_rca16_fa34_and1;
  wire f_s_dadda_rca16_fa34_or0;
  wire f_s_dadda_rca16_and_3_8;
  wire f_s_dadda_rca16_and_2_9;
  wire f_s_dadda_rca16_and_1_10;
  wire f_s_dadda_rca16_fa35_xor0;
  wire f_s_dadda_rca16_fa35_and0;
  wire f_s_dadda_rca16_fa35_xor1;
  wire f_s_dadda_rca16_fa35_and1;
  wire f_s_dadda_rca16_fa35_or0;
  wire f_s_dadda_rca16_and_0_11;
  wire f_s_dadda_rca16_fa36_xor0;
  wire f_s_dadda_rca16_fa36_and0;
  wire f_s_dadda_rca16_fa36_xor1;
  wire f_s_dadda_rca16_fa36_and1;
  wire f_s_dadda_rca16_fa36_or0;
  wire f_s_dadda_rca16_ha10_xor0;
  wire f_s_dadda_rca16_ha10_and0;
  wire f_s_dadda_rca16_fa37_xor0;
  wire f_s_dadda_rca16_fa37_and0;
  wire f_s_dadda_rca16_fa37_xor1;
  wire f_s_dadda_rca16_fa37_and1;
  wire f_s_dadda_rca16_fa37_or0;
  wire f_s_dadda_rca16_fa38_xor0;
  wire f_s_dadda_rca16_fa38_and0;
  wire f_s_dadda_rca16_fa38_xor1;
  wire f_s_dadda_rca16_fa38_and1;
  wire f_s_dadda_rca16_fa38_or0;
  wire f_s_dadda_rca16_and_12_0;
  wire f_s_dadda_rca16_fa39_xor0;
  wire f_s_dadda_rca16_fa39_and0;
  wire f_s_dadda_rca16_fa39_xor1;
  wire f_s_dadda_rca16_fa39_and1;
  wire f_s_dadda_rca16_fa39_or0;
  wire f_s_dadda_rca16_and_11_1;
  wire f_s_dadda_rca16_and_10_2;
  wire f_s_dadda_rca16_and_9_3;
  wire f_s_dadda_rca16_fa40_xor0;
  wire f_s_dadda_rca16_fa40_and0;
  wire f_s_dadda_rca16_fa40_xor1;
  wire f_s_dadda_rca16_fa40_and1;
  wire f_s_dadda_rca16_fa40_or0;
  wire f_s_dadda_rca16_and_8_4;
  wire f_s_dadda_rca16_and_7_5;
  wire f_s_dadda_rca16_and_6_6;
  wire f_s_dadda_rca16_fa41_xor0;
  wire f_s_dadda_rca16_fa41_and0;
  wire f_s_dadda_rca16_fa41_xor1;
  wire f_s_dadda_rca16_fa41_and1;
  wire f_s_dadda_rca16_fa41_or0;
  wire f_s_dadda_rca16_and_5_7;
  wire f_s_dadda_rca16_and_4_8;
  wire f_s_dadda_rca16_and_3_9;
  wire f_s_dadda_rca16_fa42_xor0;
  wire f_s_dadda_rca16_fa42_and0;
  wire f_s_dadda_rca16_fa42_xor1;
  wire f_s_dadda_rca16_fa42_and1;
  wire f_s_dadda_rca16_fa42_or0;
  wire f_s_dadda_rca16_and_2_10;
  wire f_s_dadda_rca16_and_1_11;
  wire f_s_dadda_rca16_and_0_12;
  wire f_s_dadda_rca16_fa43_xor0;
  wire f_s_dadda_rca16_fa43_and0;
  wire f_s_dadda_rca16_fa43_xor1;
  wire f_s_dadda_rca16_fa43_and1;
  wire f_s_dadda_rca16_fa43_or0;
  wire f_s_dadda_rca16_fa44_xor0;
  wire f_s_dadda_rca16_fa44_and0;
  wire f_s_dadda_rca16_fa44_xor1;
  wire f_s_dadda_rca16_fa44_and1;
  wire f_s_dadda_rca16_fa44_or0;
  wire f_s_dadda_rca16_ha11_xor0;
  wire f_s_dadda_rca16_ha11_and0;
  wire f_s_dadda_rca16_fa45_xor0;
  wire f_s_dadda_rca16_fa45_and0;
  wire f_s_dadda_rca16_fa45_xor1;
  wire f_s_dadda_rca16_fa45_and1;
  wire f_s_dadda_rca16_fa45_or0;
  wire f_s_dadda_rca16_fa46_xor0;
  wire f_s_dadda_rca16_fa46_and0;
  wire f_s_dadda_rca16_fa46_xor1;
  wire f_s_dadda_rca16_fa46_and1;
  wire f_s_dadda_rca16_fa46_or0;
  wire f_s_dadda_rca16_fa47_xor0;
  wire f_s_dadda_rca16_fa47_and0;
  wire f_s_dadda_rca16_fa47_xor1;
  wire f_s_dadda_rca16_fa47_and1;
  wire f_s_dadda_rca16_fa47_or0;
  wire f_s_dadda_rca16_and_11_2;
  wire f_s_dadda_rca16_and_10_3;
  wire f_s_dadda_rca16_and_9_4;
  wire f_s_dadda_rca16_fa48_xor0;
  wire f_s_dadda_rca16_fa48_and0;
  wire f_s_dadda_rca16_fa48_xor1;
  wire f_s_dadda_rca16_fa48_and1;
  wire f_s_dadda_rca16_fa48_or0;
  wire f_s_dadda_rca16_and_8_5;
  wire f_s_dadda_rca16_and_7_6;
  wire f_s_dadda_rca16_and_6_7;
  wire f_s_dadda_rca16_fa49_xor0;
  wire f_s_dadda_rca16_fa49_and0;
  wire f_s_dadda_rca16_fa49_xor1;
  wire f_s_dadda_rca16_fa49_and1;
  wire f_s_dadda_rca16_fa49_or0;
  wire f_s_dadda_rca16_and_5_8;
  wire f_s_dadda_rca16_and_4_9;
  wire f_s_dadda_rca16_and_3_10;
  wire f_s_dadda_rca16_fa50_xor0;
  wire f_s_dadda_rca16_fa50_and0;
  wire f_s_dadda_rca16_fa50_xor1;
  wire f_s_dadda_rca16_fa50_and1;
  wire f_s_dadda_rca16_fa50_or0;
  wire f_s_dadda_rca16_and_2_11;
  wire f_s_dadda_rca16_and_1_12;
  wire f_s_dadda_rca16_and_0_13;
  wire f_s_dadda_rca16_fa51_xor0;
  wire f_s_dadda_rca16_fa51_and0;
  wire f_s_dadda_rca16_fa51_xor1;
  wire f_s_dadda_rca16_fa51_and1;
  wire f_s_dadda_rca16_fa51_or0;
  wire f_s_dadda_rca16_fa52_xor0;
  wire f_s_dadda_rca16_fa52_and0;
  wire f_s_dadda_rca16_fa52_xor1;
  wire f_s_dadda_rca16_fa52_and1;
  wire f_s_dadda_rca16_fa52_or0;
  wire f_s_dadda_rca16_fa53_xor0;
  wire f_s_dadda_rca16_fa53_and0;
  wire f_s_dadda_rca16_fa53_xor1;
  wire f_s_dadda_rca16_fa53_and1;
  wire f_s_dadda_rca16_fa53_or0;
  wire f_s_dadda_rca16_fa54_xor0;
  wire f_s_dadda_rca16_fa54_and0;
  wire f_s_dadda_rca16_fa54_xor1;
  wire f_s_dadda_rca16_fa54_and1;
  wire f_s_dadda_rca16_fa54_or0;
  wire f_s_dadda_rca16_fa55_xor0;
  wire f_s_dadda_rca16_fa55_and0;
  wire f_s_dadda_rca16_fa55_xor1;
  wire f_s_dadda_rca16_fa55_and1;
  wire f_s_dadda_rca16_fa55_or0;
  wire f_s_dadda_rca16_fa56_xor0;
  wire f_s_dadda_rca16_fa56_and0;
  wire f_s_dadda_rca16_fa56_xor1;
  wire f_s_dadda_rca16_fa56_and1;
  wire f_s_dadda_rca16_fa56_or0;
  wire f_s_dadda_rca16_and_10_4;
  wire f_s_dadda_rca16_and_9_5;
  wire f_s_dadda_rca16_and_8_6;
  wire f_s_dadda_rca16_fa57_xor0;
  wire f_s_dadda_rca16_fa57_and0;
  wire f_s_dadda_rca16_fa57_xor1;
  wire f_s_dadda_rca16_fa57_and1;
  wire f_s_dadda_rca16_fa57_or0;
  wire f_s_dadda_rca16_and_7_7;
  wire f_s_dadda_rca16_and_6_8;
  wire f_s_dadda_rca16_and_5_9;
  wire f_s_dadda_rca16_fa58_xor0;
  wire f_s_dadda_rca16_fa58_and0;
  wire f_s_dadda_rca16_fa58_xor1;
  wire f_s_dadda_rca16_fa58_and1;
  wire f_s_dadda_rca16_fa58_or0;
  wire f_s_dadda_rca16_and_4_10;
  wire f_s_dadda_rca16_and_3_11;
  wire f_s_dadda_rca16_and_2_12;
  wire f_s_dadda_rca16_fa59_xor0;
  wire f_s_dadda_rca16_fa59_and0;
  wire f_s_dadda_rca16_fa59_xor1;
  wire f_s_dadda_rca16_fa59_and1;
  wire f_s_dadda_rca16_fa59_or0;
  wire f_s_dadda_rca16_and_1_13;
  wire f_s_dadda_rca16_and_0_14;
  wire f_s_dadda_rca16_fa60_xor0;
  wire f_s_dadda_rca16_fa60_and0;
  wire f_s_dadda_rca16_fa60_xor1;
  wire f_s_dadda_rca16_fa60_and1;
  wire f_s_dadda_rca16_fa60_or0;
  wire f_s_dadda_rca16_fa61_xor0;
  wire f_s_dadda_rca16_fa61_and0;
  wire f_s_dadda_rca16_fa61_xor1;
  wire f_s_dadda_rca16_fa61_and1;
  wire f_s_dadda_rca16_fa61_or0;
  wire f_s_dadda_rca16_fa62_xor0;
  wire f_s_dadda_rca16_fa62_and0;
  wire f_s_dadda_rca16_fa62_xor1;
  wire f_s_dadda_rca16_fa62_and1;
  wire f_s_dadda_rca16_fa62_or0;
  wire f_s_dadda_rca16_fa63_xor0;
  wire f_s_dadda_rca16_fa63_and0;
  wire f_s_dadda_rca16_fa63_xor1;
  wire f_s_dadda_rca16_fa63_and1;
  wire f_s_dadda_rca16_fa63_or0;
  wire f_s_dadda_rca16_fa64_xor0;
  wire f_s_dadda_rca16_fa64_and0;
  wire f_s_dadda_rca16_fa64_xor1;
  wire f_s_dadda_rca16_fa64_and1;
  wire f_s_dadda_rca16_fa64_or0;
  wire f_s_dadda_rca16_fa65_xor0;
  wire f_s_dadda_rca16_fa65_and0;
  wire f_s_dadda_rca16_fa65_xor1;
  wire f_s_dadda_rca16_fa65_and1;
  wire f_s_dadda_rca16_fa65_or0;
  wire f_s_dadda_rca16_and_9_6;
  wire f_s_dadda_rca16_and_8_7;
  wire f_s_dadda_rca16_and_7_8;
  wire f_s_dadda_rca16_fa66_xor0;
  wire f_s_dadda_rca16_fa66_and0;
  wire f_s_dadda_rca16_fa66_xor1;
  wire f_s_dadda_rca16_fa66_and1;
  wire f_s_dadda_rca16_fa66_or0;
  wire f_s_dadda_rca16_and_6_9;
  wire f_s_dadda_rca16_and_5_10;
  wire f_s_dadda_rca16_and_4_11;
  wire f_s_dadda_rca16_fa67_xor0;
  wire f_s_dadda_rca16_fa67_and0;
  wire f_s_dadda_rca16_fa67_xor1;
  wire f_s_dadda_rca16_fa67_and1;
  wire f_s_dadda_rca16_fa67_or0;
  wire f_s_dadda_rca16_and_3_12;
  wire f_s_dadda_rca16_and_2_13;
  wire f_s_dadda_rca16_and_1_14;
  wire f_s_dadda_rca16_fa68_xor0;
  wire f_s_dadda_rca16_fa68_and0;
  wire f_s_dadda_rca16_fa68_xor1;
  wire f_s_dadda_rca16_fa68_and1;
  wire f_s_dadda_rca16_fa68_or0;
  wire f_s_dadda_rca16_nand_0_15;
  wire f_s_dadda_rca16_fa69_xor0;
  wire f_s_dadda_rca16_fa69_and0;
  wire f_s_dadda_rca16_fa69_xor1;
  wire f_s_dadda_rca16_fa69_and1;
  wire f_s_dadda_rca16_fa69_or0;
  wire f_s_dadda_rca16_fa70_xor0;
  wire f_s_dadda_rca16_fa70_and0;
  wire f_s_dadda_rca16_fa70_xor1;
  wire f_s_dadda_rca16_fa70_and1;
  wire f_s_dadda_rca16_fa70_or0;
  wire f_s_dadda_rca16_fa71_xor0;
  wire f_s_dadda_rca16_fa71_and0;
  wire f_s_dadda_rca16_fa71_xor1;
  wire f_s_dadda_rca16_fa71_and1;
  wire f_s_dadda_rca16_fa71_or0;
  wire f_s_dadda_rca16_fa72_xor0;
  wire f_s_dadda_rca16_fa72_and0;
  wire f_s_dadda_rca16_fa72_xor1;
  wire f_s_dadda_rca16_fa72_and1;
  wire f_s_dadda_rca16_fa72_or0;
  wire f_s_dadda_rca16_fa73_xor0;
  wire f_s_dadda_rca16_fa73_and0;
  wire f_s_dadda_rca16_fa73_xor1;
  wire f_s_dadda_rca16_fa73_and1;
  wire f_s_dadda_rca16_fa73_or0;
  wire f_s_dadda_rca16_fa74_xor0;
  wire f_s_dadda_rca16_fa74_and0;
  wire f_s_dadda_rca16_fa74_xor1;
  wire f_s_dadda_rca16_fa74_and1;
  wire f_s_dadda_rca16_fa74_or0;
  wire f_s_dadda_rca16_and_10_6;
  wire f_s_dadda_rca16_and_9_7;
  wire f_s_dadda_rca16_and_8_8;
  wire f_s_dadda_rca16_fa75_xor0;
  wire f_s_dadda_rca16_fa75_and0;
  wire f_s_dadda_rca16_fa75_xor1;
  wire f_s_dadda_rca16_fa75_and1;
  wire f_s_dadda_rca16_fa75_or0;
  wire f_s_dadda_rca16_and_7_9;
  wire f_s_dadda_rca16_and_6_10;
  wire f_s_dadda_rca16_and_5_11;
  wire f_s_dadda_rca16_fa76_xor0;
  wire f_s_dadda_rca16_fa76_and0;
  wire f_s_dadda_rca16_fa76_xor1;
  wire f_s_dadda_rca16_fa76_and1;
  wire f_s_dadda_rca16_fa76_or0;
  wire f_s_dadda_rca16_and_4_12;
  wire f_s_dadda_rca16_and_3_13;
  wire f_s_dadda_rca16_and_2_14;
  wire f_s_dadda_rca16_fa77_xor0;
  wire f_s_dadda_rca16_fa77_and0;
  wire f_s_dadda_rca16_fa77_xor1;
  wire f_s_dadda_rca16_fa77_and1;
  wire f_s_dadda_rca16_fa77_or0;
  wire f_s_dadda_rca16_nand_1_15;
  wire f_s_dadda_rca16_fa78_xor0;
  wire f_s_dadda_rca16_fa78_and0;
  wire f_s_dadda_rca16_fa78_xor1;
  wire f_s_dadda_rca16_fa78_and1;
  wire f_s_dadda_rca16_fa78_or0;
  wire f_s_dadda_rca16_fa79_xor0;
  wire f_s_dadda_rca16_fa79_and0;
  wire f_s_dadda_rca16_fa79_xor1;
  wire f_s_dadda_rca16_fa79_and1;
  wire f_s_dadda_rca16_fa79_or0;
  wire f_s_dadda_rca16_fa80_xor0;
  wire f_s_dadda_rca16_fa80_and0;
  wire f_s_dadda_rca16_fa80_xor1;
  wire f_s_dadda_rca16_fa80_and1;
  wire f_s_dadda_rca16_fa80_or0;
  wire f_s_dadda_rca16_fa81_xor0;
  wire f_s_dadda_rca16_fa81_and0;
  wire f_s_dadda_rca16_fa81_xor1;
  wire f_s_dadda_rca16_fa81_and1;
  wire f_s_dadda_rca16_fa81_or0;
  wire f_s_dadda_rca16_fa82_xor0;
  wire f_s_dadda_rca16_fa82_and0;
  wire f_s_dadda_rca16_fa82_xor1;
  wire f_s_dadda_rca16_fa82_and1;
  wire f_s_dadda_rca16_fa82_or0;
  wire f_s_dadda_rca16_fa83_xor0;
  wire f_s_dadda_rca16_fa83_and0;
  wire f_s_dadda_rca16_fa83_xor1;
  wire f_s_dadda_rca16_fa83_and1;
  wire f_s_dadda_rca16_fa83_or0;
  wire f_s_dadda_rca16_and_12_5;
  wire f_s_dadda_rca16_and_11_6;
  wire f_s_dadda_rca16_and_10_7;
  wire f_s_dadda_rca16_fa84_xor0;
  wire f_s_dadda_rca16_fa84_and0;
  wire f_s_dadda_rca16_fa84_xor1;
  wire f_s_dadda_rca16_fa84_and1;
  wire f_s_dadda_rca16_fa84_or0;
  wire f_s_dadda_rca16_and_9_8;
  wire f_s_dadda_rca16_and_8_9;
  wire f_s_dadda_rca16_and_7_10;
  wire f_s_dadda_rca16_fa85_xor0;
  wire f_s_dadda_rca16_fa85_and0;
  wire f_s_dadda_rca16_fa85_xor1;
  wire f_s_dadda_rca16_fa85_and1;
  wire f_s_dadda_rca16_fa85_or0;
  wire f_s_dadda_rca16_and_6_11;
  wire f_s_dadda_rca16_and_5_12;
  wire f_s_dadda_rca16_and_4_13;
  wire f_s_dadda_rca16_fa86_xor0;
  wire f_s_dadda_rca16_fa86_and0;
  wire f_s_dadda_rca16_fa86_xor1;
  wire f_s_dadda_rca16_fa86_and1;
  wire f_s_dadda_rca16_fa86_or0;
  wire f_s_dadda_rca16_and_3_14;
  wire f_s_dadda_rca16_nand_2_15;
  wire f_s_dadda_rca16_fa87_xor0;
  wire f_s_dadda_rca16_fa87_and0;
  wire f_s_dadda_rca16_fa87_xor1;
  wire f_s_dadda_rca16_fa87_and1;
  wire f_s_dadda_rca16_fa87_or0;
  wire f_s_dadda_rca16_fa88_xor0;
  wire f_s_dadda_rca16_fa88_and0;
  wire f_s_dadda_rca16_fa88_xor1;
  wire f_s_dadda_rca16_fa88_and1;
  wire f_s_dadda_rca16_fa88_or0;
  wire f_s_dadda_rca16_fa89_xor0;
  wire f_s_dadda_rca16_fa89_and0;
  wire f_s_dadda_rca16_fa89_xor1;
  wire f_s_dadda_rca16_fa89_and1;
  wire f_s_dadda_rca16_fa89_or0;
  wire f_s_dadda_rca16_fa90_xor0;
  wire f_s_dadda_rca16_fa90_and0;
  wire f_s_dadda_rca16_fa90_xor1;
  wire f_s_dadda_rca16_fa90_and1;
  wire f_s_dadda_rca16_fa90_or0;
  wire f_s_dadda_rca16_fa91_xor0;
  wire f_s_dadda_rca16_fa91_and0;
  wire f_s_dadda_rca16_fa91_xor1;
  wire f_s_dadda_rca16_fa91_and1;
  wire f_s_dadda_rca16_fa91_or0;
  wire f_s_dadda_rca16_fa92_xor0;
  wire f_s_dadda_rca16_fa92_and0;
  wire f_s_dadda_rca16_fa92_xor1;
  wire f_s_dadda_rca16_fa92_and1;
  wire f_s_dadda_rca16_fa92_or0;
  wire f_s_dadda_rca16_and_14_4;
  wire f_s_dadda_rca16_and_13_5;
  wire f_s_dadda_rca16_and_12_6;
  wire f_s_dadda_rca16_fa93_xor0;
  wire f_s_dadda_rca16_fa93_and0;
  wire f_s_dadda_rca16_fa93_xor1;
  wire f_s_dadda_rca16_fa93_and1;
  wire f_s_dadda_rca16_fa93_or0;
  wire f_s_dadda_rca16_and_11_7;
  wire f_s_dadda_rca16_and_10_8;
  wire f_s_dadda_rca16_and_9_9;
  wire f_s_dadda_rca16_fa94_xor0;
  wire f_s_dadda_rca16_fa94_and0;
  wire f_s_dadda_rca16_fa94_xor1;
  wire f_s_dadda_rca16_fa94_and1;
  wire f_s_dadda_rca16_fa94_or0;
  wire f_s_dadda_rca16_and_8_10;
  wire f_s_dadda_rca16_and_7_11;
  wire f_s_dadda_rca16_and_6_12;
  wire f_s_dadda_rca16_fa95_xor0;
  wire f_s_dadda_rca16_fa95_and0;
  wire f_s_dadda_rca16_fa95_xor1;
  wire f_s_dadda_rca16_fa95_and1;
  wire f_s_dadda_rca16_fa95_or0;
  wire f_s_dadda_rca16_and_5_13;
  wire f_s_dadda_rca16_and_4_14;
  wire f_s_dadda_rca16_nand_3_15;
  wire f_s_dadda_rca16_fa96_xor0;
  wire f_s_dadda_rca16_fa96_and0;
  wire f_s_dadda_rca16_fa96_xor1;
  wire f_s_dadda_rca16_fa96_and1;
  wire f_s_dadda_rca16_fa96_or0;
  wire f_s_dadda_rca16_fa97_xor0;
  wire f_s_dadda_rca16_fa97_and0;
  wire f_s_dadda_rca16_fa97_xor1;
  wire f_s_dadda_rca16_fa97_and1;
  wire f_s_dadda_rca16_fa97_or0;
  wire f_s_dadda_rca16_fa98_xor0;
  wire f_s_dadda_rca16_fa98_and0;
  wire f_s_dadda_rca16_fa98_xor1;
  wire f_s_dadda_rca16_fa98_and1;
  wire f_s_dadda_rca16_fa98_or0;
  wire f_s_dadda_rca16_fa99_xor0;
  wire f_s_dadda_rca16_fa99_and0;
  wire f_s_dadda_rca16_fa99_xor1;
  wire f_s_dadda_rca16_fa99_and1;
  wire f_s_dadda_rca16_fa99_or0;
  wire f_s_dadda_rca16_fa100_xor0;
  wire f_s_dadda_rca16_fa100_and0;
  wire f_s_dadda_rca16_fa100_xor1;
  wire f_s_dadda_rca16_fa100_and1;
  wire f_s_dadda_rca16_fa100_or0;
  wire f_s_dadda_rca16_fa101_xor0;
  wire f_s_dadda_rca16_fa101_and0;
  wire f_s_dadda_rca16_fa101_xor1;
  wire f_s_dadda_rca16_fa101_and1;
  wire f_s_dadda_rca16_fa101_or0;
  wire f_s_dadda_rca16_nand_15_4;
  wire f_s_dadda_rca16_and_14_5;
  wire f_s_dadda_rca16_fa102_xor0;
  wire f_s_dadda_rca16_fa102_and0;
  wire f_s_dadda_rca16_fa102_xor1;
  wire f_s_dadda_rca16_fa102_and1;
  wire f_s_dadda_rca16_fa102_or0;
  wire f_s_dadda_rca16_and_13_6;
  wire f_s_dadda_rca16_and_12_7;
  wire f_s_dadda_rca16_and_11_8;
  wire f_s_dadda_rca16_fa103_xor0;
  wire f_s_dadda_rca16_fa103_and0;
  wire f_s_dadda_rca16_fa103_xor1;
  wire f_s_dadda_rca16_fa103_and1;
  wire f_s_dadda_rca16_fa103_or0;
  wire f_s_dadda_rca16_and_10_9;
  wire f_s_dadda_rca16_and_9_10;
  wire f_s_dadda_rca16_and_8_11;
  wire f_s_dadda_rca16_fa104_xor0;
  wire f_s_dadda_rca16_fa104_and0;
  wire f_s_dadda_rca16_fa104_xor1;
  wire f_s_dadda_rca16_fa104_and1;
  wire f_s_dadda_rca16_fa104_or0;
  wire f_s_dadda_rca16_and_7_12;
  wire f_s_dadda_rca16_and_6_13;
  wire f_s_dadda_rca16_and_5_14;
  wire f_s_dadda_rca16_fa105_xor0;
  wire f_s_dadda_rca16_fa105_and0;
  wire f_s_dadda_rca16_fa105_xor1;
  wire f_s_dadda_rca16_fa105_and1;
  wire f_s_dadda_rca16_fa105_or0;
  wire f_s_dadda_rca16_nand_4_15;
  wire f_s_dadda_rca16_fa106_xor0;
  wire f_s_dadda_rca16_fa106_and0;
  wire f_s_dadda_rca16_fa106_xor1;
  wire f_s_dadda_rca16_fa106_and1;
  wire f_s_dadda_rca16_fa106_or0;
  wire f_s_dadda_rca16_fa107_xor0;
  wire f_s_dadda_rca16_fa107_and0;
  wire f_s_dadda_rca16_fa107_xor1;
  wire f_s_dadda_rca16_fa107_and1;
  wire f_s_dadda_rca16_fa107_or0;
  wire f_s_dadda_rca16_fa108_xor0;
  wire f_s_dadda_rca16_fa108_and0;
  wire f_s_dadda_rca16_fa108_xor1;
  wire f_s_dadda_rca16_fa108_and1;
  wire f_s_dadda_rca16_fa108_or0;
  wire f_s_dadda_rca16_fa109_xor0;
  wire f_s_dadda_rca16_fa109_and0;
  wire f_s_dadda_rca16_fa109_xor1;
  wire f_s_dadda_rca16_fa109_and1;
  wire f_s_dadda_rca16_fa109_or0;
  wire f_s_dadda_rca16_fa110_xor0;
  wire f_s_dadda_rca16_fa110_and0;
  wire f_s_dadda_rca16_fa110_xor1;
  wire f_s_dadda_rca16_fa110_and1;
  wire f_s_dadda_rca16_fa110_or0;
  wire f_s_dadda_rca16_nand_15_5;
  wire f_s_dadda_rca16_and_14_6;
  wire f_s_dadda_rca16_and_13_7;
  wire f_s_dadda_rca16_fa111_xor0;
  wire f_s_dadda_rca16_fa111_and0;
  wire f_s_dadda_rca16_fa111_xor1;
  wire f_s_dadda_rca16_fa111_and1;
  wire f_s_dadda_rca16_fa111_or0;
  wire f_s_dadda_rca16_and_12_8;
  wire f_s_dadda_rca16_and_11_9;
  wire f_s_dadda_rca16_and_10_10;
  wire f_s_dadda_rca16_fa112_xor0;
  wire f_s_dadda_rca16_fa112_and0;
  wire f_s_dadda_rca16_fa112_xor1;
  wire f_s_dadda_rca16_fa112_and1;
  wire f_s_dadda_rca16_fa112_or0;
  wire f_s_dadda_rca16_and_9_11;
  wire f_s_dadda_rca16_and_8_12;
  wire f_s_dadda_rca16_and_7_13;
  wire f_s_dadda_rca16_fa113_xor0;
  wire f_s_dadda_rca16_fa113_and0;
  wire f_s_dadda_rca16_fa113_xor1;
  wire f_s_dadda_rca16_fa113_and1;
  wire f_s_dadda_rca16_fa113_or0;
  wire f_s_dadda_rca16_and_6_14;
  wire f_s_dadda_rca16_nand_5_15;
  wire f_s_dadda_rca16_fa114_xor0;
  wire f_s_dadda_rca16_fa114_and0;
  wire f_s_dadda_rca16_fa114_xor1;
  wire f_s_dadda_rca16_fa114_and1;
  wire f_s_dadda_rca16_fa114_or0;
  wire f_s_dadda_rca16_fa115_xor0;
  wire f_s_dadda_rca16_fa115_and0;
  wire f_s_dadda_rca16_fa115_xor1;
  wire f_s_dadda_rca16_fa115_and1;
  wire f_s_dadda_rca16_fa115_or0;
  wire f_s_dadda_rca16_fa116_xor0;
  wire f_s_dadda_rca16_fa116_and0;
  wire f_s_dadda_rca16_fa116_xor1;
  wire f_s_dadda_rca16_fa116_and1;
  wire f_s_dadda_rca16_fa116_or0;
  wire f_s_dadda_rca16_fa117_xor0;
  wire f_s_dadda_rca16_fa117_and0;
  wire f_s_dadda_rca16_fa117_xor1;
  wire f_s_dadda_rca16_fa117_and1;
  wire f_s_dadda_rca16_fa117_or0;
  wire f_s_dadda_rca16_nand_15_6;
  wire f_s_dadda_rca16_fa118_xor0;
  wire f_s_dadda_rca16_fa118_and0;
  wire f_s_dadda_rca16_fa118_xor1;
  wire f_s_dadda_rca16_fa118_and1;
  wire f_s_dadda_rca16_fa118_or0;
  wire f_s_dadda_rca16_and_14_7;
  wire f_s_dadda_rca16_and_13_8;
  wire f_s_dadda_rca16_and_12_9;
  wire f_s_dadda_rca16_fa119_xor0;
  wire f_s_dadda_rca16_fa119_and0;
  wire f_s_dadda_rca16_fa119_xor1;
  wire f_s_dadda_rca16_fa119_and1;
  wire f_s_dadda_rca16_fa119_or0;
  wire f_s_dadda_rca16_and_11_10;
  wire f_s_dadda_rca16_and_10_11;
  wire f_s_dadda_rca16_and_9_12;
  wire f_s_dadda_rca16_fa120_xor0;
  wire f_s_dadda_rca16_fa120_and0;
  wire f_s_dadda_rca16_fa120_xor1;
  wire f_s_dadda_rca16_fa120_and1;
  wire f_s_dadda_rca16_fa120_or0;
  wire f_s_dadda_rca16_and_8_13;
  wire f_s_dadda_rca16_and_7_14;
  wire f_s_dadda_rca16_nand_6_15;
  wire f_s_dadda_rca16_fa121_xor0;
  wire f_s_dadda_rca16_fa121_and0;
  wire f_s_dadda_rca16_fa121_xor1;
  wire f_s_dadda_rca16_fa121_and1;
  wire f_s_dadda_rca16_fa121_or0;
  wire f_s_dadda_rca16_fa122_xor0;
  wire f_s_dadda_rca16_fa122_and0;
  wire f_s_dadda_rca16_fa122_xor1;
  wire f_s_dadda_rca16_fa122_and1;
  wire f_s_dadda_rca16_fa122_or0;
  wire f_s_dadda_rca16_fa123_xor0;
  wire f_s_dadda_rca16_fa123_and0;
  wire f_s_dadda_rca16_fa123_xor1;
  wire f_s_dadda_rca16_fa123_and1;
  wire f_s_dadda_rca16_fa123_or0;
  wire f_s_dadda_rca16_fa124_xor0;
  wire f_s_dadda_rca16_fa124_and0;
  wire f_s_dadda_rca16_fa124_xor1;
  wire f_s_dadda_rca16_fa124_and1;
  wire f_s_dadda_rca16_fa124_or0;
  wire f_s_dadda_rca16_nand_15_7;
  wire f_s_dadda_rca16_and_14_8;
  wire f_s_dadda_rca16_fa125_xor0;
  wire f_s_dadda_rca16_fa125_and0;
  wire f_s_dadda_rca16_fa125_xor1;
  wire f_s_dadda_rca16_fa125_and1;
  wire f_s_dadda_rca16_fa125_or0;
  wire f_s_dadda_rca16_and_13_9;
  wire f_s_dadda_rca16_and_12_10;
  wire f_s_dadda_rca16_and_11_11;
  wire f_s_dadda_rca16_fa126_xor0;
  wire f_s_dadda_rca16_fa126_and0;
  wire f_s_dadda_rca16_fa126_xor1;
  wire f_s_dadda_rca16_fa126_and1;
  wire f_s_dadda_rca16_fa126_or0;
  wire f_s_dadda_rca16_and_10_12;
  wire f_s_dadda_rca16_and_9_13;
  wire f_s_dadda_rca16_and_8_14;
  wire f_s_dadda_rca16_fa127_xor0;
  wire f_s_dadda_rca16_fa127_and0;
  wire f_s_dadda_rca16_fa127_xor1;
  wire f_s_dadda_rca16_fa127_and1;
  wire f_s_dadda_rca16_fa127_or0;
  wire f_s_dadda_rca16_nand_7_15;
  wire f_s_dadda_rca16_fa128_xor0;
  wire f_s_dadda_rca16_fa128_and0;
  wire f_s_dadda_rca16_fa128_xor1;
  wire f_s_dadda_rca16_fa128_and1;
  wire f_s_dadda_rca16_fa128_or0;
  wire f_s_dadda_rca16_fa129_xor0;
  wire f_s_dadda_rca16_fa129_and0;
  wire f_s_dadda_rca16_fa129_xor1;
  wire f_s_dadda_rca16_fa129_and1;
  wire f_s_dadda_rca16_fa129_or0;
  wire f_s_dadda_rca16_fa130_xor0;
  wire f_s_dadda_rca16_fa130_and0;
  wire f_s_dadda_rca16_fa130_xor1;
  wire f_s_dadda_rca16_fa130_and1;
  wire f_s_dadda_rca16_fa130_or0;
  wire f_s_dadda_rca16_nand_15_8;
  wire f_s_dadda_rca16_and_14_9;
  wire f_s_dadda_rca16_and_13_10;
  wire f_s_dadda_rca16_fa131_xor0;
  wire f_s_dadda_rca16_fa131_and0;
  wire f_s_dadda_rca16_fa131_xor1;
  wire f_s_dadda_rca16_fa131_and1;
  wire f_s_dadda_rca16_fa131_or0;
  wire f_s_dadda_rca16_and_12_11;
  wire f_s_dadda_rca16_and_11_12;
  wire f_s_dadda_rca16_and_10_13;
  wire f_s_dadda_rca16_fa132_xor0;
  wire f_s_dadda_rca16_fa132_and0;
  wire f_s_dadda_rca16_fa132_xor1;
  wire f_s_dadda_rca16_fa132_and1;
  wire f_s_dadda_rca16_fa132_or0;
  wire f_s_dadda_rca16_and_9_14;
  wire f_s_dadda_rca16_nand_8_15;
  wire f_s_dadda_rca16_fa133_xor0;
  wire f_s_dadda_rca16_fa133_and0;
  wire f_s_dadda_rca16_fa133_xor1;
  wire f_s_dadda_rca16_fa133_and1;
  wire f_s_dadda_rca16_fa133_or0;
  wire f_s_dadda_rca16_fa134_xor0;
  wire f_s_dadda_rca16_fa134_and0;
  wire f_s_dadda_rca16_fa134_xor1;
  wire f_s_dadda_rca16_fa134_and1;
  wire f_s_dadda_rca16_fa134_or0;
  wire f_s_dadda_rca16_nand_15_9;
  wire f_s_dadda_rca16_fa135_xor0;
  wire f_s_dadda_rca16_fa135_and0;
  wire f_s_dadda_rca16_fa135_xor1;
  wire f_s_dadda_rca16_fa135_and1;
  wire f_s_dadda_rca16_fa135_or0;
  wire f_s_dadda_rca16_and_14_10;
  wire f_s_dadda_rca16_and_13_11;
  wire f_s_dadda_rca16_and_12_12;
  wire f_s_dadda_rca16_fa136_xor0;
  wire f_s_dadda_rca16_fa136_and0;
  wire f_s_dadda_rca16_fa136_xor1;
  wire f_s_dadda_rca16_fa136_and1;
  wire f_s_dadda_rca16_fa136_or0;
  wire f_s_dadda_rca16_and_11_13;
  wire f_s_dadda_rca16_and_10_14;
  wire f_s_dadda_rca16_nand_9_15;
  wire f_s_dadda_rca16_fa137_xor0;
  wire f_s_dadda_rca16_fa137_and0;
  wire f_s_dadda_rca16_fa137_xor1;
  wire f_s_dadda_rca16_fa137_and1;
  wire f_s_dadda_rca16_fa137_or0;
  wire f_s_dadda_rca16_fa138_xor0;
  wire f_s_dadda_rca16_fa138_and0;
  wire f_s_dadda_rca16_fa138_xor1;
  wire f_s_dadda_rca16_fa138_and1;
  wire f_s_dadda_rca16_fa138_or0;
  wire f_s_dadda_rca16_nand_15_10;
  wire f_s_dadda_rca16_and_14_11;
  wire f_s_dadda_rca16_fa139_xor0;
  wire f_s_dadda_rca16_fa139_and0;
  wire f_s_dadda_rca16_fa139_xor1;
  wire f_s_dadda_rca16_fa139_and1;
  wire f_s_dadda_rca16_fa139_or0;
  wire f_s_dadda_rca16_and_13_12;
  wire f_s_dadda_rca16_and_12_13;
  wire f_s_dadda_rca16_and_11_14;
  wire f_s_dadda_rca16_fa140_xor0;
  wire f_s_dadda_rca16_fa140_and0;
  wire f_s_dadda_rca16_fa140_xor1;
  wire f_s_dadda_rca16_fa140_and1;
  wire f_s_dadda_rca16_fa140_or0;
  wire f_s_dadda_rca16_fa141_xor0;
  wire f_s_dadda_rca16_fa141_and0;
  wire f_s_dadda_rca16_fa141_xor1;
  wire f_s_dadda_rca16_fa141_and1;
  wire f_s_dadda_rca16_fa141_or0;
  wire f_s_dadda_rca16_nand_15_11;
  wire f_s_dadda_rca16_and_14_12;
  wire f_s_dadda_rca16_and_13_13;
  wire f_s_dadda_rca16_fa142_xor0;
  wire f_s_dadda_rca16_fa142_and0;
  wire f_s_dadda_rca16_fa142_xor1;
  wire f_s_dadda_rca16_fa142_and1;
  wire f_s_dadda_rca16_fa142_or0;
  wire f_s_dadda_rca16_nand_15_12;
  wire f_s_dadda_rca16_fa143_xor0;
  wire f_s_dadda_rca16_fa143_and0;
  wire f_s_dadda_rca16_fa143_xor1;
  wire f_s_dadda_rca16_fa143_and1;
  wire f_s_dadda_rca16_fa143_or0;
  wire f_s_dadda_rca16_and_3_0;
  wire f_s_dadda_rca16_and_2_1;
  wire f_s_dadda_rca16_ha12_xor0;
  wire f_s_dadda_rca16_ha12_and0;
  wire f_s_dadda_rca16_and_2_2;
  wire f_s_dadda_rca16_and_1_3;
  wire f_s_dadda_rca16_fa144_xor0;
  wire f_s_dadda_rca16_fa144_and0;
  wire f_s_dadda_rca16_fa144_xor1;
  wire f_s_dadda_rca16_fa144_and1;
  wire f_s_dadda_rca16_fa144_or0;
  wire f_s_dadda_rca16_and_1_4;
  wire f_s_dadda_rca16_and_0_5;
  wire f_s_dadda_rca16_fa145_xor0;
  wire f_s_dadda_rca16_fa145_and0;
  wire f_s_dadda_rca16_fa145_xor1;
  wire f_s_dadda_rca16_fa145_and1;
  wire f_s_dadda_rca16_fa145_or0;
  wire f_s_dadda_rca16_and_0_6;
  wire f_s_dadda_rca16_fa146_xor0;
  wire f_s_dadda_rca16_fa146_and0;
  wire f_s_dadda_rca16_fa146_xor1;
  wire f_s_dadda_rca16_fa146_and1;
  wire f_s_dadda_rca16_fa146_or0;
  wire f_s_dadda_rca16_fa147_xor0;
  wire f_s_dadda_rca16_fa147_and0;
  wire f_s_dadda_rca16_fa147_xor1;
  wire f_s_dadda_rca16_fa147_and1;
  wire f_s_dadda_rca16_fa147_or0;
  wire f_s_dadda_rca16_fa148_xor0;
  wire f_s_dadda_rca16_fa148_and0;
  wire f_s_dadda_rca16_fa148_xor1;
  wire f_s_dadda_rca16_fa148_and1;
  wire f_s_dadda_rca16_fa148_or0;
  wire f_s_dadda_rca16_fa149_xor0;
  wire f_s_dadda_rca16_fa149_and0;
  wire f_s_dadda_rca16_fa149_xor1;
  wire f_s_dadda_rca16_fa149_and1;
  wire f_s_dadda_rca16_fa149_or0;
  wire f_s_dadda_rca16_fa150_xor0;
  wire f_s_dadda_rca16_fa150_and0;
  wire f_s_dadda_rca16_fa150_xor1;
  wire f_s_dadda_rca16_fa150_and1;
  wire f_s_dadda_rca16_fa150_or0;
  wire f_s_dadda_rca16_fa151_xor0;
  wire f_s_dadda_rca16_fa151_and0;
  wire f_s_dadda_rca16_fa151_xor1;
  wire f_s_dadda_rca16_fa151_and1;
  wire f_s_dadda_rca16_fa151_or0;
  wire f_s_dadda_rca16_fa152_xor0;
  wire f_s_dadda_rca16_fa152_and0;
  wire f_s_dadda_rca16_fa152_xor1;
  wire f_s_dadda_rca16_fa152_and1;
  wire f_s_dadda_rca16_fa152_or0;
  wire f_s_dadda_rca16_fa153_xor0;
  wire f_s_dadda_rca16_fa153_and0;
  wire f_s_dadda_rca16_fa153_xor1;
  wire f_s_dadda_rca16_fa153_and1;
  wire f_s_dadda_rca16_fa153_or0;
  wire f_s_dadda_rca16_fa154_xor0;
  wire f_s_dadda_rca16_fa154_and0;
  wire f_s_dadda_rca16_fa154_xor1;
  wire f_s_dadda_rca16_fa154_and1;
  wire f_s_dadda_rca16_fa154_or0;
  wire f_s_dadda_rca16_fa155_xor0;
  wire f_s_dadda_rca16_fa155_and0;
  wire f_s_dadda_rca16_fa155_xor1;
  wire f_s_dadda_rca16_fa155_and1;
  wire f_s_dadda_rca16_fa155_or0;
  wire f_s_dadda_rca16_fa156_xor0;
  wire f_s_dadda_rca16_fa156_and0;
  wire f_s_dadda_rca16_fa156_xor1;
  wire f_s_dadda_rca16_fa156_and1;
  wire f_s_dadda_rca16_fa156_or0;
  wire f_s_dadda_rca16_fa157_xor0;
  wire f_s_dadda_rca16_fa157_and0;
  wire f_s_dadda_rca16_fa157_xor1;
  wire f_s_dadda_rca16_fa157_and1;
  wire f_s_dadda_rca16_fa157_or0;
  wire f_s_dadda_rca16_fa158_xor0;
  wire f_s_dadda_rca16_fa158_and0;
  wire f_s_dadda_rca16_fa158_xor1;
  wire f_s_dadda_rca16_fa158_and1;
  wire f_s_dadda_rca16_fa158_or0;
  wire f_s_dadda_rca16_fa159_xor0;
  wire f_s_dadda_rca16_fa159_and0;
  wire f_s_dadda_rca16_fa159_xor1;
  wire f_s_dadda_rca16_fa159_and1;
  wire f_s_dadda_rca16_fa159_or0;
  wire f_s_dadda_rca16_fa160_xor0;
  wire f_s_dadda_rca16_fa160_and0;
  wire f_s_dadda_rca16_fa160_xor1;
  wire f_s_dadda_rca16_fa160_and1;
  wire f_s_dadda_rca16_fa160_or0;
  wire f_s_dadda_rca16_fa161_xor0;
  wire f_s_dadda_rca16_fa161_and0;
  wire f_s_dadda_rca16_fa161_xor1;
  wire f_s_dadda_rca16_fa161_and1;
  wire f_s_dadda_rca16_fa161_or0;
  wire f_s_dadda_rca16_fa162_xor0;
  wire f_s_dadda_rca16_fa162_and0;
  wire f_s_dadda_rca16_fa162_xor1;
  wire f_s_dadda_rca16_fa162_and1;
  wire f_s_dadda_rca16_fa162_or0;
  wire f_s_dadda_rca16_fa163_xor0;
  wire f_s_dadda_rca16_fa163_and0;
  wire f_s_dadda_rca16_fa163_xor1;
  wire f_s_dadda_rca16_fa163_and1;
  wire f_s_dadda_rca16_fa163_or0;
  wire f_s_dadda_rca16_fa164_xor0;
  wire f_s_dadda_rca16_fa164_and0;
  wire f_s_dadda_rca16_fa164_xor1;
  wire f_s_dadda_rca16_fa164_and1;
  wire f_s_dadda_rca16_fa164_or0;
  wire f_s_dadda_rca16_nand_10_15;
  wire f_s_dadda_rca16_fa165_xor0;
  wire f_s_dadda_rca16_fa165_and0;
  wire f_s_dadda_rca16_fa165_xor1;
  wire f_s_dadda_rca16_fa165_and1;
  wire f_s_dadda_rca16_fa165_or0;
  wire f_s_dadda_rca16_and_12_14;
  wire f_s_dadda_rca16_nand_11_15;
  wire f_s_dadda_rca16_fa166_xor0;
  wire f_s_dadda_rca16_fa166_and0;
  wire f_s_dadda_rca16_fa166_xor1;
  wire f_s_dadda_rca16_fa166_and1;
  wire f_s_dadda_rca16_fa166_or0;
  wire f_s_dadda_rca16_and_14_13;
  wire f_s_dadda_rca16_and_13_14;
  wire f_s_dadda_rca16_fa167_xor0;
  wire f_s_dadda_rca16_fa167_and0;
  wire f_s_dadda_rca16_fa167_xor1;
  wire f_s_dadda_rca16_fa167_and1;
  wire f_s_dadda_rca16_fa167_or0;
  wire f_s_dadda_rca16_nand_15_13;
  wire f_s_dadda_rca16_fa168_xor0;
  wire f_s_dadda_rca16_fa168_and0;
  wire f_s_dadda_rca16_fa168_xor1;
  wire f_s_dadda_rca16_fa168_and1;
  wire f_s_dadda_rca16_fa168_or0;
  wire f_s_dadda_rca16_and_2_0;
  wire f_s_dadda_rca16_and_1_1;
  wire f_s_dadda_rca16_ha13_xor0;
  wire f_s_dadda_rca16_ha13_and0;
  wire f_s_dadda_rca16_and_1_2;
  wire f_s_dadda_rca16_and_0_3;
  wire f_s_dadda_rca16_fa169_xor0;
  wire f_s_dadda_rca16_fa169_and0;
  wire f_s_dadda_rca16_fa169_xor1;
  wire f_s_dadda_rca16_fa169_and1;
  wire f_s_dadda_rca16_fa169_or0;
  wire f_s_dadda_rca16_and_0_4;
  wire f_s_dadda_rca16_fa170_xor0;
  wire f_s_dadda_rca16_fa170_and0;
  wire f_s_dadda_rca16_fa170_xor1;
  wire f_s_dadda_rca16_fa170_and1;
  wire f_s_dadda_rca16_fa170_or0;
  wire f_s_dadda_rca16_fa171_xor0;
  wire f_s_dadda_rca16_fa171_and0;
  wire f_s_dadda_rca16_fa171_xor1;
  wire f_s_dadda_rca16_fa171_and1;
  wire f_s_dadda_rca16_fa171_or0;
  wire f_s_dadda_rca16_fa172_xor0;
  wire f_s_dadda_rca16_fa172_and0;
  wire f_s_dadda_rca16_fa172_xor1;
  wire f_s_dadda_rca16_fa172_and1;
  wire f_s_dadda_rca16_fa172_or0;
  wire f_s_dadda_rca16_fa173_xor0;
  wire f_s_dadda_rca16_fa173_and0;
  wire f_s_dadda_rca16_fa173_xor1;
  wire f_s_dadda_rca16_fa173_and1;
  wire f_s_dadda_rca16_fa173_or0;
  wire f_s_dadda_rca16_fa174_xor0;
  wire f_s_dadda_rca16_fa174_and0;
  wire f_s_dadda_rca16_fa174_xor1;
  wire f_s_dadda_rca16_fa174_and1;
  wire f_s_dadda_rca16_fa174_or0;
  wire f_s_dadda_rca16_fa175_xor0;
  wire f_s_dadda_rca16_fa175_and0;
  wire f_s_dadda_rca16_fa175_xor1;
  wire f_s_dadda_rca16_fa175_and1;
  wire f_s_dadda_rca16_fa175_or0;
  wire f_s_dadda_rca16_fa176_xor0;
  wire f_s_dadda_rca16_fa176_and0;
  wire f_s_dadda_rca16_fa176_xor1;
  wire f_s_dadda_rca16_fa176_and1;
  wire f_s_dadda_rca16_fa176_or0;
  wire f_s_dadda_rca16_fa177_xor0;
  wire f_s_dadda_rca16_fa177_and0;
  wire f_s_dadda_rca16_fa177_xor1;
  wire f_s_dadda_rca16_fa177_and1;
  wire f_s_dadda_rca16_fa177_or0;
  wire f_s_dadda_rca16_fa178_xor0;
  wire f_s_dadda_rca16_fa178_and0;
  wire f_s_dadda_rca16_fa178_xor1;
  wire f_s_dadda_rca16_fa178_and1;
  wire f_s_dadda_rca16_fa178_or0;
  wire f_s_dadda_rca16_fa179_xor0;
  wire f_s_dadda_rca16_fa179_and0;
  wire f_s_dadda_rca16_fa179_xor1;
  wire f_s_dadda_rca16_fa179_and1;
  wire f_s_dadda_rca16_fa179_or0;
  wire f_s_dadda_rca16_fa180_xor0;
  wire f_s_dadda_rca16_fa180_and0;
  wire f_s_dadda_rca16_fa180_xor1;
  wire f_s_dadda_rca16_fa180_and1;
  wire f_s_dadda_rca16_fa180_or0;
  wire f_s_dadda_rca16_fa181_xor0;
  wire f_s_dadda_rca16_fa181_and0;
  wire f_s_dadda_rca16_fa181_xor1;
  wire f_s_dadda_rca16_fa181_and1;
  wire f_s_dadda_rca16_fa181_or0;
  wire f_s_dadda_rca16_fa182_xor0;
  wire f_s_dadda_rca16_fa182_and0;
  wire f_s_dadda_rca16_fa182_xor1;
  wire f_s_dadda_rca16_fa182_and1;
  wire f_s_dadda_rca16_fa182_or0;
  wire f_s_dadda_rca16_fa183_xor0;
  wire f_s_dadda_rca16_fa183_and0;
  wire f_s_dadda_rca16_fa183_xor1;
  wire f_s_dadda_rca16_fa183_and1;
  wire f_s_dadda_rca16_fa183_or0;
  wire f_s_dadda_rca16_fa184_xor0;
  wire f_s_dadda_rca16_fa184_and0;
  wire f_s_dadda_rca16_fa184_xor1;
  wire f_s_dadda_rca16_fa184_and1;
  wire f_s_dadda_rca16_fa184_or0;
  wire f_s_dadda_rca16_fa185_xor0;
  wire f_s_dadda_rca16_fa185_and0;
  wire f_s_dadda_rca16_fa185_xor1;
  wire f_s_dadda_rca16_fa185_and1;
  wire f_s_dadda_rca16_fa185_or0;
  wire f_s_dadda_rca16_fa186_xor0;
  wire f_s_dadda_rca16_fa186_and0;
  wire f_s_dadda_rca16_fa186_xor1;
  wire f_s_dadda_rca16_fa186_and1;
  wire f_s_dadda_rca16_fa186_or0;
  wire f_s_dadda_rca16_fa187_xor0;
  wire f_s_dadda_rca16_fa187_and0;
  wire f_s_dadda_rca16_fa187_xor1;
  wire f_s_dadda_rca16_fa187_and1;
  wire f_s_dadda_rca16_fa187_or0;
  wire f_s_dadda_rca16_fa188_xor0;
  wire f_s_dadda_rca16_fa188_and0;
  wire f_s_dadda_rca16_fa188_xor1;
  wire f_s_dadda_rca16_fa188_and1;
  wire f_s_dadda_rca16_fa188_or0;
  wire f_s_dadda_rca16_fa189_xor0;
  wire f_s_dadda_rca16_fa189_and0;
  wire f_s_dadda_rca16_fa189_xor1;
  wire f_s_dadda_rca16_fa189_and1;
  wire f_s_dadda_rca16_fa189_or0;
  wire f_s_dadda_rca16_fa190_xor0;
  wire f_s_dadda_rca16_fa190_and0;
  wire f_s_dadda_rca16_fa190_xor1;
  wire f_s_dadda_rca16_fa190_and1;
  wire f_s_dadda_rca16_fa190_or0;
  wire f_s_dadda_rca16_fa191_xor0;
  wire f_s_dadda_rca16_fa191_and0;
  wire f_s_dadda_rca16_fa191_xor1;
  wire f_s_dadda_rca16_fa191_and1;
  wire f_s_dadda_rca16_fa191_or0;
  wire f_s_dadda_rca16_fa192_xor0;
  wire f_s_dadda_rca16_fa192_and0;
  wire f_s_dadda_rca16_fa192_xor1;
  wire f_s_dadda_rca16_fa192_and1;
  wire f_s_dadda_rca16_fa192_or0;
  wire f_s_dadda_rca16_nand_12_15;
  wire f_s_dadda_rca16_fa193_xor0;
  wire f_s_dadda_rca16_fa193_and0;
  wire f_s_dadda_rca16_fa193_xor1;
  wire f_s_dadda_rca16_fa193_and1;
  wire f_s_dadda_rca16_fa193_or0;
  wire f_s_dadda_rca16_and_14_14;
  wire f_s_dadda_rca16_nand_13_15;
  wire f_s_dadda_rca16_fa194_xor0;
  wire f_s_dadda_rca16_fa194_and0;
  wire f_s_dadda_rca16_fa194_xor1;
  wire f_s_dadda_rca16_fa194_and1;
  wire f_s_dadda_rca16_fa194_or0;
  wire f_s_dadda_rca16_nand_15_14;
  wire f_s_dadda_rca16_fa195_xor0;
  wire f_s_dadda_rca16_fa195_and0;
  wire f_s_dadda_rca16_fa195_xor1;
  wire f_s_dadda_rca16_fa195_and1;
  wire f_s_dadda_rca16_fa195_or0;
  wire f_s_dadda_rca16_and_0_0;
  wire f_s_dadda_rca16_and_1_0;
  wire f_s_dadda_rca16_and_0_2;
  wire f_s_dadda_rca16_nand_14_15;
  wire f_s_dadda_rca16_and_0_1;
  wire f_s_dadda_rca16_and_15_15;
  wire f_s_dadda_rca16_u_rca30_ha_xor0;
  wire f_s_dadda_rca16_u_rca30_ha_and0;
  wire f_s_dadda_rca16_u_rca30_fa1_xor0;
  wire f_s_dadda_rca16_u_rca30_fa1_and0;
  wire f_s_dadda_rca16_u_rca30_fa1_xor1;
  wire f_s_dadda_rca16_u_rca30_fa1_and1;
  wire f_s_dadda_rca16_u_rca30_fa1_or0;
  wire f_s_dadda_rca16_u_rca30_fa2_xor0;
  wire f_s_dadda_rca16_u_rca30_fa2_and0;
  wire f_s_dadda_rca16_u_rca30_fa2_xor1;
  wire f_s_dadda_rca16_u_rca30_fa2_and1;
  wire f_s_dadda_rca16_u_rca30_fa2_or0;
  wire f_s_dadda_rca16_u_rca30_fa3_xor0;
  wire f_s_dadda_rca16_u_rca30_fa3_and0;
  wire f_s_dadda_rca16_u_rca30_fa3_xor1;
  wire f_s_dadda_rca16_u_rca30_fa3_and1;
  wire f_s_dadda_rca16_u_rca30_fa3_or0;
  wire f_s_dadda_rca16_u_rca30_fa4_xor0;
  wire f_s_dadda_rca16_u_rca30_fa4_and0;
  wire f_s_dadda_rca16_u_rca30_fa4_xor1;
  wire f_s_dadda_rca16_u_rca30_fa4_and1;
  wire f_s_dadda_rca16_u_rca30_fa4_or0;
  wire f_s_dadda_rca16_u_rca30_fa5_xor0;
  wire f_s_dadda_rca16_u_rca30_fa5_and0;
  wire f_s_dadda_rca16_u_rca30_fa5_xor1;
  wire f_s_dadda_rca16_u_rca30_fa5_and1;
  wire f_s_dadda_rca16_u_rca30_fa5_or0;
  wire f_s_dadda_rca16_u_rca30_fa6_xor0;
  wire f_s_dadda_rca16_u_rca30_fa6_and0;
  wire f_s_dadda_rca16_u_rca30_fa6_xor1;
  wire f_s_dadda_rca16_u_rca30_fa6_and1;
  wire f_s_dadda_rca16_u_rca30_fa6_or0;
  wire f_s_dadda_rca16_u_rca30_fa7_xor0;
  wire f_s_dadda_rca16_u_rca30_fa7_and0;
  wire f_s_dadda_rca16_u_rca30_fa7_xor1;
  wire f_s_dadda_rca16_u_rca30_fa7_and1;
  wire f_s_dadda_rca16_u_rca30_fa7_or0;
  wire f_s_dadda_rca16_u_rca30_fa8_xor0;
  wire f_s_dadda_rca16_u_rca30_fa8_and0;
  wire f_s_dadda_rca16_u_rca30_fa8_xor1;
  wire f_s_dadda_rca16_u_rca30_fa8_and1;
  wire f_s_dadda_rca16_u_rca30_fa8_or0;
  wire f_s_dadda_rca16_u_rca30_fa9_xor0;
  wire f_s_dadda_rca16_u_rca30_fa9_and0;
  wire f_s_dadda_rca16_u_rca30_fa9_xor1;
  wire f_s_dadda_rca16_u_rca30_fa9_and1;
  wire f_s_dadda_rca16_u_rca30_fa9_or0;
  wire f_s_dadda_rca16_u_rca30_fa10_xor0;
  wire f_s_dadda_rca16_u_rca30_fa10_and0;
  wire f_s_dadda_rca16_u_rca30_fa10_xor1;
  wire f_s_dadda_rca16_u_rca30_fa10_and1;
  wire f_s_dadda_rca16_u_rca30_fa10_or0;
  wire f_s_dadda_rca16_u_rca30_fa11_xor0;
  wire f_s_dadda_rca16_u_rca30_fa11_and0;
  wire f_s_dadda_rca16_u_rca30_fa11_xor1;
  wire f_s_dadda_rca16_u_rca30_fa11_and1;
  wire f_s_dadda_rca16_u_rca30_fa11_or0;
  wire f_s_dadda_rca16_u_rca30_fa12_xor0;
  wire f_s_dadda_rca16_u_rca30_fa12_and0;
  wire f_s_dadda_rca16_u_rca30_fa12_xor1;
  wire f_s_dadda_rca16_u_rca30_fa12_and1;
  wire f_s_dadda_rca16_u_rca30_fa12_or0;
  wire f_s_dadda_rca16_u_rca30_fa13_xor0;
  wire f_s_dadda_rca16_u_rca30_fa13_and0;
  wire f_s_dadda_rca16_u_rca30_fa13_xor1;
  wire f_s_dadda_rca16_u_rca30_fa13_and1;
  wire f_s_dadda_rca16_u_rca30_fa13_or0;
  wire f_s_dadda_rca16_u_rca30_fa14_xor0;
  wire f_s_dadda_rca16_u_rca30_fa14_and0;
  wire f_s_dadda_rca16_u_rca30_fa14_xor1;
  wire f_s_dadda_rca16_u_rca30_fa14_and1;
  wire f_s_dadda_rca16_u_rca30_fa14_or0;
  wire f_s_dadda_rca16_u_rca30_fa15_xor0;
  wire f_s_dadda_rca16_u_rca30_fa15_and0;
  wire f_s_dadda_rca16_u_rca30_fa15_xor1;
  wire f_s_dadda_rca16_u_rca30_fa15_and1;
  wire f_s_dadda_rca16_u_rca30_fa15_or0;
  wire f_s_dadda_rca16_u_rca30_fa16_xor0;
  wire f_s_dadda_rca16_u_rca30_fa16_and0;
  wire f_s_dadda_rca16_u_rca30_fa16_xor1;
  wire f_s_dadda_rca16_u_rca30_fa16_and1;
  wire f_s_dadda_rca16_u_rca30_fa16_or0;
  wire f_s_dadda_rca16_u_rca30_fa17_xor0;
  wire f_s_dadda_rca16_u_rca30_fa17_and0;
  wire f_s_dadda_rca16_u_rca30_fa17_xor1;
  wire f_s_dadda_rca16_u_rca30_fa17_and1;
  wire f_s_dadda_rca16_u_rca30_fa17_or0;
  wire f_s_dadda_rca16_u_rca30_fa18_xor0;
  wire f_s_dadda_rca16_u_rca30_fa18_and0;
  wire f_s_dadda_rca16_u_rca30_fa18_xor1;
  wire f_s_dadda_rca16_u_rca30_fa18_and1;
  wire f_s_dadda_rca16_u_rca30_fa18_or0;
  wire f_s_dadda_rca16_u_rca30_fa19_xor0;
  wire f_s_dadda_rca16_u_rca30_fa19_and0;
  wire f_s_dadda_rca16_u_rca30_fa19_xor1;
  wire f_s_dadda_rca16_u_rca30_fa19_and1;
  wire f_s_dadda_rca16_u_rca30_fa19_or0;
  wire f_s_dadda_rca16_u_rca30_fa20_xor0;
  wire f_s_dadda_rca16_u_rca30_fa20_and0;
  wire f_s_dadda_rca16_u_rca30_fa20_xor1;
  wire f_s_dadda_rca16_u_rca30_fa20_and1;
  wire f_s_dadda_rca16_u_rca30_fa20_or0;
  wire f_s_dadda_rca16_u_rca30_fa21_xor0;
  wire f_s_dadda_rca16_u_rca30_fa21_and0;
  wire f_s_dadda_rca16_u_rca30_fa21_xor1;
  wire f_s_dadda_rca16_u_rca30_fa21_and1;
  wire f_s_dadda_rca16_u_rca30_fa21_or0;
  wire f_s_dadda_rca16_u_rca30_fa22_xor0;
  wire f_s_dadda_rca16_u_rca30_fa22_and0;
  wire f_s_dadda_rca16_u_rca30_fa22_xor1;
  wire f_s_dadda_rca16_u_rca30_fa22_and1;
  wire f_s_dadda_rca16_u_rca30_fa22_or0;
  wire f_s_dadda_rca16_u_rca30_fa23_xor0;
  wire f_s_dadda_rca16_u_rca30_fa23_and0;
  wire f_s_dadda_rca16_u_rca30_fa23_xor1;
  wire f_s_dadda_rca16_u_rca30_fa23_and1;
  wire f_s_dadda_rca16_u_rca30_fa23_or0;
  wire f_s_dadda_rca16_u_rca30_fa24_xor0;
  wire f_s_dadda_rca16_u_rca30_fa24_and0;
  wire f_s_dadda_rca16_u_rca30_fa24_xor1;
  wire f_s_dadda_rca16_u_rca30_fa24_and1;
  wire f_s_dadda_rca16_u_rca30_fa24_or0;
  wire f_s_dadda_rca16_u_rca30_fa25_xor0;
  wire f_s_dadda_rca16_u_rca30_fa25_and0;
  wire f_s_dadda_rca16_u_rca30_fa25_xor1;
  wire f_s_dadda_rca16_u_rca30_fa25_and1;
  wire f_s_dadda_rca16_u_rca30_fa25_or0;
  wire f_s_dadda_rca16_u_rca30_fa26_xor0;
  wire f_s_dadda_rca16_u_rca30_fa26_and0;
  wire f_s_dadda_rca16_u_rca30_fa26_xor1;
  wire f_s_dadda_rca16_u_rca30_fa26_and1;
  wire f_s_dadda_rca16_u_rca30_fa26_or0;
  wire f_s_dadda_rca16_u_rca30_fa27_xor0;
  wire f_s_dadda_rca16_u_rca30_fa27_and0;
  wire f_s_dadda_rca16_u_rca30_fa27_xor1;
  wire f_s_dadda_rca16_u_rca30_fa27_and1;
  wire f_s_dadda_rca16_u_rca30_fa27_or0;
  wire f_s_dadda_rca16_u_rca30_fa28_xor0;
  wire f_s_dadda_rca16_u_rca30_fa28_and0;
  wire f_s_dadda_rca16_u_rca30_fa28_xor1;
  wire f_s_dadda_rca16_u_rca30_fa28_and1;
  wire f_s_dadda_rca16_u_rca30_fa28_or0;
  wire f_s_dadda_rca16_u_rca30_fa29_xor0;
  wire f_s_dadda_rca16_u_rca30_fa29_and0;
  wire f_s_dadda_rca16_u_rca30_fa29_xor1;
  wire f_s_dadda_rca16_u_rca30_fa29_and1;
  wire f_s_dadda_rca16_u_rca30_fa29_or0;
  wire f_s_dadda_rca16_xor0;

  assign f_s_dadda_rca16_and_13_0 = a[13] & b[0];
  assign f_s_dadda_rca16_and_12_1 = a[12] & b[1];
  assign f_s_dadda_rca16_ha0_xor0 = f_s_dadda_rca16_and_13_0 ^ f_s_dadda_rca16_and_12_1;
  assign f_s_dadda_rca16_ha0_and0 = f_s_dadda_rca16_and_13_0 & f_s_dadda_rca16_and_12_1;
  assign f_s_dadda_rca16_and_14_0 = a[14] & b[0];
  assign f_s_dadda_rca16_and_13_1 = a[13] & b[1];
  assign f_s_dadda_rca16_fa0_xor0 = f_s_dadda_rca16_ha0_and0 ^ f_s_dadda_rca16_and_14_0;
  assign f_s_dadda_rca16_fa0_and0 = f_s_dadda_rca16_ha0_and0 & f_s_dadda_rca16_and_14_0;
  assign f_s_dadda_rca16_fa0_xor1 = f_s_dadda_rca16_fa0_xor0 ^ f_s_dadda_rca16_and_13_1;
  assign f_s_dadda_rca16_fa0_and1 = f_s_dadda_rca16_fa0_xor0 & f_s_dadda_rca16_and_13_1;
  assign f_s_dadda_rca16_fa0_or0 = f_s_dadda_rca16_fa0_and0 | f_s_dadda_rca16_fa0_and1;
  assign f_s_dadda_rca16_and_12_2 = a[12] & b[2];
  assign f_s_dadda_rca16_and_11_3 = a[11] & b[3];
  assign f_s_dadda_rca16_ha1_xor0 = f_s_dadda_rca16_and_12_2 ^ f_s_dadda_rca16_and_11_3;
  assign f_s_dadda_rca16_ha1_and0 = f_s_dadda_rca16_and_12_2 & f_s_dadda_rca16_and_11_3;
  assign f_s_dadda_rca16_nand_15_0 = ~(a[15] & b[0]);
  assign f_s_dadda_rca16_fa1_xor0 = f_s_dadda_rca16_ha1_and0 ^ f_s_dadda_rca16_fa0_or0;
  assign f_s_dadda_rca16_fa1_and0 = f_s_dadda_rca16_ha1_and0 & f_s_dadda_rca16_fa0_or0;
  assign f_s_dadda_rca16_fa1_xor1 = f_s_dadda_rca16_fa1_xor0 ^ f_s_dadda_rca16_nand_15_0;
  assign f_s_dadda_rca16_fa1_and1 = f_s_dadda_rca16_fa1_xor0 & f_s_dadda_rca16_nand_15_0;
  assign f_s_dadda_rca16_fa1_or0 = f_s_dadda_rca16_fa1_and0 | f_s_dadda_rca16_fa1_and1;
  assign f_s_dadda_rca16_and_14_1 = a[14] & b[1];
  assign f_s_dadda_rca16_and_13_2 = a[13] & b[2];
  assign f_s_dadda_rca16_and_12_3 = a[12] & b[3];
  assign f_s_dadda_rca16_fa2_xor0 = f_s_dadda_rca16_and_14_1 ^ f_s_dadda_rca16_and_13_2;
  assign f_s_dadda_rca16_fa2_and0 = f_s_dadda_rca16_and_14_1 & f_s_dadda_rca16_and_13_2;
  assign f_s_dadda_rca16_fa2_xor1 = f_s_dadda_rca16_fa2_xor0 ^ f_s_dadda_rca16_and_12_3;
  assign f_s_dadda_rca16_fa2_and1 = f_s_dadda_rca16_fa2_xor0 & f_s_dadda_rca16_and_12_3;
  assign f_s_dadda_rca16_fa2_or0 = f_s_dadda_rca16_fa2_and0 | f_s_dadda_rca16_fa2_and1;
  assign f_s_dadda_rca16_and_11_4 = a[11] & b[4];
  assign f_s_dadda_rca16_and_10_5 = a[10] & b[5];
  assign f_s_dadda_rca16_ha2_xor0 = f_s_dadda_rca16_and_11_4 ^ f_s_dadda_rca16_and_10_5;
  assign f_s_dadda_rca16_ha2_and0 = f_s_dadda_rca16_and_11_4 & f_s_dadda_rca16_and_10_5;
  assign f_s_dadda_rca16_fa3_xor0 = f_s_dadda_rca16_ha2_and0 ^ f_s_dadda_rca16_fa2_or0;
  assign f_s_dadda_rca16_fa3_and0 = f_s_dadda_rca16_ha2_and0 & f_s_dadda_rca16_fa2_or0;
  assign f_s_dadda_rca16_fa3_xor1 = f_s_dadda_rca16_fa3_xor0 ^ f_s_dadda_rca16_fa1_or0;
  assign f_s_dadda_rca16_fa3_and1 = f_s_dadda_rca16_fa3_xor0 & f_s_dadda_rca16_fa1_or0;
  assign f_s_dadda_rca16_fa3_or0 = f_s_dadda_rca16_fa3_and0 | f_s_dadda_rca16_fa3_and1;
  assign f_s_dadda_rca16_nand_15_1 = ~(a[15] & b[1]);
  assign f_s_dadda_rca16_and_14_2 = a[14] & b[2];
  assign f_s_dadda_rca16_fa4_xor0 = ~f_s_dadda_rca16_nand_15_1;
  assign f_s_dadda_rca16_fa4_xor1 = f_s_dadda_rca16_fa4_xor0 ^ f_s_dadda_rca16_and_14_2;
  assign f_s_dadda_rca16_fa4_and1 = f_s_dadda_rca16_fa4_xor0 & f_s_dadda_rca16_and_14_2;
  assign f_s_dadda_rca16_fa4_or0 = f_s_dadda_rca16_nand_15_1 | f_s_dadda_rca16_fa4_and1;
  assign f_s_dadda_rca16_and_13_3 = a[13] & b[3];
  assign f_s_dadda_rca16_and_12_4 = a[12] & b[4];
  assign f_s_dadda_rca16_and_11_5 = a[11] & b[5];
  assign f_s_dadda_rca16_fa5_xor0 = f_s_dadda_rca16_and_13_3 ^ f_s_dadda_rca16_and_12_4;
  assign f_s_dadda_rca16_fa5_and0 = f_s_dadda_rca16_and_13_3 & f_s_dadda_rca16_and_12_4;
  assign f_s_dadda_rca16_fa5_xor1 = f_s_dadda_rca16_fa5_xor0 ^ f_s_dadda_rca16_and_11_5;
  assign f_s_dadda_rca16_fa5_and1 = f_s_dadda_rca16_fa5_xor0 & f_s_dadda_rca16_and_11_5;
  assign f_s_dadda_rca16_fa5_or0 = f_s_dadda_rca16_fa5_and0 | f_s_dadda_rca16_fa5_and1;
  assign f_s_dadda_rca16_fa6_xor0 = f_s_dadda_rca16_fa5_or0 ^ f_s_dadda_rca16_fa4_or0;
  assign f_s_dadda_rca16_fa6_and0 = f_s_dadda_rca16_fa5_or0 & f_s_dadda_rca16_fa4_or0;
  assign f_s_dadda_rca16_fa6_xor1 = f_s_dadda_rca16_fa6_xor0 ^ f_s_dadda_rca16_fa3_or0;
  assign f_s_dadda_rca16_fa6_and1 = f_s_dadda_rca16_fa6_xor0 & f_s_dadda_rca16_fa3_or0;
  assign f_s_dadda_rca16_fa6_or0 = f_s_dadda_rca16_fa6_and0 | f_s_dadda_rca16_fa6_and1;
  assign f_s_dadda_rca16_nand_15_2 = ~(a[15] & b[2]);
  assign f_s_dadda_rca16_and_14_3 = a[14] & b[3];
  assign f_s_dadda_rca16_and_13_4 = a[13] & b[4];
  assign f_s_dadda_rca16_fa7_xor0 = f_s_dadda_rca16_nand_15_2 ^ f_s_dadda_rca16_and_14_3;
  assign f_s_dadda_rca16_fa7_and0 = f_s_dadda_rca16_nand_15_2 & f_s_dadda_rca16_and_14_3;
  assign f_s_dadda_rca16_fa7_xor1 = f_s_dadda_rca16_fa7_xor0 ^ f_s_dadda_rca16_and_13_4;
  assign f_s_dadda_rca16_fa7_and1 = f_s_dadda_rca16_fa7_xor0 & f_s_dadda_rca16_and_13_4;
  assign f_s_dadda_rca16_fa7_or0 = f_s_dadda_rca16_fa7_and0 | f_s_dadda_rca16_fa7_and1;
  assign f_s_dadda_rca16_nand_15_3 = ~(a[15] & b[3]);
  assign f_s_dadda_rca16_fa8_xor0 = f_s_dadda_rca16_fa7_or0 ^ f_s_dadda_rca16_fa6_or0;
  assign f_s_dadda_rca16_fa8_and0 = f_s_dadda_rca16_fa7_or0 & f_s_dadda_rca16_fa6_or0;
  assign f_s_dadda_rca16_fa8_xor1 = f_s_dadda_rca16_fa8_xor0 ^ f_s_dadda_rca16_nand_15_3;
  assign f_s_dadda_rca16_fa8_and1 = f_s_dadda_rca16_fa8_xor0 & f_s_dadda_rca16_nand_15_3;
  assign f_s_dadda_rca16_fa8_or0 = f_s_dadda_rca16_fa8_and0 | f_s_dadda_rca16_fa8_and1;
  assign f_s_dadda_rca16_and_4_0 = a[4] & b[0];
  assign f_s_dadda_rca16_and_3_1 = a[3] & b[1];
  assign f_s_dadda_rca16_ha3_xor0 = f_s_dadda_rca16_and_4_0 ^ f_s_dadda_rca16_and_3_1;
  assign f_s_dadda_rca16_ha3_and0 = f_s_dadda_rca16_and_4_0 & f_s_dadda_rca16_and_3_1;
  assign f_s_dadda_rca16_and_5_0 = a[5] & b[0];
  assign f_s_dadda_rca16_and_4_1 = a[4] & b[1];
  assign f_s_dadda_rca16_fa9_xor0 = f_s_dadda_rca16_ha3_and0 ^ f_s_dadda_rca16_and_5_0;
  assign f_s_dadda_rca16_fa9_and0 = f_s_dadda_rca16_ha3_and0 & f_s_dadda_rca16_and_5_0;
  assign f_s_dadda_rca16_fa9_xor1 = f_s_dadda_rca16_fa9_xor0 ^ f_s_dadda_rca16_and_4_1;
  assign f_s_dadda_rca16_fa9_and1 = f_s_dadda_rca16_fa9_xor0 & f_s_dadda_rca16_and_4_1;
  assign f_s_dadda_rca16_fa9_or0 = f_s_dadda_rca16_fa9_and0 | f_s_dadda_rca16_fa9_and1;
  assign f_s_dadda_rca16_and_3_2 = a[3] & b[2];
  assign f_s_dadda_rca16_and_2_3 = a[2] & b[3];
  assign f_s_dadda_rca16_ha4_xor0 = f_s_dadda_rca16_and_3_2 ^ f_s_dadda_rca16_and_2_3;
  assign f_s_dadda_rca16_ha4_and0 = f_s_dadda_rca16_and_3_2 & f_s_dadda_rca16_and_2_3;
  assign f_s_dadda_rca16_and_6_0 = a[6] & b[0];
  assign f_s_dadda_rca16_fa10_xor0 = f_s_dadda_rca16_ha4_and0 ^ f_s_dadda_rca16_fa9_or0;
  assign f_s_dadda_rca16_fa10_and0 = f_s_dadda_rca16_ha4_and0 & f_s_dadda_rca16_fa9_or0;
  assign f_s_dadda_rca16_fa10_xor1 = f_s_dadda_rca16_fa10_xor0 ^ f_s_dadda_rca16_and_6_0;
  assign f_s_dadda_rca16_fa10_and1 = f_s_dadda_rca16_fa10_xor0 & f_s_dadda_rca16_and_6_0;
  assign f_s_dadda_rca16_fa10_or0 = f_s_dadda_rca16_fa10_and0 | f_s_dadda_rca16_fa10_and1;
  assign f_s_dadda_rca16_and_5_1 = a[5] & b[1];
  assign f_s_dadda_rca16_and_4_2 = a[4] & b[2];
  assign f_s_dadda_rca16_and_3_3 = a[3] & b[3];
  assign f_s_dadda_rca16_fa11_xor0 = f_s_dadda_rca16_and_5_1 ^ f_s_dadda_rca16_and_4_2;
  assign f_s_dadda_rca16_fa11_and0 = f_s_dadda_rca16_and_5_1 & f_s_dadda_rca16_and_4_2;
  assign f_s_dadda_rca16_fa11_xor1 = f_s_dadda_rca16_fa11_xor0 ^ f_s_dadda_rca16_and_3_3;
  assign f_s_dadda_rca16_fa11_and1 = f_s_dadda_rca16_fa11_xor0 & f_s_dadda_rca16_and_3_3;
  assign f_s_dadda_rca16_fa11_or0 = f_s_dadda_rca16_fa11_and0 | f_s_dadda_rca16_fa11_and1;
  assign f_s_dadda_rca16_and_2_4 = a[2] & b[4];
  assign f_s_dadda_rca16_and_1_5 = a[1] & b[5];
  assign f_s_dadda_rca16_ha5_xor0 = f_s_dadda_rca16_and_2_4 ^ f_s_dadda_rca16_and_1_5;
  assign f_s_dadda_rca16_ha5_and0 = f_s_dadda_rca16_and_2_4 & f_s_dadda_rca16_and_1_5;
  assign f_s_dadda_rca16_fa12_xor0 = f_s_dadda_rca16_ha5_and0 ^ f_s_dadda_rca16_fa11_or0;
  assign f_s_dadda_rca16_fa12_and0 = f_s_dadda_rca16_ha5_and0 & f_s_dadda_rca16_fa11_or0;
  assign f_s_dadda_rca16_fa12_xor1 = f_s_dadda_rca16_fa12_xor0 ^ f_s_dadda_rca16_fa10_or0;
  assign f_s_dadda_rca16_fa12_and1 = f_s_dadda_rca16_fa12_xor0 & f_s_dadda_rca16_fa10_or0;
  assign f_s_dadda_rca16_fa12_or0 = f_s_dadda_rca16_fa12_and0 | f_s_dadda_rca16_fa12_and1;
  assign f_s_dadda_rca16_and_7_0 = a[7] & b[0];
  assign f_s_dadda_rca16_and_6_1 = a[6] & b[1];
  assign f_s_dadda_rca16_and_5_2 = a[5] & b[2];
  assign f_s_dadda_rca16_fa13_xor0 = f_s_dadda_rca16_and_7_0 ^ f_s_dadda_rca16_and_6_1;
  assign f_s_dadda_rca16_fa13_and0 = f_s_dadda_rca16_and_7_0 & f_s_dadda_rca16_and_6_1;
  assign f_s_dadda_rca16_fa13_xor1 = f_s_dadda_rca16_fa13_xor0 ^ f_s_dadda_rca16_and_5_2;
  assign f_s_dadda_rca16_fa13_and1 = f_s_dadda_rca16_fa13_xor0 & f_s_dadda_rca16_and_5_2;
  assign f_s_dadda_rca16_fa13_or0 = f_s_dadda_rca16_fa13_and0 | f_s_dadda_rca16_fa13_and1;
  assign f_s_dadda_rca16_and_4_3 = a[4] & b[3];
  assign f_s_dadda_rca16_and_3_4 = a[3] & b[4];
  assign f_s_dadda_rca16_and_2_5 = a[2] & b[5];
  assign f_s_dadda_rca16_fa14_xor0 = f_s_dadda_rca16_and_4_3 ^ f_s_dadda_rca16_and_3_4;
  assign f_s_dadda_rca16_fa14_and0 = f_s_dadda_rca16_and_4_3 & f_s_dadda_rca16_and_3_4;
  assign f_s_dadda_rca16_fa14_xor1 = f_s_dadda_rca16_fa14_xor0 ^ f_s_dadda_rca16_and_2_5;
  assign f_s_dadda_rca16_fa14_and1 = f_s_dadda_rca16_fa14_xor0 & f_s_dadda_rca16_and_2_5;
  assign f_s_dadda_rca16_fa14_or0 = f_s_dadda_rca16_fa14_and0 | f_s_dadda_rca16_fa14_and1;
  assign f_s_dadda_rca16_and_1_6 = a[1] & b[6];
  assign f_s_dadda_rca16_and_0_7 = a[0] & b[7];
  assign f_s_dadda_rca16_ha6_xor0 = f_s_dadda_rca16_and_1_6 ^ f_s_dadda_rca16_and_0_7;
  assign f_s_dadda_rca16_ha6_and0 = f_s_dadda_rca16_and_1_6 & f_s_dadda_rca16_and_0_7;
  assign f_s_dadda_rca16_fa15_xor0 = f_s_dadda_rca16_ha6_and0 ^ f_s_dadda_rca16_fa14_or0;
  assign f_s_dadda_rca16_fa15_and0 = f_s_dadda_rca16_ha6_and0 & f_s_dadda_rca16_fa14_or0;
  assign f_s_dadda_rca16_fa15_xor1 = f_s_dadda_rca16_fa15_xor0 ^ f_s_dadda_rca16_fa13_or0;
  assign f_s_dadda_rca16_fa15_and1 = f_s_dadda_rca16_fa15_xor0 & f_s_dadda_rca16_fa13_or0;
  assign f_s_dadda_rca16_fa15_or0 = f_s_dadda_rca16_fa15_and0 | f_s_dadda_rca16_fa15_and1;
  assign f_s_dadda_rca16_and_8_0 = a[8] & b[0];
  assign f_s_dadda_rca16_and_7_1 = a[7] & b[1];
  assign f_s_dadda_rca16_fa16_xor0 = f_s_dadda_rca16_fa12_or0 ^ f_s_dadda_rca16_and_8_0;
  assign f_s_dadda_rca16_fa16_and0 = f_s_dadda_rca16_fa12_or0 & f_s_dadda_rca16_and_8_0;
  assign f_s_dadda_rca16_fa16_xor1 = f_s_dadda_rca16_fa16_xor0 ^ f_s_dadda_rca16_and_7_1;
  assign f_s_dadda_rca16_fa16_and1 = f_s_dadda_rca16_fa16_xor0 & f_s_dadda_rca16_and_7_1;
  assign f_s_dadda_rca16_fa16_or0 = f_s_dadda_rca16_fa16_and0 | f_s_dadda_rca16_fa16_and1;
  assign f_s_dadda_rca16_and_6_2 = a[6] & b[2];
  assign f_s_dadda_rca16_and_5_3 = a[5] & b[3];
  assign f_s_dadda_rca16_and_4_4 = a[4] & b[4];
  assign f_s_dadda_rca16_fa17_xor0 = f_s_dadda_rca16_and_6_2 ^ f_s_dadda_rca16_and_5_3;
  assign f_s_dadda_rca16_fa17_and0 = f_s_dadda_rca16_and_6_2 & f_s_dadda_rca16_and_5_3;
  assign f_s_dadda_rca16_fa17_xor1 = f_s_dadda_rca16_fa17_xor0 ^ f_s_dadda_rca16_and_4_4;
  assign f_s_dadda_rca16_fa17_and1 = f_s_dadda_rca16_fa17_xor0 & f_s_dadda_rca16_and_4_4;
  assign f_s_dadda_rca16_fa17_or0 = f_s_dadda_rca16_fa17_and0 | f_s_dadda_rca16_fa17_and1;
  assign f_s_dadda_rca16_and_3_5 = a[3] & b[5];
  assign f_s_dadda_rca16_and_2_6 = a[2] & b[6];
  assign f_s_dadda_rca16_and_1_7 = a[1] & b[7];
  assign f_s_dadda_rca16_fa18_xor0 = f_s_dadda_rca16_and_3_5 ^ f_s_dadda_rca16_and_2_6;
  assign f_s_dadda_rca16_fa18_and0 = f_s_dadda_rca16_and_3_5 & f_s_dadda_rca16_and_2_6;
  assign f_s_dadda_rca16_fa18_xor1 = f_s_dadda_rca16_fa18_xor0 ^ f_s_dadda_rca16_and_1_7;
  assign f_s_dadda_rca16_fa18_and1 = f_s_dadda_rca16_fa18_xor0 & f_s_dadda_rca16_and_1_7;
  assign f_s_dadda_rca16_fa18_or0 = f_s_dadda_rca16_fa18_and0 | f_s_dadda_rca16_fa18_and1;
  assign f_s_dadda_rca16_and_0_8 = a[0] & b[8];
  assign f_s_dadda_rca16_ha7_xor0 = f_s_dadda_rca16_and_0_8 ^ f_s_dadda_rca16_fa15_xor1;
  assign f_s_dadda_rca16_ha7_and0 = f_s_dadda_rca16_and_0_8 & f_s_dadda_rca16_fa15_xor1;
  assign f_s_dadda_rca16_fa19_xor0 = f_s_dadda_rca16_ha7_and0 ^ f_s_dadda_rca16_fa18_or0;
  assign f_s_dadda_rca16_fa19_and0 = f_s_dadda_rca16_ha7_and0 & f_s_dadda_rca16_fa18_or0;
  assign f_s_dadda_rca16_fa19_xor1 = f_s_dadda_rca16_fa19_xor0 ^ f_s_dadda_rca16_fa17_or0;
  assign f_s_dadda_rca16_fa19_and1 = f_s_dadda_rca16_fa19_xor0 & f_s_dadda_rca16_fa17_or0;
  assign f_s_dadda_rca16_fa19_or0 = f_s_dadda_rca16_fa19_and0 | f_s_dadda_rca16_fa19_and1;
  assign f_s_dadda_rca16_and_9_0 = a[9] & b[0];
  assign f_s_dadda_rca16_fa20_xor0 = f_s_dadda_rca16_fa16_or0 ^ f_s_dadda_rca16_fa15_or0;
  assign f_s_dadda_rca16_fa20_and0 = f_s_dadda_rca16_fa16_or0 & f_s_dadda_rca16_fa15_or0;
  assign f_s_dadda_rca16_fa20_xor1 = f_s_dadda_rca16_fa20_xor0 ^ f_s_dadda_rca16_and_9_0;
  assign f_s_dadda_rca16_fa20_and1 = f_s_dadda_rca16_fa20_xor0 & f_s_dadda_rca16_and_9_0;
  assign f_s_dadda_rca16_fa20_or0 = f_s_dadda_rca16_fa20_and0 | f_s_dadda_rca16_fa20_and1;
  assign f_s_dadda_rca16_and_8_1 = a[8] & b[1];
  assign f_s_dadda_rca16_and_7_2 = a[7] & b[2];
  assign f_s_dadda_rca16_and_6_3 = a[6] & b[3];
  assign f_s_dadda_rca16_fa21_xor0 = f_s_dadda_rca16_and_8_1 ^ f_s_dadda_rca16_and_7_2;
  assign f_s_dadda_rca16_fa21_and0 = f_s_dadda_rca16_and_8_1 & f_s_dadda_rca16_and_7_2;
  assign f_s_dadda_rca16_fa21_xor1 = f_s_dadda_rca16_fa21_xor0 ^ f_s_dadda_rca16_and_6_3;
  assign f_s_dadda_rca16_fa21_and1 = f_s_dadda_rca16_fa21_xor0 & f_s_dadda_rca16_and_6_3;
  assign f_s_dadda_rca16_fa21_or0 = f_s_dadda_rca16_fa21_and0 | f_s_dadda_rca16_fa21_and1;
  assign f_s_dadda_rca16_and_5_4 = a[5] & b[4];
  assign f_s_dadda_rca16_and_4_5 = a[4] & b[5];
  assign f_s_dadda_rca16_and_3_6 = a[3] & b[6];
  assign f_s_dadda_rca16_fa22_xor0 = f_s_dadda_rca16_and_5_4 ^ f_s_dadda_rca16_and_4_5;
  assign f_s_dadda_rca16_fa22_and0 = f_s_dadda_rca16_and_5_4 & f_s_dadda_rca16_and_4_5;
  assign f_s_dadda_rca16_fa22_xor1 = f_s_dadda_rca16_fa22_xor0 ^ f_s_dadda_rca16_and_3_6;
  assign f_s_dadda_rca16_fa22_and1 = f_s_dadda_rca16_fa22_xor0 & f_s_dadda_rca16_and_3_6;
  assign f_s_dadda_rca16_fa22_or0 = f_s_dadda_rca16_fa22_and0 | f_s_dadda_rca16_fa22_and1;
  assign f_s_dadda_rca16_and_2_7 = a[2] & b[7];
  assign f_s_dadda_rca16_and_1_8 = a[1] & b[8];
  assign f_s_dadda_rca16_and_0_9 = a[0] & b[9];
  assign f_s_dadda_rca16_fa23_xor0 = f_s_dadda_rca16_and_2_7 ^ f_s_dadda_rca16_and_1_8;
  assign f_s_dadda_rca16_fa23_and0 = f_s_dadda_rca16_and_2_7 & f_s_dadda_rca16_and_1_8;
  assign f_s_dadda_rca16_fa23_xor1 = f_s_dadda_rca16_fa23_xor0 ^ f_s_dadda_rca16_and_0_9;
  assign f_s_dadda_rca16_fa23_and1 = f_s_dadda_rca16_fa23_xor0 & f_s_dadda_rca16_and_0_9;
  assign f_s_dadda_rca16_fa23_or0 = f_s_dadda_rca16_fa23_and0 | f_s_dadda_rca16_fa23_and1;
  assign f_s_dadda_rca16_ha8_xor0 = f_s_dadda_rca16_fa19_xor1 ^ f_s_dadda_rca16_fa20_xor1;
  assign f_s_dadda_rca16_ha8_and0 = f_s_dadda_rca16_fa19_xor1 & f_s_dadda_rca16_fa20_xor1;
  assign f_s_dadda_rca16_fa24_xor0 = f_s_dadda_rca16_ha8_and0 ^ f_s_dadda_rca16_fa23_or0;
  assign f_s_dadda_rca16_fa24_and0 = f_s_dadda_rca16_ha8_and0 & f_s_dadda_rca16_fa23_or0;
  assign f_s_dadda_rca16_fa24_xor1 = f_s_dadda_rca16_fa24_xor0 ^ f_s_dadda_rca16_fa22_or0;
  assign f_s_dadda_rca16_fa24_and1 = f_s_dadda_rca16_fa24_xor0 & f_s_dadda_rca16_fa22_or0;
  assign f_s_dadda_rca16_fa24_or0 = f_s_dadda_rca16_fa24_and0 | f_s_dadda_rca16_fa24_and1;
  assign f_s_dadda_rca16_fa25_xor0 = f_s_dadda_rca16_fa21_or0 ^ f_s_dadda_rca16_fa20_or0;
  assign f_s_dadda_rca16_fa25_and0 = f_s_dadda_rca16_fa21_or0 & f_s_dadda_rca16_fa20_or0;
  assign f_s_dadda_rca16_fa25_xor1 = f_s_dadda_rca16_fa25_xor0 ^ f_s_dadda_rca16_fa19_or0;
  assign f_s_dadda_rca16_fa25_and1 = f_s_dadda_rca16_fa25_xor0 & f_s_dadda_rca16_fa19_or0;
  assign f_s_dadda_rca16_fa25_or0 = f_s_dadda_rca16_fa25_and0 | f_s_dadda_rca16_fa25_and1;
  assign f_s_dadda_rca16_and_10_0 = a[10] & b[0];
  assign f_s_dadda_rca16_and_9_1 = a[9] & b[1];
  assign f_s_dadda_rca16_and_8_2 = a[8] & b[2];
  assign f_s_dadda_rca16_fa26_xor0 = f_s_dadda_rca16_and_10_0 ^ f_s_dadda_rca16_and_9_1;
  assign f_s_dadda_rca16_fa26_and0 = f_s_dadda_rca16_and_10_0 & f_s_dadda_rca16_and_9_1;
  assign f_s_dadda_rca16_fa26_xor1 = f_s_dadda_rca16_fa26_xor0 ^ f_s_dadda_rca16_and_8_2;
  assign f_s_dadda_rca16_fa26_and1 = f_s_dadda_rca16_fa26_xor0 & f_s_dadda_rca16_and_8_2;
  assign f_s_dadda_rca16_fa26_or0 = f_s_dadda_rca16_fa26_and0 | f_s_dadda_rca16_fa26_and1;
  assign f_s_dadda_rca16_and_7_3 = a[7] & b[3];
  assign f_s_dadda_rca16_and_6_4 = a[6] & b[4];
  assign f_s_dadda_rca16_and_5_5 = a[5] & b[5];
  assign f_s_dadda_rca16_fa27_xor0 = f_s_dadda_rca16_and_7_3 ^ f_s_dadda_rca16_and_6_4;
  assign f_s_dadda_rca16_fa27_and0 = f_s_dadda_rca16_and_7_3 & f_s_dadda_rca16_and_6_4;
  assign f_s_dadda_rca16_fa27_xor1 = f_s_dadda_rca16_fa27_xor0 ^ f_s_dadda_rca16_and_5_5;
  assign f_s_dadda_rca16_fa27_and1 = f_s_dadda_rca16_fa27_xor0 & f_s_dadda_rca16_and_5_5;
  assign f_s_dadda_rca16_fa27_or0 = f_s_dadda_rca16_fa27_and0 | f_s_dadda_rca16_fa27_and1;
  assign f_s_dadda_rca16_and_4_6 = a[4] & b[6];
  assign f_s_dadda_rca16_and_3_7 = a[3] & b[7];
  assign f_s_dadda_rca16_and_2_8 = a[2] & b[8];
  assign f_s_dadda_rca16_fa28_xor0 = f_s_dadda_rca16_and_4_6 ^ f_s_dadda_rca16_and_3_7;
  assign f_s_dadda_rca16_fa28_and0 = f_s_dadda_rca16_and_4_6 & f_s_dadda_rca16_and_3_7;
  assign f_s_dadda_rca16_fa28_xor1 = f_s_dadda_rca16_fa28_xor0 ^ f_s_dadda_rca16_and_2_8;
  assign f_s_dadda_rca16_fa28_and1 = f_s_dadda_rca16_fa28_xor0 & f_s_dadda_rca16_and_2_8;
  assign f_s_dadda_rca16_fa28_or0 = f_s_dadda_rca16_fa28_and0 | f_s_dadda_rca16_fa28_and1;
  assign f_s_dadda_rca16_and_1_9 = a[1] & b[9];
  assign f_s_dadda_rca16_and_0_10 = a[0] & b[10];
  assign f_s_dadda_rca16_fa29_xor0 = f_s_dadda_rca16_and_1_9 ^ f_s_dadda_rca16_and_0_10;
  assign f_s_dadda_rca16_fa29_and0 = f_s_dadda_rca16_and_1_9 & f_s_dadda_rca16_and_0_10;
  assign f_s_dadda_rca16_fa29_xor1 = f_s_dadda_rca16_fa29_xor0 ^ f_s_dadda_rca16_fa24_xor1;
  assign f_s_dadda_rca16_fa29_and1 = f_s_dadda_rca16_fa29_xor0 & f_s_dadda_rca16_fa24_xor1;
  assign f_s_dadda_rca16_fa29_or0 = f_s_dadda_rca16_fa29_and0 | f_s_dadda_rca16_fa29_and1;
  assign f_s_dadda_rca16_ha9_xor0 = f_s_dadda_rca16_fa25_xor1 ^ f_s_dadda_rca16_fa26_xor1;
  assign f_s_dadda_rca16_ha9_and0 = f_s_dadda_rca16_fa25_xor1 & f_s_dadda_rca16_fa26_xor1;
  assign f_s_dadda_rca16_fa30_xor0 = f_s_dadda_rca16_ha9_and0 ^ f_s_dadda_rca16_fa29_or0;
  assign f_s_dadda_rca16_fa30_and0 = f_s_dadda_rca16_ha9_and0 & f_s_dadda_rca16_fa29_or0;
  assign f_s_dadda_rca16_fa30_xor1 = f_s_dadda_rca16_fa30_xor0 ^ f_s_dadda_rca16_fa28_or0;
  assign f_s_dadda_rca16_fa30_and1 = f_s_dadda_rca16_fa30_xor0 & f_s_dadda_rca16_fa28_or0;
  assign f_s_dadda_rca16_fa30_or0 = f_s_dadda_rca16_fa30_and0 | f_s_dadda_rca16_fa30_and1;
  assign f_s_dadda_rca16_fa31_xor0 = f_s_dadda_rca16_fa27_or0 ^ f_s_dadda_rca16_fa26_or0;
  assign f_s_dadda_rca16_fa31_and0 = f_s_dadda_rca16_fa27_or0 & f_s_dadda_rca16_fa26_or0;
  assign f_s_dadda_rca16_fa31_xor1 = f_s_dadda_rca16_fa31_xor0 ^ f_s_dadda_rca16_fa25_or0;
  assign f_s_dadda_rca16_fa31_and1 = f_s_dadda_rca16_fa31_xor0 & f_s_dadda_rca16_fa25_or0;
  assign f_s_dadda_rca16_fa31_or0 = f_s_dadda_rca16_fa31_and0 | f_s_dadda_rca16_fa31_and1;
  assign f_s_dadda_rca16_and_11_0 = a[11] & b[0];
  assign f_s_dadda_rca16_and_10_1 = a[10] & b[1];
  assign f_s_dadda_rca16_fa32_xor0 = f_s_dadda_rca16_fa24_or0 ^ f_s_dadda_rca16_and_11_0;
  assign f_s_dadda_rca16_fa32_and0 = f_s_dadda_rca16_fa24_or0 & f_s_dadda_rca16_and_11_0;
  assign f_s_dadda_rca16_fa32_xor1 = f_s_dadda_rca16_fa32_xor0 ^ f_s_dadda_rca16_and_10_1;
  assign f_s_dadda_rca16_fa32_and1 = f_s_dadda_rca16_fa32_xor0 & f_s_dadda_rca16_and_10_1;
  assign f_s_dadda_rca16_fa32_or0 = f_s_dadda_rca16_fa32_and0 | f_s_dadda_rca16_fa32_and1;
  assign f_s_dadda_rca16_and_9_2 = a[9] & b[2];
  assign f_s_dadda_rca16_and_8_3 = a[8] & b[3];
  assign f_s_dadda_rca16_and_7_4 = a[7] & b[4];
  assign f_s_dadda_rca16_fa33_xor0 = f_s_dadda_rca16_and_9_2 ^ f_s_dadda_rca16_and_8_3;
  assign f_s_dadda_rca16_fa33_and0 = f_s_dadda_rca16_and_9_2 & f_s_dadda_rca16_and_8_3;
  assign f_s_dadda_rca16_fa33_xor1 = f_s_dadda_rca16_fa33_xor0 ^ f_s_dadda_rca16_and_7_4;
  assign f_s_dadda_rca16_fa33_and1 = f_s_dadda_rca16_fa33_xor0 & f_s_dadda_rca16_and_7_4;
  assign f_s_dadda_rca16_fa33_or0 = f_s_dadda_rca16_fa33_and0 | f_s_dadda_rca16_fa33_and1;
  assign f_s_dadda_rca16_and_6_5 = a[6] & b[5];
  assign f_s_dadda_rca16_and_5_6 = a[5] & b[6];
  assign f_s_dadda_rca16_and_4_7 = a[4] & b[7];
  assign f_s_dadda_rca16_fa34_xor0 = f_s_dadda_rca16_and_6_5 ^ f_s_dadda_rca16_and_5_6;
  assign f_s_dadda_rca16_fa34_and0 = f_s_dadda_rca16_and_6_5 & f_s_dadda_rca16_and_5_6;
  assign f_s_dadda_rca16_fa34_xor1 = f_s_dadda_rca16_fa34_xor0 ^ f_s_dadda_rca16_and_4_7;
  assign f_s_dadda_rca16_fa34_and1 = f_s_dadda_rca16_fa34_xor0 & f_s_dadda_rca16_and_4_7;
  assign f_s_dadda_rca16_fa34_or0 = f_s_dadda_rca16_fa34_and0 | f_s_dadda_rca16_fa34_and1;
  assign f_s_dadda_rca16_and_3_8 = a[3] & b[8];
  assign f_s_dadda_rca16_and_2_9 = a[2] & b[9];
  assign f_s_dadda_rca16_and_1_10 = a[1] & b[10];
  assign f_s_dadda_rca16_fa35_xor0 = f_s_dadda_rca16_and_3_8 ^ f_s_dadda_rca16_and_2_9;
  assign f_s_dadda_rca16_fa35_and0 = f_s_dadda_rca16_and_3_8 & f_s_dadda_rca16_and_2_9;
  assign f_s_dadda_rca16_fa35_xor1 = f_s_dadda_rca16_fa35_xor0 ^ f_s_dadda_rca16_and_1_10;
  assign f_s_dadda_rca16_fa35_and1 = f_s_dadda_rca16_fa35_xor0 & f_s_dadda_rca16_and_1_10;
  assign f_s_dadda_rca16_fa35_or0 = f_s_dadda_rca16_fa35_and0 | f_s_dadda_rca16_fa35_and1;
  assign f_s_dadda_rca16_and_0_11 = a[0] & b[11];
  assign f_s_dadda_rca16_fa36_xor0 = f_s_dadda_rca16_and_0_11 ^ f_s_dadda_rca16_fa30_xor1;
  assign f_s_dadda_rca16_fa36_and0 = f_s_dadda_rca16_and_0_11 & f_s_dadda_rca16_fa30_xor1;
  assign f_s_dadda_rca16_fa36_xor1 = f_s_dadda_rca16_fa36_xor0 ^ f_s_dadda_rca16_fa31_xor1;
  assign f_s_dadda_rca16_fa36_and1 = f_s_dadda_rca16_fa36_xor0 & f_s_dadda_rca16_fa31_xor1;
  assign f_s_dadda_rca16_fa36_or0 = f_s_dadda_rca16_fa36_and0 | f_s_dadda_rca16_fa36_and1;
  assign f_s_dadda_rca16_ha10_xor0 = f_s_dadda_rca16_fa32_xor1 ^ f_s_dadda_rca16_fa33_xor1;
  assign f_s_dadda_rca16_ha10_and0 = f_s_dadda_rca16_fa32_xor1 & f_s_dadda_rca16_fa33_xor1;
  assign f_s_dadda_rca16_fa37_xor0 = f_s_dadda_rca16_ha10_and0 ^ f_s_dadda_rca16_fa36_or0;
  assign f_s_dadda_rca16_fa37_and0 = f_s_dadda_rca16_ha10_and0 & f_s_dadda_rca16_fa36_or0;
  assign f_s_dadda_rca16_fa37_xor1 = f_s_dadda_rca16_fa37_xor0 ^ f_s_dadda_rca16_fa35_or0;
  assign f_s_dadda_rca16_fa37_and1 = f_s_dadda_rca16_fa37_xor0 & f_s_dadda_rca16_fa35_or0;
  assign f_s_dadda_rca16_fa37_or0 = f_s_dadda_rca16_fa37_and0 | f_s_dadda_rca16_fa37_and1;
  assign f_s_dadda_rca16_fa38_xor0 = f_s_dadda_rca16_fa34_or0 ^ f_s_dadda_rca16_fa33_or0;
  assign f_s_dadda_rca16_fa38_and0 = f_s_dadda_rca16_fa34_or0 & f_s_dadda_rca16_fa33_or0;
  assign f_s_dadda_rca16_fa38_xor1 = f_s_dadda_rca16_fa38_xor0 ^ f_s_dadda_rca16_fa32_or0;
  assign f_s_dadda_rca16_fa38_and1 = f_s_dadda_rca16_fa38_xor0 & f_s_dadda_rca16_fa32_or0;
  assign f_s_dadda_rca16_fa38_or0 = f_s_dadda_rca16_fa38_and0 | f_s_dadda_rca16_fa38_and1;
  assign f_s_dadda_rca16_and_12_0 = a[12] & b[0];
  assign f_s_dadda_rca16_fa39_xor0 = f_s_dadda_rca16_fa31_or0 ^ f_s_dadda_rca16_fa30_or0;
  assign f_s_dadda_rca16_fa39_and0 = f_s_dadda_rca16_fa31_or0 & f_s_dadda_rca16_fa30_or0;
  assign f_s_dadda_rca16_fa39_xor1 = f_s_dadda_rca16_fa39_xor0 ^ f_s_dadda_rca16_and_12_0;
  assign f_s_dadda_rca16_fa39_and1 = f_s_dadda_rca16_fa39_xor0 & f_s_dadda_rca16_and_12_0;
  assign f_s_dadda_rca16_fa39_or0 = f_s_dadda_rca16_fa39_and0 | f_s_dadda_rca16_fa39_and1;
  assign f_s_dadda_rca16_and_11_1 = a[11] & b[1];
  assign f_s_dadda_rca16_and_10_2 = a[10] & b[2];
  assign f_s_dadda_rca16_and_9_3 = a[9] & b[3];
  assign f_s_dadda_rca16_fa40_xor0 = f_s_dadda_rca16_and_11_1 ^ f_s_dadda_rca16_and_10_2;
  assign f_s_dadda_rca16_fa40_and0 = f_s_dadda_rca16_and_11_1 & f_s_dadda_rca16_and_10_2;
  assign f_s_dadda_rca16_fa40_xor1 = f_s_dadda_rca16_fa40_xor0 ^ f_s_dadda_rca16_and_9_3;
  assign f_s_dadda_rca16_fa40_and1 = f_s_dadda_rca16_fa40_xor0 & f_s_dadda_rca16_and_9_3;
  assign f_s_dadda_rca16_fa40_or0 = f_s_dadda_rca16_fa40_and0 | f_s_dadda_rca16_fa40_and1;
  assign f_s_dadda_rca16_and_8_4 = a[8] & b[4];
  assign f_s_dadda_rca16_and_7_5 = a[7] & b[5];
  assign f_s_dadda_rca16_and_6_6 = a[6] & b[6];
  assign f_s_dadda_rca16_fa41_xor0 = f_s_dadda_rca16_and_8_4 ^ f_s_dadda_rca16_and_7_5;
  assign f_s_dadda_rca16_fa41_and0 = f_s_dadda_rca16_and_8_4 & f_s_dadda_rca16_and_7_5;
  assign f_s_dadda_rca16_fa41_xor1 = f_s_dadda_rca16_fa41_xor0 ^ f_s_dadda_rca16_and_6_6;
  assign f_s_dadda_rca16_fa41_and1 = f_s_dadda_rca16_fa41_xor0 & f_s_dadda_rca16_and_6_6;
  assign f_s_dadda_rca16_fa41_or0 = f_s_dadda_rca16_fa41_and0 | f_s_dadda_rca16_fa41_and1;
  assign f_s_dadda_rca16_and_5_7 = a[5] & b[7];
  assign f_s_dadda_rca16_and_4_8 = a[4] & b[8];
  assign f_s_dadda_rca16_and_3_9 = a[3] & b[9];
  assign f_s_dadda_rca16_fa42_xor0 = f_s_dadda_rca16_and_5_7 ^ f_s_dadda_rca16_and_4_8;
  assign f_s_dadda_rca16_fa42_and0 = f_s_dadda_rca16_and_5_7 & f_s_dadda_rca16_and_4_8;
  assign f_s_dadda_rca16_fa42_xor1 = f_s_dadda_rca16_fa42_xor0 ^ f_s_dadda_rca16_and_3_9;
  assign f_s_dadda_rca16_fa42_and1 = f_s_dadda_rca16_fa42_xor0 & f_s_dadda_rca16_and_3_9;
  assign f_s_dadda_rca16_fa42_or0 = f_s_dadda_rca16_fa42_and0 | f_s_dadda_rca16_fa42_and1;
  assign f_s_dadda_rca16_and_2_10 = a[2] & b[10];
  assign f_s_dadda_rca16_and_1_11 = a[1] & b[11];
  assign f_s_dadda_rca16_and_0_12 = a[0] & b[12];
  assign f_s_dadda_rca16_fa43_xor0 = f_s_dadda_rca16_and_2_10 ^ f_s_dadda_rca16_and_1_11;
  assign f_s_dadda_rca16_fa43_and0 = f_s_dadda_rca16_and_2_10 & f_s_dadda_rca16_and_1_11;
  assign f_s_dadda_rca16_fa43_xor1 = f_s_dadda_rca16_fa43_xor0 ^ f_s_dadda_rca16_and_0_12;
  assign f_s_dadda_rca16_fa43_and1 = f_s_dadda_rca16_fa43_xor0 & f_s_dadda_rca16_and_0_12;
  assign f_s_dadda_rca16_fa43_or0 = f_s_dadda_rca16_fa43_and0 | f_s_dadda_rca16_fa43_and1;
  assign f_s_dadda_rca16_fa44_xor0 = f_s_dadda_rca16_fa37_xor1 ^ f_s_dadda_rca16_fa38_xor1;
  assign f_s_dadda_rca16_fa44_and0 = f_s_dadda_rca16_fa37_xor1 & f_s_dadda_rca16_fa38_xor1;
  assign f_s_dadda_rca16_fa44_xor1 = f_s_dadda_rca16_fa44_xor0 ^ f_s_dadda_rca16_fa39_xor1;
  assign f_s_dadda_rca16_fa44_and1 = f_s_dadda_rca16_fa44_xor0 & f_s_dadda_rca16_fa39_xor1;
  assign f_s_dadda_rca16_fa44_or0 = f_s_dadda_rca16_fa44_and0 | f_s_dadda_rca16_fa44_and1;
  assign f_s_dadda_rca16_ha11_xor0 = f_s_dadda_rca16_fa40_xor1 ^ f_s_dadda_rca16_fa41_xor1;
  assign f_s_dadda_rca16_ha11_and0 = f_s_dadda_rca16_fa40_xor1 & f_s_dadda_rca16_fa41_xor1;
  assign f_s_dadda_rca16_fa45_xor0 = f_s_dadda_rca16_ha11_and0 ^ f_s_dadda_rca16_fa44_or0;
  assign f_s_dadda_rca16_fa45_and0 = f_s_dadda_rca16_ha11_and0 & f_s_dadda_rca16_fa44_or0;
  assign f_s_dadda_rca16_fa45_xor1 = f_s_dadda_rca16_fa45_xor0 ^ f_s_dadda_rca16_fa43_or0;
  assign f_s_dadda_rca16_fa45_and1 = f_s_dadda_rca16_fa45_xor0 & f_s_dadda_rca16_fa43_or0;
  assign f_s_dadda_rca16_fa45_or0 = f_s_dadda_rca16_fa45_and0 | f_s_dadda_rca16_fa45_and1;
  assign f_s_dadda_rca16_fa46_xor0 = f_s_dadda_rca16_fa42_or0 ^ f_s_dadda_rca16_fa41_or0;
  assign f_s_dadda_rca16_fa46_and0 = f_s_dadda_rca16_fa42_or0 & f_s_dadda_rca16_fa41_or0;
  assign f_s_dadda_rca16_fa46_xor1 = f_s_dadda_rca16_fa46_xor0 ^ f_s_dadda_rca16_fa40_or0;
  assign f_s_dadda_rca16_fa46_and1 = f_s_dadda_rca16_fa46_xor0 & f_s_dadda_rca16_fa40_or0;
  assign f_s_dadda_rca16_fa46_or0 = f_s_dadda_rca16_fa46_and0 | f_s_dadda_rca16_fa46_and1;
  assign f_s_dadda_rca16_fa47_xor0 = f_s_dadda_rca16_fa39_or0 ^ f_s_dadda_rca16_fa38_or0;
  assign f_s_dadda_rca16_fa47_and0 = f_s_dadda_rca16_fa39_or0 & f_s_dadda_rca16_fa38_or0;
  assign f_s_dadda_rca16_fa47_xor1 = f_s_dadda_rca16_fa47_xor0 ^ f_s_dadda_rca16_fa37_or0;
  assign f_s_dadda_rca16_fa47_and1 = f_s_dadda_rca16_fa47_xor0 & f_s_dadda_rca16_fa37_or0;
  assign f_s_dadda_rca16_fa47_or0 = f_s_dadda_rca16_fa47_and0 | f_s_dadda_rca16_fa47_and1;
  assign f_s_dadda_rca16_and_11_2 = a[11] & b[2];
  assign f_s_dadda_rca16_and_10_3 = a[10] & b[3];
  assign f_s_dadda_rca16_and_9_4 = a[9] & b[4];
  assign f_s_dadda_rca16_fa48_xor0 = f_s_dadda_rca16_and_11_2 ^ f_s_dadda_rca16_and_10_3;
  assign f_s_dadda_rca16_fa48_and0 = f_s_dadda_rca16_and_11_2 & f_s_dadda_rca16_and_10_3;
  assign f_s_dadda_rca16_fa48_xor1 = f_s_dadda_rca16_fa48_xor0 ^ f_s_dadda_rca16_and_9_4;
  assign f_s_dadda_rca16_fa48_and1 = f_s_dadda_rca16_fa48_xor0 & f_s_dadda_rca16_and_9_4;
  assign f_s_dadda_rca16_fa48_or0 = f_s_dadda_rca16_fa48_and0 | f_s_dadda_rca16_fa48_and1;
  assign f_s_dadda_rca16_and_8_5 = a[8] & b[5];
  assign f_s_dadda_rca16_and_7_6 = a[7] & b[6];
  assign f_s_dadda_rca16_and_6_7 = a[6] & b[7];
  assign f_s_dadda_rca16_fa49_xor0 = f_s_dadda_rca16_and_8_5 ^ f_s_dadda_rca16_and_7_6;
  assign f_s_dadda_rca16_fa49_and0 = f_s_dadda_rca16_and_8_5 & f_s_dadda_rca16_and_7_6;
  assign f_s_dadda_rca16_fa49_xor1 = f_s_dadda_rca16_fa49_xor0 ^ f_s_dadda_rca16_and_6_7;
  assign f_s_dadda_rca16_fa49_and1 = f_s_dadda_rca16_fa49_xor0 & f_s_dadda_rca16_and_6_7;
  assign f_s_dadda_rca16_fa49_or0 = f_s_dadda_rca16_fa49_and0 | f_s_dadda_rca16_fa49_and1;
  assign f_s_dadda_rca16_and_5_8 = a[5] & b[8];
  assign f_s_dadda_rca16_and_4_9 = a[4] & b[9];
  assign f_s_dadda_rca16_and_3_10 = a[3] & b[10];
  assign f_s_dadda_rca16_fa50_xor0 = f_s_dadda_rca16_and_5_8 ^ f_s_dadda_rca16_and_4_9;
  assign f_s_dadda_rca16_fa50_and0 = f_s_dadda_rca16_and_5_8 & f_s_dadda_rca16_and_4_9;
  assign f_s_dadda_rca16_fa50_xor1 = f_s_dadda_rca16_fa50_xor0 ^ f_s_dadda_rca16_and_3_10;
  assign f_s_dadda_rca16_fa50_and1 = f_s_dadda_rca16_fa50_xor0 & f_s_dadda_rca16_and_3_10;
  assign f_s_dadda_rca16_fa50_or0 = f_s_dadda_rca16_fa50_and0 | f_s_dadda_rca16_fa50_and1;
  assign f_s_dadda_rca16_and_2_11 = a[2] & b[11];
  assign f_s_dadda_rca16_and_1_12 = a[1] & b[12];
  assign f_s_dadda_rca16_and_0_13 = a[0] & b[13];
  assign f_s_dadda_rca16_fa51_xor0 = f_s_dadda_rca16_and_2_11 ^ f_s_dadda_rca16_and_1_12;
  assign f_s_dadda_rca16_fa51_and0 = f_s_dadda_rca16_and_2_11 & f_s_dadda_rca16_and_1_12;
  assign f_s_dadda_rca16_fa51_xor1 = f_s_dadda_rca16_fa51_xor0 ^ f_s_dadda_rca16_and_0_13;
  assign f_s_dadda_rca16_fa51_and1 = f_s_dadda_rca16_fa51_xor0 & f_s_dadda_rca16_and_0_13;
  assign f_s_dadda_rca16_fa51_or0 = f_s_dadda_rca16_fa51_and0 | f_s_dadda_rca16_fa51_and1;
  assign f_s_dadda_rca16_fa52_xor0 = f_s_dadda_rca16_ha0_xor0 ^ f_s_dadda_rca16_fa45_xor1;
  assign f_s_dadda_rca16_fa52_and0 = f_s_dadda_rca16_ha0_xor0 & f_s_dadda_rca16_fa45_xor1;
  assign f_s_dadda_rca16_fa52_xor1 = f_s_dadda_rca16_fa52_xor0 ^ f_s_dadda_rca16_fa46_xor1;
  assign f_s_dadda_rca16_fa52_and1 = f_s_dadda_rca16_fa52_xor0 & f_s_dadda_rca16_fa46_xor1;
  assign f_s_dadda_rca16_fa52_or0 = f_s_dadda_rca16_fa52_and0 | f_s_dadda_rca16_fa52_and1;
  assign f_s_dadda_rca16_fa53_xor0 = f_s_dadda_rca16_fa47_xor1 ^ f_s_dadda_rca16_fa48_xor1;
  assign f_s_dadda_rca16_fa53_and0 = f_s_dadda_rca16_fa47_xor1 & f_s_dadda_rca16_fa48_xor1;
  assign f_s_dadda_rca16_fa53_xor1 = f_s_dadda_rca16_fa53_xor0 ^ f_s_dadda_rca16_fa49_xor1;
  assign f_s_dadda_rca16_fa53_and1 = f_s_dadda_rca16_fa53_xor0 & f_s_dadda_rca16_fa49_xor1;
  assign f_s_dadda_rca16_fa53_or0 = f_s_dadda_rca16_fa53_and0 | f_s_dadda_rca16_fa53_and1;
  assign f_s_dadda_rca16_fa54_xor0 = f_s_dadda_rca16_fa53_or0 ^ f_s_dadda_rca16_fa52_or0;
  assign f_s_dadda_rca16_fa54_and0 = f_s_dadda_rca16_fa53_or0 & f_s_dadda_rca16_fa52_or0;
  assign f_s_dadda_rca16_fa54_xor1 = f_s_dadda_rca16_fa54_xor0 ^ f_s_dadda_rca16_fa51_or0;
  assign f_s_dadda_rca16_fa54_and1 = f_s_dadda_rca16_fa54_xor0 & f_s_dadda_rca16_fa51_or0;
  assign f_s_dadda_rca16_fa54_or0 = f_s_dadda_rca16_fa54_and0 | f_s_dadda_rca16_fa54_and1;
  assign f_s_dadda_rca16_fa55_xor0 = f_s_dadda_rca16_fa50_or0 ^ f_s_dadda_rca16_fa49_or0;
  assign f_s_dadda_rca16_fa55_and0 = f_s_dadda_rca16_fa50_or0 & f_s_dadda_rca16_fa49_or0;
  assign f_s_dadda_rca16_fa55_xor1 = f_s_dadda_rca16_fa55_xor0 ^ f_s_dadda_rca16_fa48_or0;
  assign f_s_dadda_rca16_fa55_and1 = f_s_dadda_rca16_fa55_xor0 & f_s_dadda_rca16_fa48_or0;
  assign f_s_dadda_rca16_fa55_or0 = f_s_dadda_rca16_fa55_and0 | f_s_dadda_rca16_fa55_and1;
  assign f_s_dadda_rca16_fa56_xor0 = f_s_dadda_rca16_fa47_or0 ^ f_s_dadda_rca16_fa46_or0;
  assign f_s_dadda_rca16_fa56_and0 = f_s_dadda_rca16_fa47_or0 & f_s_dadda_rca16_fa46_or0;
  assign f_s_dadda_rca16_fa56_xor1 = f_s_dadda_rca16_fa56_xor0 ^ f_s_dadda_rca16_fa45_or0;
  assign f_s_dadda_rca16_fa56_and1 = f_s_dadda_rca16_fa56_xor0 & f_s_dadda_rca16_fa45_or0;
  assign f_s_dadda_rca16_fa56_or0 = f_s_dadda_rca16_fa56_and0 | f_s_dadda_rca16_fa56_and1;
  assign f_s_dadda_rca16_and_10_4 = a[10] & b[4];
  assign f_s_dadda_rca16_and_9_5 = a[9] & b[5];
  assign f_s_dadda_rca16_and_8_6 = a[8] & b[6];
  assign f_s_dadda_rca16_fa57_xor0 = f_s_dadda_rca16_and_10_4 ^ f_s_dadda_rca16_and_9_5;
  assign f_s_dadda_rca16_fa57_and0 = f_s_dadda_rca16_and_10_4 & f_s_dadda_rca16_and_9_5;
  assign f_s_dadda_rca16_fa57_xor1 = f_s_dadda_rca16_fa57_xor0 ^ f_s_dadda_rca16_and_8_6;
  assign f_s_dadda_rca16_fa57_and1 = f_s_dadda_rca16_fa57_xor0 & f_s_dadda_rca16_and_8_6;
  assign f_s_dadda_rca16_fa57_or0 = f_s_dadda_rca16_fa57_and0 | f_s_dadda_rca16_fa57_and1;
  assign f_s_dadda_rca16_and_7_7 = a[7] & b[7];
  assign f_s_dadda_rca16_and_6_8 = a[6] & b[8];
  assign f_s_dadda_rca16_and_5_9 = a[5] & b[9];
  assign f_s_dadda_rca16_fa58_xor0 = f_s_dadda_rca16_and_7_7 ^ f_s_dadda_rca16_and_6_8;
  assign f_s_dadda_rca16_fa58_and0 = f_s_dadda_rca16_and_7_7 & f_s_dadda_rca16_and_6_8;
  assign f_s_dadda_rca16_fa58_xor1 = f_s_dadda_rca16_fa58_xor0 ^ f_s_dadda_rca16_and_5_9;
  assign f_s_dadda_rca16_fa58_and1 = f_s_dadda_rca16_fa58_xor0 & f_s_dadda_rca16_and_5_9;
  assign f_s_dadda_rca16_fa58_or0 = f_s_dadda_rca16_fa58_and0 | f_s_dadda_rca16_fa58_and1;
  assign f_s_dadda_rca16_and_4_10 = a[4] & b[10];
  assign f_s_dadda_rca16_and_3_11 = a[3] & b[11];
  assign f_s_dadda_rca16_and_2_12 = a[2] & b[12];
  assign f_s_dadda_rca16_fa59_xor0 = f_s_dadda_rca16_and_4_10 ^ f_s_dadda_rca16_and_3_11;
  assign f_s_dadda_rca16_fa59_and0 = f_s_dadda_rca16_and_4_10 & f_s_dadda_rca16_and_3_11;
  assign f_s_dadda_rca16_fa59_xor1 = f_s_dadda_rca16_fa59_xor0 ^ f_s_dadda_rca16_and_2_12;
  assign f_s_dadda_rca16_fa59_and1 = f_s_dadda_rca16_fa59_xor0 & f_s_dadda_rca16_and_2_12;
  assign f_s_dadda_rca16_fa59_or0 = f_s_dadda_rca16_fa59_and0 | f_s_dadda_rca16_fa59_and1;
  assign f_s_dadda_rca16_and_1_13 = a[1] & b[13];
  assign f_s_dadda_rca16_and_0_14 = a[0] & b[14];
  assign f_s_dadda_rca16_fa60_xor0 = f_s_dadda_rca16_and_1_13 ^ f_s_dadda_rca16_and_0_14;
  assign f_s_dadda_rca16_fa60_and0 = f_s_dadda_rca16_and_1_13 & f_s_dadda_rca16_and_0_14;
  assign f_s_dadda_rca16_fa60_xor1 = f_s_dadda_rca16_fa60_xor0 ^ f_s_dadda_rca16_fa0_xor1;
  assign f_s_dadda_rca16_fa60_and1 = f_s_dadda_rca16_fa60_xor0 & f_s_dadda_rca16_fa0_xor1;
  assign f_s_dadda_rca16_fa60_or0 = f_s_dadda_rca16_fa60_and0 | f_s_dadda_rca16_fa60_and1;
  assign f_s_dadda_rca16_fa61_xor0 = f_s_dadda_rca16_ha1_xor0 ^ f_s_dadda_rca16_fa54_xor1;
  assign f_s_dadda_rca16_fa61_and0 = f_s_dadda_rca16_ha1_xor0 & f_s_dadda_rca16_fa54_xor1;
  assign f_s_dadda_rca16_fa61_xor1 = f_s_dadda_rca16_fa61_xor0 ^ f_s_dadda_rca16_fa55_xor1;
  assign f_s_dadda_rca16_fa61_and1 = f_s_dadda_rca16_fa61_xor0 & f_s_dadda_rca16_fa55_xor1;
  assign f_s_dadda_rca16_fa61_or0 = f_s_dadda_rca16_fa61_and0 | f_s_dadda_rca16_fa61_and1;
  assign f_s_dadda_rca16_fa62_xor0 = f_s_dadda_rca16_fa56_xor1 ^ f_s_dadda_rca16_fa57_xor1;
  assign f_s_dadda_rca16_fa62_and0 = f_s_dadda_rca16_fa56_xor1 & f_s_dadda_rca16_fa57_xor1;
  assign f_s_dadda_rca16_fa62_xor1 = f_s_dadda_rca16_fa62_xor0 ^ f_s_dadda_rca16_fa58_xor1;
  assign f_s_dadda_rca16_fa62_and1 = f_s_dadda_rca16_fa62_xor0 & f_s_dadda_rca16_fa58_xor1;
  assign f_s_dadda_rca16_fa62_or0 = f_s_dadda_rca16_fa62_and0 | f_s_dadda_rca16_fa62_and1;
  assign f_s_dadda_rca16_fa63_xor0 = f_s_dadda_rca16_fa62_or0 ^ f_s_dadda_rca16_fa61_or0;
  assign f_s_dadda_rca16_fa63_and0 = f_s_dadda_rca16_fa62_or0 & f_s_dadda_rca16_fa61_or0;
  assign f_s_dadda_rca16_fa63_xor1 = f_s_dadda_rca16_fa63_xor0 ^ f_s_dadda_rca16_fa60_or0;
  assign f_s_dadda_rca16_fa63_and1 = f_s_dadda_rca16_fa63_xor0 & f_s_dadda_rca16_fa60_or0;
  assign f_s_dadda_rca16_fa63_or0 = f_s_dadda_rca16_fa63_and0 | f_s_dadda_rca16_fa63_and1;
  assign f_s_dadda_rca16_fa64_xor0 = f_s_dadda_rca16_fa59_or0 ^ f_s_dadda_rca16_fa58_or0;
  assign f_s_dadda_rca16_fa64_and0 = f_s_dadda_rca16_fa59_or0 & f_s_dadda_rca16_fa58_or0;
  assign f_s_dadda_rca16_fa64_xor1 = f_s_dadda_rca16_fa64_xor0 ^ f_s_dadda_rca16_fa57_or0;
  assign f_s_dadda_rca16_fa64_and1 = f_s_dadda_rca16_fa64_xor0 & f_s_dadda_rca16_fa57_or0;
  assign f_s_dadda_rca16_fa64_or0 = f_s_dadda_rca16_fa64_and0 | f_s_dadda_rca16_fa64_and1;
  assign f_s_dadda_rca16_fa65_xor0 = f_s_dadda_rca16_fa56_or0 ^ f_s_dadda_rca16_fa55_or0;
  assign f_s_dadda_rca16_fa65_and0 = f_s_dadda_rca16_fa56_or0 & f_s_dadda_rca16_fa55_or0;
  assign f_s_dadda_rca16_fa65_xor1 = f_s_dadda_rca16_fa65_xor0 ^ f_s_dadda_rca16_fa54_or0;
  assign f_s_dadda_rca16_fa65_and1 = f_s_dadda_rca16_fa65_xor0 & f_s_dadda_rca16_fa54_or0;
  assign f_s_dadda_rca16_fa65_or0 = f_s_dadda_rca16_fa65_and0 | f_s_dadda_rca16_fa65_and1;
  assign f_s_dadda_rca16_and_9_6 = a[9] & b[6];
  assign f_s_dadda_rca16_and_8_7 = a[8] & b[7];
  assign f_s_dadda_rca16_and_7_8 = a[7] & b[8];
  assign f_s_dadda_rca16_fa66_xor0 = f_s_dadda_rca16_and_9_6 ^ f_s_dadda_rca16_and_8_7;
  assign f_s_dadda_rca16_fa66_and0 = f_s_dadda_rca16_and_9_6 & f_s_dadda_rca16_and_8_7;
  assign f_s_dadda_rca16_fa66_xor1 = f_s_dadda_rca16_fa66_xor0 ^ f_s_dadda_rca16_and_7_8;
  assign f_s_dadda_rca16_fa66_and1 = f_s_dadda_rca16_fa66_xor0 & f_s_dadda_rca16_and_7_8;
  assign f_s_dadda_rca16_fa66_or0 = f_s_dadda_rca16_fa66_and0 | f_s_dadda_rca16_fa66_and1;
  assign f_s_dadda_rca16_and_6_9 = a[6] & b[9];
  assign f_s_dadda_rca16_and_5_10 = a[5] & b[10];
  assign f_s_dadda_rca16_and_4_11 = a[4] & b[11];
  assign f_s_dadda_rca16_fa67_xor0 = f_s_dadda_rca16_and_6_9 ^ f_s_dadda_rca16_and_5_10;
  assign f_s_dadda_rca16_fa67_and0 = f_s_dadda_rca16_and_6_9 & f_s_dadda_rca16_and_5_10;
  assign f_s_dadda_rca16_fa67_xor1 = f_s_dadda_rca16_fa67_xor0 ^ f_s_dadda_rca16_and_4_11;
  assign f_s_dadda_rca16_fa67_and1 = f_s_dadda_rca16_fa67_xor0 & f_s_dadda_rca16_and_4_11;
  assign f_s_dadda_rca16_fa67_or0 = f_s_dadda_rca16_fa67_and0 | f_s_dadda_rca16_fa67_and1;
  assign f_s_dadda_rca16_and_3_12 = a[3] & b[12];
  assign f_s_dadda_rca16_and_2_13 = a[2] & b[13];
  assign f_s_dadda_rca16_and_1_14 = a[1] & b[14];
  assign f_s_dadda_rca16_fa68_xor0 = f_s_dadda_rca16_and_3_12 ^ f_s_dadda_rca16_and_2_13;
  assign f_s_dadda_rca16_fa68_and0 = f_s_dadda_rca16_and_3_12 & f_s_dadda_rca16_and_2_13;
  assign f_s_dadda_rca16_fa68_xor1 = f_s_dadda_rca16_fa68_xor0 ^ f_s_dadda_rca16_and_1_14;
  assign f_s_dadda_rca16_fa68_and1 = f_s_dadda_rca16_fa68_xor0 & f_s_dadda_rca16_and_1_14;
  assign f_s_dadda_rca16_fa68_or0 = f_s_dadda_rca16_fa68_and0 | f_s_dadda_rca16_fa68_and1;
  assign f_s_dadda_rca16_nand_0_15 = ~(a[0] & b[15]);
  assign f_s_dadda_rca16_fa69_xor0 = f_s_dadda_rca16_nand_0_15 ^ f_s_dadda_rca16_fa1_xor1;
  assign f_s_dadda_rca16_fa69_and0 = f_s_dadda_rca16_nand_0_15 & f_s_dadda_rca16_fa1_xor1;
  assign f_s_dadda_rca16_fa69_xor1 = f_s_dadda_rca16_fa69_xor0 ^ f_s_dadda_rca16_fa2_xor1;
  assign f_s_dadda_rca16_fa69_and1 = f_s_dadda_rca16_fa69_xor0 & f_s_dadda_rca16_fa2_xor1;
  assign f_s_dadda_rca16_fa69_or0 = f_s_dadda_rca16_fa69_and0 | f_s_dadda_rca16_fa69_and1;
  assign f_s_dadda_rca16_fa70_xor0 = f_s_dadda_rca16_ha2_xor0 ^ f_s_dadda_rca16_fa63_xor1;
  assign f_s_dadda_rca16_fa70_and0 = f_s_dadda_rca16_ha2_xor0 & f_s_dadda_rca16_fa63_xor1;
  assign f_s_dadda_rca16_fa70_xor1 = f_s_dadda_rca16_fa70_xor0 ^ f_s_dadda_rca16_fa64_xor1;
  assign f_s_dadda_rca16_fa70_and1 = f_s_dadda_rca16_fa70_xor0 & f_s_dadda_rca16_fa64_xor1;
  assign f_s_dadda_rca16_fa70_or0 = f_s_dadda_rca16_fa70_and0 | f_s_dadda_rca16_fa70_and1;
  assign f_s_dadda_rca16_fa71_xor0 = f_s_dadda_rca16_fa65_xor1 ^ f_s_dadda_rca16_fa66_xor1;
  assign f_s_dadda_rca16_fa71_and0 = f_s_dadda_rca16_fa65_xor1 & f_s_dadda_rca16_fa66_xor1;
  assign f_s_dadda_rca16_fa71_xor1 = f_s_dadda_rca16_fa71_xor0 ^ f_s_dadda_rca16_fa67_xor1;
  assign f_s_dadda_rca16_fa71_and1 = f_s_dadda_rca16_fa71_xor0 & f_s_dadda_rca16_fa67_xor1;
  assign f_s_dadda_rca16_fa71_or0 = f_s_dadda_rca16_fa71_and0 | f_s_dadda_rca16_fa71_and1;
  assign f_s_dadda_rca16_fa72_xor0 = f_s_dadda_rca16_fa71_or0 ^ f_s_dadda_rca16_fa70_or0;
  assign f_s_dadda_rca16_fa72_and0 = f_s_dadda_rca16_fa71_or0 & f_s_dadda_rca16_fa70_or0;
  assign f_s_dadda_rca16_fa72_xor1 = f_s_dadda_rca16_fa72_xor0 ^ f_s_dadda_rca16_fa69_or0;
  assign f_s_dadda_rca16_fa72_and1 = f_s_dadda_rca16_fa72_xor0 & f_s_dadda_rca16_fa69_or0;
  assign f_s_dadda_rca16_fa72_or0 = f_s_dadda_rca16_fa72_and0 | f_s_dadda_rca16_fa72_and1;
  assign f_s_dadda_rca16_fa73_xor0 = f_s_dadda_rca16_fa68_or0 ^ f_s_dadda_rca16_fa67_or0;
  assign f_s_dadda_rca16_fa73_and0 = f_s_dadda_rca16_fa68_or0 & f_s_dadda_rca16_fa67_or0;
  assign f_s_dadda_rca16_fa73_xor1 = f_s_dadda_rca16_fa73_xor0 ^ f_s_dadda_rca16_fa66_or0;
  assign f_s_dadda_rca16_fa73_and1 = f_s_dadda_rca16_fa73_xor0 & f_s_dadda_rca16_fa66_or0;
  assign f_s_dadda_rca16_fa73_or0 = f_s_dadda_rca16_fa73_and0 | f_s_dadda_rca16_fa73_and1;
  assign f_s_dadda_rca16_fa74_xor0 = f_s_dadda_rca16_fa65_or0 ^ f_s_dadda_rca16_fa64_or0;
  assign f_s_dadda_rca16_fa74_and0 = f_s_dadda_rca16_fa65_or0 & f_s_dadda_rca16_fa64_or0;
  assign f_s_dadda_rca16_fa74_xor1 = f_s_dadda_rca16_fa74_xor0 ^ f_s_dadda_rca16_fa63_or0;
  assign f_s_dadda_rca16_fa74_and1 = f_s_dadda_rca16_fa74_xor0 & f_s_dadda_rca16_fa63_or0;
  assign f_s_dadda_rca16_fa74_or0 = f_s_dadda_rca16_fa74_and0 | f_s_dadda_rca16_fa74_and1;
  assign f_s_dadda_rca16_and_10_6 = a[10] & b[6];
  assign f_s_dadda_rca16_and_9_7 = a[9] & b[7];
  assign f_s_dadda_rca16_and_8_8 = a[8] & b[8];
  assign f_s_dadda_rca16_fa75_xor0 = f_s_dadda_rca16_and_10_6 ^ f_s_dadda_rca16_and_9_7;
  assign f_s_dadda_rca16_fa75_and0 = f_s_dadda_rca16_and_10_6 & f_s_dadda_rca16_and_9_7;
  assign f_s_dadda_rca16_fa75_xor1 = f_s_dadda_rca16_fa75_xor0 ^ f_s_dadda_rca16_and_8_8;
  assign f_s_dadda_rca16_fa75_and1 = f_s_dadda_rca16_fa75_xor0 & f_s_dadda_rca16_and_8_8;
  assign f_s_dadda_rca16_fa75_or0 = f_s_dadda_rca16_fa75_and0 | f_s_dadda_rca16_fa75_and1;
  assign f_s_dadda_rca16_and_7_9 = a[7] & b[9];
  assign f_s_dadda_rca16_and_6_10 = a[6] & b[10];
  assign f_s_dadda_rca16_and_5_11 = a[5] & b[11];
  assign f_s_dadda_rca16_fa76_xor0 = f_s_dadda_rca16_and_7_9 ^ f_s_dadda_rca16_and_6_10;
  assign f_s_dadda_rca16_fa76_and0 = f_s_dadda_rca16_and_7_9 & f_s_dadda_rca16_and_6_10;
  assign f_s_dadda_rca16_fa76_xor1 = f_s_dadda_rca16_fa76_xor0 ^ f_s_dadda_rca16_and_5_11;
  assign f_s_dadda_rca16_fa76_and1 = f_s_dadda_rca16_fa76_xor0 & f_s_dadda_rca16_and_5_11;
  assign f_s_dadda_rca16_fa76_or0 = f_s_dadda_rca16_fa76_and0 | f_s_dadda_rca16_fa76_and1;
  assign f_s_dadda_rca16_and_4_12 = a[4] & b[12];
  assign f_s_dadda_rca16_and_3_13 = a[3] & b[13];
  assign f_s_dadda_rca16_and_2_14 = a[2] & b[14];
  assign f_s_dadda_rca16_fa77_xor0 = f_s_dadda_rca16_and_4_12 ^ f_s_dadda_rca16_and_3_13;
  assign f_s_dadda_rca16_fa77_and0 = f_s_dadda_rca16_and_4_12 & f_s_dadda_rca16_and_3_13;
  assign f_s_dadda_rca16_fa77_xor1 = f_s_dadda_rca16_fa77_xor0 ^ f_s_dadda_rca16_and_2_14;
  assign f_s_dadda_rca16_fa77_and1 = f_s_dadda_rca16_fa77_xor0 & f_s_dadda_rca16_and_2_14;
  assign f_s_dadda_rca16_fa77_or0 = f_s_dadda_rca16_fa77_and0 | f_s_dadda_rca16_fa77_and1;
  assign f_s_dadda_rca16_nand_1_15 = ~(a[1] & b[15]);
  assign f_s_dadda_rca16_fa78_xor0 = f_s_dadda_rca16_nand_1_15 ^ f_s_dadda_rca16_fa3_xor1;
  assign f_s_dadda_rca16_fa78_and0 = f_s_dadda_rca16_nand_1_15 & f_s_dadda_rca16_fa3_xor1;
  assign f_s_dadda_rca16_fa78_xor1 = f_s_dadda_rca16_fa78_xor0 ^ f_s_dadda_rca16_fa4_xor1;
  assign f_s_dadda_rca16_fa78_and1 = f_s_dadda_rca16_fa78_xor0 & f_s_dadda_rca16_fa4_xor1;
  assign f_s_dadda_rca16_fa78_or0 = f_s_dadda_rca16_fa78_and0 | f_s_dadda_rca16_fa78_and1;
  assign f_s_dadda_rca16_fa79_xor0 = f_s_dadda_rca16_fa5_xor1 ^ f_s_dadda_rca16_fa72_xor1;
  assign f_s_dadda_rca16_fa79_and0 = f_s_dadda_rca16_fa5_xor1 & f_s_dadda_rca16_fa72_xor1;
  assign f_s_dadda_rca16_fa79_xor1 = f_s_dadda_rca16_fa79_xor0 ^ f_s_dadda_rca16_fa73_xor1;
  assign f_s_dadda_rca16_fa79_and1 = f_s_dadda_rca16_fa79_xor0 & f_s_dadda_rca16_fa73_xor1;
  assign f_s_dadda_rca16_fa79_or0 = f_s_dadda_rca16_fa79_and0 | f_s_dadda_rca16_fa79_and1;
  assign f_s_dadda_rca16_fa80_xor0 = f_s_dadda_rca16_fa74_xor1 ^ f_s_dadda_rca16_fa75_xor1;
  assign f_s_dadda_rca16_fa80_and0 = f_s_dadda_rca16_fa74_xor1 & f_s_dadda_rca16_fa75_xor1;
  assign f_s_dadda_rca16_fa80_xor1 = f_s_dadda_rca16_fa80_xor0 ^ f_s_dadda_rca16_fa76_xor1;
  assign f_s_dadda_rca16_fa80_and1 = f_s_dadda_rca16_fa80_xor0 & f_s_dadda_rca16_fa76_xor1;
  assign f_s_dadda_rca16_fa80_or0 = f_s_dadda_rca16_fa80_and0 | f_s_dadda_rca16_fa80_and1;
  assign f_s_dadda_rca16_fa81_xor0 = f_s_dadda_rca16_fa80_or0 ^ f_s_dadda_rca16_fa79_or0;
  assign f_s_dadda_rca16_fa81_and0 = f_s_dadda_rca16_fa80_or0 & f_s_dadda_rca16_fa79_or0;
  assign f_s_dadda_rca16_fa81_xor1 = f_s_dadda_rca16_fa81_xor0 ^ f_s_dadda_rca16_fa78_or0;
  assign f_s_dadda_rca16_fa81_and1 = f_s_dadda_rca16_fa81_xor0 & f_s_dadda_rca16_fa78_or0;
  assign f_s_dadda_rca16_fa81_or0 = f_s_dadda_rca16_fa81_and0 | f_s_dadda_rca16_fa81_and1;
  assign f_s_dadda_rca16_fa82_xor0 = f_s_dadda_rca16_fa77_or0 ^ f_s_dadda_rca16_fa76_or0;
  assign f_s_dadda_rca16_fa82_and0 = f_s_dadda_rca16_fa77_or0 & f_s_dadda_rca16_fa76_or0;
  assign f_s_dadda_rca16_fa82_xor1 = f_s_dadda_rca16_fa82_xor0 ^ f_s_dadda_rca16_fa75_or0;
  assign f_s_dadda_rca16_fa82_and1 = f_s_dadda_rca16_fa82_xor0 & f_s_dadda_rca16_fa75_or0;
  assign f_s_dadda_rca16_fa82_or0 = f_s_dadda_rca16_fa82_and0 | f_s_dadda_rca16_fa82_and1;
  assign f_s_dadda_rca16_fa83_xor0 = f_s_dadda_rca16_fa74_or0 ^ f_s_dadda_rca16_fa73_or0;
  assign f_s_dadda_rca16_fa83_and0 = f_s_dadda_rca16_fa74_or0 & f_s_dadda_rca16_fa73_or0;
  assign f_s_dadda_rca16_fa83_xor1 = f_s_dadda_rca16_fa83_xor0 ^ f_s_dadda_rca16_fa72_or0;
  assign f_s_dadda_rca16_fa83_and1 = f_s_dadda_rca16_fa83_xor0 & f_s_dadda_rca16_fa72_or0;
  assign f_s_dadda_rca16_fa83_or0 = f_s_dadda_rca16_fa83_and0 | f_s_dadda_rca16_fa83_and1;
  assign f_s_dadda_rca16_and_12_5 = a[12] & b[5];
  assign f_s_dadda_rca16_and_11_6 = a[11] & b[6];
  assign f_s_dadda_rca16_and_10_7 = a[10] & b[7];
  assign f_s_dadda_rca16_fa84_xor0 = f_s_dadda_rca16_and_12_5 ^ f_s_dadda_rca16_and_11_6;
  assign f_s_dadda_rca16_fa84_and0 = f_s_dadda_rca16_and_12_5 & f_s_dadda_rca16_and_11_6;
  assign f_s_dadda_rca16_fa84_xor1 = f_s_dadda_rca16_fa84_xor0 ^ f_s_dadda_rca16_and_10_7;
  assign f_s_dadda_rca16_fa84_and1 = f_s_dadda_rca16_fa84_xor0 & f_s_dadda_rca16_and_10_7;
  assign f_s_dadda_rca16_fa84_or0 = f_s_dadda_rca16_fa84_and0 | f_s_dadda_rca16_fa84_and1;
  assign f_s_dadda_rca16_and_9_8 = a[9] & b[8];
  assign f_s_dadda_rca16_and_8_9 = a[8] & b[9];
  assign f_s_dadda_rca16_and_7_10 = a[7] & b[10];
  assign f_s_dadda_rca16_fa85_xor0 = f_s_dadda_rca16_and_9_8 ^ f_s_dadda_rca16_and_8_9;
  assign f_s_dadda_rca16_fa85_and0 = f_s_dadda_rca16_and_9_8 & f_s_dadda_rca16_and_8_9;
  assign f_s_dadda_rca16_fa85_xor1 = f_s_dadda_rca16_fa85_xor0 ^ f_s_dadda_rca16_and_7_10;
  assign f_s_dadda_rca16_fa85_and1 = f_s_dadda_rca16_fa85_xor0 & f_s_dadda_rca16_and_7_10;
  assign f_s_dadda_rca16_fa85_or0 = f_s_dadda_rca16_fa85_and0 | f_s_dadda_rca16_fa85_and1;
  assign f_s_dadda_rca16_and_6_11 = a[6] & b[11];
  assign f_s_dadda_rca16_and_5_12 = a[5] & b[12];
  assign f_s_dadda_rca16_and_4_13 = a[4] & b[13];
  assign f_s_dadda_rca16_fa86_xor0 = f_s_dadda_rca16_and_6_11 ^ f_s_dadda_rca16_and_5_12;
  assign f_s_dadda_rca16_fa86_and0 = f_s_dadda_rca16_and_6_11 & f_s_dadda_rca16_and_5_12;
  assign f_s_dadda_rca16_fa86_xor1 = f_s_dadda_rca16_fa86_xor0 ^ f_s_dadda_rca16_and_4_13;
  assign f_s_dadda_rca16_fa86_and1 = f_s_dadda_rca16_fa86_xor0 & f_s_dadda_rca16_and_4_13;
  assign f_s_dadda_rca16_fa86_or0 = f_s_dadda_rca16_fa86_and0 | f_s_dadda_rca16_fa86_and1;
  assign f_s_dadda_rca16_and_3_14 = a[3] & b[14];
  assign f_s_dadda_rca16_nand_2_15 = ~(a[2] & b[15]);
  assign f_s_dadda_rca16_fa87_xor0 = f_s_dadda_rca16_and_3_14 ^ f_s_dadda_rca16_nand_2_15;
  assign f_s_dadda_rca16_fa87_and0 = f_s_dadda_rca16_and_3_14 & f_s_dadda_rca16_nand_2_15;
  assign f_s_dadda_rca16_fa87_xor1 = f_s_dadda_rca16_fa87_xor0 ^ f_s_dadda_rca16_fa6_xor1;
  assign f_s_dadda_rca16_fa87_and1 = f_s_dadda_rca16_fa87_xor0 & f_s_dadda_rca16_fa6_xor1;
  assign f_s_dadda_rca16_fa87_or0 = f_s_dadda_rca16_fa87_and0 | f_s_dadda_rca16_fa87_and1;
  assign f_s_dadda_rca16_fa88_xor0 = f_s_dadda_rca16_fa7_xor1 ^ f_s_dadda_rca16_fa81_xor1;
  assign f_s_dadda_rca16_fa88_and0 = f_s_dadda_rca16_fa7_xor1 & f_s_dadda_rca16_fa81_xor1;
  assign f_s_dadda_rca16_fa88_xor1 = f_s_dadda_rca16_fa88_xor0 ^ f_s_dadda_rca16_fa82_xor1;
  assign f_s_dadda_rca16_fa88_and1 = f_s_dadda_rca16_fa88_xor0 & f_s_dadda_rca16_fa82_xor1;
  assign f_s_dadda_rca16_fa88_or0 = f_s_dadda_rca16_fa88_and0 | f_s_dadda_rca16_fa88_and1;
  assign f_s_dadda_rca16_fa89_xor0 = f_s_dadda_rca16_fa83_xor1 ^ f_s_dadda_rca16_fa84_xor1;
  assign f_s_dadda_rca16_fa89_and0 = f_s_dadda_rca16_fa83_xor1 & f_s_dadda_rca16_fa84_xor1;
  assign f_s_dadda_rca16_fa89_xor1 = f_s_dadda_rca16_fa89_xor0 ^ f_s_dadda_rca16_fa85_xor1;
  assign f_s_dadda_rca16_fa89_and1 = f_s_dadda_rca16_fa89_xor0 & f_s_dadda_rca16_fa85_xor1;
  assign f_s_dadda_rca16_fa89_or0 = f_s_dadda_rca16_fa89_and0 | f_s_dadda_rca16_fa89_and1;
  assign f_s_dadda_rca16_fa90_xor0 = f_s_dadda_rca16_fa89_or0 ^ f_s_dadda_rca16_fa88_or0;
  assign f_s_dadda_rca16_fa90_and0 = f_s_dadda_rca16_fa89_or0 & f_s_dadda_rca16_fa88_or0;
  assign f_s_dadda_rca16_fa90_xor1 = f_s_dadda_rca16_fa90_xor0 ^ f_s_dadda_rca16_fa87_or0;
  assign f_s_dadda_rca16_fa90_and1 = f_s_dadda_rca16_fa90_xor0 & f_s_dadda_rca16_fa87_or0;
  assign f_s_dadda_rca16_fa90_or0 = f_s_dadda_rca16_fa90_and0 | f_s_dadda_rca16_fa90_and1;
  assign f_s_dadda_rca16_fa91_xor0 = f_s_dadda_rca16_fa86_or0 ^ f_s_dadda_rca16_fa85_or0;
  assign f_s_dadda_rca16_fa91_and0 = f_s_dadda_rca16_fa86_or0 & f_s_dadda_rca16_fa85_or0;
  assign f_s_dadda_rca16_fa91_xor1 = f_s_dadda_rca16_fa91_xor0 ^ f_s_dadda_rca16_fa84_or0;
  assign f_s_dadda_rca16_fa91_and1 = f_s_dadda_rca16_fa91_xor0 & f_s_dadda_rca16_fa84_or0;
  assign f_s_dadda_rca16_fa91_or0 = f_s_dadda_rca16_fa91_and0 | f_s_dadda_rca16_fa91_and1;
  assign f_s_dadda_rca16_fa92_xor0 = f_s_dadda_rca16_fa83_or0 ^ f_s_dadda_rca16_fa82_or0;
  assign f_s_dadda_rca16_fa92_and0 = f_s_dadda_rca16_fa83_or0 & f_s_dadda_rca16_fa82_or0;
  assign f_s_dadda_rca16_fa92_xor1 = f_s_dadda_rca16_fa92_xor0 ^ f_s_dadda_rca16_fa81_or0;
  assign f_s_dadda_rca16_fa92_and1 = f_s_dadda_rca16_fa92_xor0 & f_s_dadda_rca16_fa81_or0;
  assign f_s_dadda_rca16_fa92_or0 = f_s_dadda_rca16_fa92_and0 | f_s_dadda_rca16_fa92_and1;
  assign f_s_dadda_rca16_and_14_4 = a[14] & b[4];
  assign f_s_dadda_rca16_and_13_5 = a[13] & b[5];
  assign f_s_dadda_rca16_and_12_6 = a[12] & b[6];
  assign f_s_dadda_rca16_fa93_xor0 = f_s_dadda_rca16_and_14_4 ^ f_s_dadda_rca16_and_13_5;
  assign f_s_dadda_rca16_fa93_and0 = f_s_dadda_rca16_and_14_4 & f_s_dadda_rca16_and_13_5;
  assign f_s_dadda_rca16_fa93_xor1 = f_s_dadda_rca16_fa93_xor0 ^ f_s_dadda_rca16_and_12_6;
  assign f_s_dadda_rca16_fa93_and1 = f_s_dadda_rca16_fa93_xor0 & f_s_dadda_rca16_and_12_6;
  assign f_s_dadda_rca16_fa93_or0 = f_s_dadda_rca16_fa93_and0 | f_s_dadda_rca16_fa93_and1;
  assign f_s_dadda_rca16_and_11_7 = a[11] & b[7];
  assign f_s_dadda_rca16_and_10_8 = a[10] & b[8];
  assign f_s_dadda_rca16_and_9_9 = a[9] & b[9];
  assign f_s_dadda_rca16_fa94_xor0 = f_s_dadda_rca16_and_11_7 ^ f_s_dadda_rca16_and_10_8;
  assign f_s_dadda_rca16_fa94_and0 = f_s_dadda_rca16_and_11_7 & f_s_dadda_rca16_and_10_8;
  assign f_s_dadda_rca16_fa94_xor1 = f_s_dadda_rca16_fa94_xor0 ^ f_s_dadda_rca16_and_9_9;
  assign f_s_dadda_rca16_fa94_and1 = f_s_dadda_rca16_fa94_xor0 & f_s_dadda_rca16_and_9_9;
  assign f_s_dadda_rca16_fa94_or0 = f_s_dadda_rca16_fa94_and0 | f_s_dadda_rca16_fa94_and1;
  assign f_s_dadda_rca16_and_8_10 = a[8] & b[10];
  assign f_s_dadda_rca16_and_7_11 = a[7] & b[11];
  assign f_s_dadda_rca16_and_6_12 = a[6] & b[12];
  assign f_s_dadda_rca16_fa95_xor0 = f_s_dadda_rca16_and_8_10 ^ f_s_dadda_rca16_and_7_11;
  assign f_s_dadda_rca16_fa95_and0 = f_s_dadda_rca16_and_8_10 & f_s_dadda_rca16_and_7_11;
  assign f_s_dadda_rca16_fa95_xor1 = f_s_dadda_rca16_fa95_xor0 ^ f_s_dadda_rca16_and_6_12;
  assign f_s_dadda_rca16_fa95_and1 = f_s_dadda_rca16_fa95_xor0 & f_s_dadda_rca16_and_6_12;
  assign f_s_dadda_rca16_fa95_or0 = f_s_dadda_rca16_fa95_and0 | f_s_dadda_rca16_fa95_and1;
  assign f_s_dadda_rca16_and_5_13 = a[5] & b[13];
  assign f_s_dadda_rca16_and_4_14 = a[4] & b[14];
  assign f_s_dadda_rca16_nand_3_15 = ~(a[3] & b[15]);
  assign f_s_dadda_rca16_fa96_xor0 = f_s_dadda_rca16_and_5_13 ^ f_s_dadda_rca16_and_4_14;
  assign f_s_dadda_rca16_fa96_and0 = f_s_dadda_rca16_and_5_13 & f_s_dadda_rca16_and_4_14;
  assign f_s_dadda_rca16_fa96_xor1 = f_s_dadda_rca16_fa96_xor0 ^ f_s_dadda_rca16_nand_3_15;
  assign f_s_dadda_rca16_fa96_and1 = f_s_dadda_rca16_fa96_xor0 & f_s_dadda_rca16_nand_3_15;
  assign f_s_dadda_rca16_fa96_or0 = f_s_dadda_rca16_fa96_and0 | f_s_dadda_rca16_fa96_and1;
  assign f_s_dadda_rca16_fa97_xor0 = f_s_dadda_rca16_fa8_xor1 ^ f_s_dadda_rca16_fa90_xor1;
  assign f_s_dadda_rca16_fa97_and0 = f_s_dadda_rca16_fa8_xor1 & f_s_dadda_rca16_fa90_xor1;
  assign f_s_dadda_rca16_fa97_xor1 = f_s_dadda_rca16_fa97_xor0 ^ f_s_dadda_rca16_fa91_xor1;
  assign f_s_dadda_rca16_fa97_and1 = f_s_dadda_rca16_fa97_xor0 & f_s_dadda_rca16_fa91_xor1;
  assign f_s_dadda_rca16_fa97_or0 = f_s_dadda_rca16_fa97_and0 | f_s_dadda_rca16_fa97_and1;
  assign f_s_dadda_rca16_fa98_xor0 = f_s_dadda_rca16_fa92_xor1 ^ f_s_dadda_rca16_fa93_xor1;
  assign f_s_dadda_rca16_fa98_and0 = f_s_dadda_rca16_fa92_xor1 & f_s_dadda_rca16_fa93_xor1;
  assign f_s_dadda_rca16_fa98_xor1 = f_s_dadda_rca16_fa98_xor0 ^ f_s_dadda_rca16_fa94_xor1;
  assign f_s_dadda_rca16_fa98_and1 = f_s_dadda_rca16_fa98_xor0 & f_s_dadda_rca16_fa94_xor1;
  assign f_s_dadda_rca16_fa98_or0 = f_s_dadda_rca16_fa98_and0 | f_s_dadda_rca16_fa98_and1;
  assign f_s_dadda_rca16_fa99_xor0 = f_s_dadda_rca16_fa98_or0 ^ f_s_dadda_rca16_fa97_or0;
  assign f_s_dadda_rca16_fa99_and0 = f_s_dadda_rca16_fa98_or0 & f_s_dadda_rca16_fa97_or0;
  assign f_s_dadda_rca16_fa99_xor1 = f_s_dadda_rca16_fa99_xor0 ^ f_s_dadda_rca16_fa96_or0;
  assign f_s_dadda_rca16_fa99_and1 = f_s_dadda_rca16_fa99_xor0 & f_s_dadda_rca16_fa96_or0;
  assign f_s_dadda_rca16_fa99_or0 = f_s_dadda_rca16_fa99_and0 | f_s_dadda_rca16_fa99_and1;
  assign f_s_dadda_rca16_fa100_xor0 = f_s_dadda_rca16_fa95_or0 ^ f_s_dadda_rca16_fa94_or0;
  assign f_s_dadda_rca16_fa100_and0 = f_s_dadda_rca16_fa95_or0 & f_s_dadda_rca16_fa94_or0;
  assign f_s_dadda_rca16_fa100_xor1 = f_s_dadda_rca16_fa100_xor0 ^ f_s_dadda_rca16_fa93_or0;
  assign f_s_dadda_rca16_fa100_and1 = f_s_dadda_rca16_fa100_xor0 & f_s_dadda_rca16_fa93_or0;
  assign f_s_dadda_rca16_fa100_or0 = f_s_dadda_rca16_fa100_and0 | f_s_dadda_rca16_fa100_and1;
  assign f_s_dadda_rca16_fa101_xor0 = f_s_dadda_rca16_fa92_or0 ^ f_s_dadda_rca16_fa91_or0;
  assign f_s_dadda_rca16_fa101_and0 = f_s_dadda_rca16_fa92_or0 & f_s_dadda_rca16_fa91_or0;
  assign f_s_dadda_rca16_fa101_xor1 = f_s_dadda_rca16_fa101_xor0 ^ f_s_dadda_rca16_fa90_or0;
  assign f_s_dadda_rca16_fa101_and1 = f_s_dadda_rca16_fa101_xor0 & f_s_dadda_rca16_fa90_or0;
  assign f_s_dadda_rca16_fa101_or0 = f_s_dadda_rca16_fa101_and0 | f_s_dadda_rca16_fa101_and1;
  assign f_s_dadda_rca16_nand_15_4 = ~(a[15] & b[4]);
  assign f_s_dadda_rca16_and_14_5 = a[14] & b[5];
  assign f_s_dadda_rca16_fa102_xor0 = f_s_dadda_rca16_fa8_or0 ^ f_s_dadda_rca16_nand_15_4;
  assign f_s_dadda_rca16_fa102_and0 = f_s_dadda_rca16_fa8_or0 & f_s_dadda_rca16_nand_15_4;
  assign f_s_dadda_rca16_fa102_xor1 = f_s_dadda_rca16_fa102_xor0 ^ f_s_dadda_rca16_and_14_5;
  assign f_s_dadda_rca16_fa102_and1 = f_s_dadda_rca16_fa102_xor0 & f_s_dadda_rca16_and_14_5;
  assign f_s_dadda_rca16_fa102_or0 = f_s_dadda_rca16_fa102_and0 | f_s_dadda_rca16_fa102_and1;
  assign f_s_dadda_rca16_and_13_6 = a[13] & b[6];
  assign f_s_dadda_rca16_and_12_7 = a[12] & b[7];
  assign f_s_dadda_rca16_and_11_8 = a[11] & b[8];
  assign f_s_dadda_rca16_fa103_xor0 = f_s_dadda_rca16_and_13_6 ^ f_s_dadda_rca16_and_12_7;
  assign f_s_dadda_rca16_fa103_and0 = f_s_dadda_rca16_and_13_6 & f_s_dadda_rca16_and_12_7;
  assign f_s_dadda_rca16_fa103_xor1 = f_s_dadda_rca16_fa103_xor0 ^ f_s_dadda_rca16_and_11_8;
  assign f_s_dadda_rca16_fa103_and1 = f_s_dadda_rca16_fa103_xor0 & f_s_dadda_rca16_and_11_8;
  assign f_s_dadda_rca16_fa103_or0 = f_s_dadda_rca16_fa103_and0 | f_s_dadda_rca16_fa103_and1;
  assign f_s_dadda_rca16_and_10_9 = a[10] & b[9];
  assign f_s_dadda_rca16_and_9_10 = a[9] & b[10];
  assign f_s_dadda_rca16_and_8_11 = a[8] & b[11];
  assign f_s_dadda_rca16_fa104_xor0 = f_s_dadda_rca16_and_10_9 ^ f_s_dadda_rca16_and_9_10;
  assign f_s_dadda_rca16_fa104_and0 = f_s_dadda_rca16_and_10_9 & f_s_dadda_rca16_and_9_10;
  assign f_s_dadda_rca16_fa104_xor1 = f_s_dadda_rca16_fa104_xor0 ^ f_s_dadda_rca16_and_8_11;
  assign f_s_dadda_rca16_fa104_and1 = f_s_dadda_rca16_fa104_xor0 & f_s_dadda_rca16_and_8_11;
  assign f_s_dadda_rca16_fa104_or0 = f_s_dadda_rca16_fa104_and0 | f_s_dadda_rca16_fa104_and1;
  assign f_s_dadda_rca16_and_7_12 = a[7] & b[12];
  assign f_s_dadda_rca16_and_6_13 = a[6] & b[13];
  assign f_s_dadda_rca16_and_5_14 = a[5] & b[14];
  assign f_s_dadda_rca16_fa105_xor0 = f_s_dadda_rca16_and_7_12 ^ f_s_dadda_rca16_and_6_13;
  assign f_s_dadda_rca16_fa105_and0 = f_s_dadda_rca16_and_7_12 & f_s_dadda_rca16_and_6_13;
  assign f_s_dadda_rca16_fa105_xor1 = f_s_dadda_rca16_fa105_xor0 ^ f_s_dadda_rca16_and_5_14;
  assign f_s_dadda_rca16_fa105_and1 = f_s_dadda_rca16_fa105_xor0 & f_s_dadda_rca16_and_5_14;
  assign f_s_dadda_rca16_fa105_or0 = f_s_dadda_rca16_fa105_and0 | f_s_dadda_rca16_fa105_and1;
  assign f_s_dadda_rca16_nand_4_15 = ~(a[4] & b[15]);
  assign f_s_dadda_rca16_fa106_xor0 = f_s_dadda_rca16_nand_4_15 ^ f_s_dadda_rca16_fa99_xor1;
  assign f_s_dadda_rca16_fa106_and0 = f_s_dadda_rca16_nand_4_15 & f_s_dadda_rca16_fa99_xor1;
  assign f_s_dadda_rca16_fa106_xor1 = f_s_dadda_rca16_fa106_xor0 ^ f_s_dadda_rca16_fa100_xor1;
  assign f_s_dadda_rca16_fa106_and1 = f_s_dadda_rca16_fa106_xor0 & f_s_dadda_rca16_fa100_xor1;
  assign f_s_dadda_rca16_fa106_or0 = f_s_dadda_rca16_fa106_and0 | f_s_dadda_rca16_fa106_and1;
  assign f_s_dadda_rca16_fa107_xor0 = f_s_dadda_rca16_fa101_xor1 ^ f_s_dadda_rca16_fa102_xor1;
  assign f_s_dadda_rca16_fa107_and0 = f_s_dadda_rca16_fa101_xor1 & f_s_dadda_rca16_fa102_xor1;
  assign f_s_dadda_rca16_fa107_xor1 = f_s_dadda_rca16_fa107_xor0 ^ f_s_dadda_rca16_fa103_xor1;
  assign f_s_dadda_rca16_fa107_and1 = f_s_dadda_rca16_fa107_xor0 & f_s_dadda_rca16_fa103_xor1;
  assign f_s_dadda_rca16_fa107_or0 = f_s_dadda_rca16_fa107_and0 | f_s_dadda_rca16_fa107_and1;
  assign f_s_dadda_rca16_fa108_xor0 = f_s_dadda_rca16_fa107_or0 ^ f_s_dadda_rca16_fa106_or0;
  assign f_s_dadda_rca16_fa108_and0 = f_s_dadda_rca16_fa107_or0 & f_s_dadda_rca16_fa106_or0;
  assign f_s_dadda_rca16_fa108_xor1 = f_s_dadda_rca16_fa108_xor0 ^ f_s_dadda_rca16_fa105_or0;
  assign f_s_dadda_rca16_fa108_and1 = f_s_dadda_rca16_fa108_xor0 & f_s_dadda_rca16_fa105_or0;
  assign f_s_dadda_rca16_fa108_or0 = f_s_dadda_rca16_fa108_and0 | f_s_dadda_rca16_fa108_and1;
  assign f_s_dadda_rca16_fa109_xor0 = f_s_dadda_rca16_fa104_or0 ^ f_s_dadda_rca16_fa103_or0;
  assign f_s_dadda_rca16_fa109_and0 = f_s_dadda_rca16_fa104_or0 & f_s_dadda_rca16_fa103_or0;
  assign f_s_dadda_rca16_fa109_xor1 = f_s_dadda_rca16_fa109_xor0 ^ f_s_dadda_rca16_fa102_or0;
  assign f_s_dadda_rca16_fa109_and1 = f_s_dadda_rca16_fa109_xor0 & f_s_dadda_rca16_fa102_or0;
  assign f_s_dadda_rca16_fa109_or0 = f_s_dadda_rca16_fa109_and0 | f_s_dadda_rca16_fa109_and1;
  assign f_s_dadda_rca16_fa110_xor0 = f_s_dadda_rca16_fa101_or0 ^ f_s_dadda_rca16_fa100_or0;
  assign f_s_dadda_rca16_fa110_and0 = f_s_dadda_rca16_fa101_or0 & f_s_dadda_rca16_fa100_or0;
  assign f_s_dadda_rca16_fa110_xor1 = f_s_dadda_rca16_fa110_xor0 ^ f_s_dadda_rca16_fa99_or0;
  assign f_s_dadda_rca16_fa110_and1 = f_s_dadda_rca16_fa110_xor0 & f_s_dadda_rca16_fa99_or0;
  assign f_s_dadda_rca16_fa110_or0 = f_s_dadda_rca16_fa110_and0 | f_s_dadda_rca16_fa110_and1;
  assign f_s_dadda_rca16_nand_15_5 = ~(a[15] & b[5]);
  assign f_s_dadda_rca16_and_14_6 = a[14] & b[6];
  assign f_s_dadda_rca16_and_13_7 = a[13] & b[7];
  assign f_s_dadda_rca16_fa111_xor0 = f_s_dadda_rca16_nand_15_5 ^ f_s_dadda_rca16_and_14_6;
  assign f_s_dadda_rca16_fa111_and0 = f_s_dadda_rca16_nand_15_5 & f_s_dadda_rca16_and_14_6;
  assign f_s_dadda_rca16_fa111_xor1 = f_s_dadda_rca16_fa111_xor0 ^ f_s_dadda_rca16_and_13_7;
  assign f_s_dadda_rca16_fa111_and1 = f_s_dadda_rca16_fa111_xor0 & f_s_dadda_rca16_and_13_7;
  assign f_s_dadda_rca16_fa111_or0 = f_s_dadda_rca16_fa111_and0 | f_s_dadda_rca16_fa111_and1;
  assign f_s_dadda_rca16_and_12_8 = a[12] & b[8];
  assign f_s_dadda_rca16_and_11_9 = a[11] & b[9];
  assign f_s_dadda_rca16_and_10_10 = a[10] & b[10];
  assign f_s_dadda_rca16_fa112_xor0 = f_s_dadda_rca16_and_12_8 ^ f_s_dadda_rca16_and_11_9;
  assign f_s_dadda_rca16_fa112_and0 = f_s_dadda_rca16_and_12_8 & f_s_dadda_rca16_and_11_9;
  assign f_s_dadda_rca16_fa112_xor1 = f_s_dadda_rca16_fa112_xor0 ^ f_s_dadda_rca16_and_10_10;
  assign f_s_dadda_rca16_fa112_and1 = f_s_dadda_rca16_fa112_xor0 & f_s_dadda_rca16_and_10_10;
  assign f_s_dadda_rca16_fa112_or0 = f_s_dadda_rca16_fa112_and0 | f_s_dadda_rca16_fa112_and1;
  assign f_s_dadda_rca16_and_9_11 = a[9] & b[11];
  assign f_s_dadda_rca16_and_8_12 = a[8] & b[12];
  assign f_s_dadda_rca16_and_7_13 = a[7] & b[13];
  assign f_s_dadda_rca16_fa113_xor0 = f_s_dadda_rca16_and_9_11 ^ f_s_dadda_rca16_and_8_12;
  assign f_s_dadda_rca16_fa113_and0 = f_s_dadda_rca16_and_9_11 & f_s_dadda_rca16_and_8_12;
  assign f_s_dadda_rca16_fa113_xor1 = f_s_dadda_rca16_fa113_xor0 ^ f_s_dadda_rca16_and_7_13;
  assign f_s_dadda_rca16_fa113_and1 = f_s_dadda_rca16_fa113_xor0 & f_s_dadda_rca16_and_7_13;
  assign f_s_dadda_rca16_fa113_or0 = f_s_dadda_rca16_fa113_and0 | f_s_dadda_rca16_fa113_and1;
  assign f_s_dadda_rca16_and_6_14 = a[6] & b[14];
  assign f_s_dadda_rca16_nand_5_15 = ~(a[5] & b[15]);
  assign f_s_dadda_rca16_fa114_xor0 = f_s_dadda_rca16_and_6_14 ^ f_s_dadda_rca16_nand_5_15;
  assign f_s_dadda_rca16_fa114_and0 = f_s_dadda_rca16_and_6_14 & f_s_dadda_rca16_nand_5_15;
  assign f_s_dadda_rca16_fa114_xor1 = f_s_dadda_rca16_fa114_xor0 ^ f_s_dadda_rca16_fa108_xor1;
  assign f_s_dadda_rca16_fa114_and1 = f_s_dadda_rca16_fa114_xor0 & f_s_dadda_rca16_fa108_xor1;
  assign f_s_dadda_rca16_fa114_or0 = f_s_dadda_rca16_fa114_and0 | f_s_dadda_rca16_fa114_and1;
  assign f_s_dadda_rca16_fa115_xor0 = f_s_dadda_rca16_fa109_xor1 ^ f_s_dadda_rca16_fa110_xor1;
  assign f_s_dadda_rca16_fa115_and0 = f_s_dadda_rca16_fa109_xor1 & f_s_dadda_rca16_fa110_xor1;
  assign f_s_dadda_rca16_fa115_xor1 = f_s_dadda_rca16_fa115_xor0 ^ f_s_dadda_rca16_fa111_xor1;
  assign f_s_dadda_rca16_fa115_and1 = f_s_dadda_rca16_fa115_xor0 & f_s_dadda_rca16_fa111_xor1;
  assign f_s_dadda_rca16_fa115_or0 = f_s_dadda_rca16_fa115_and0 | f_s_dadda_rca16_fa115_and1;
  assign f_s_dadda_rca16_fa116_xor0 = f_s_dadda_rca16_fa115_or0 ^ f_s_dadda_rca16_fa114_or0;
  assign f_s_dadda_rca16_fa116_and0 = f_s_dadda_rca16_fa115_or0 & f_s_dadda_rca16_fa114_or0;
  assign f_s_dadda_rca16_fa116_xor1 = f_s_dadda_rca16_fa116_xor0 ^ f_s_dadda_rca16_fa113_or0;
  assign f_s_dadda_rca16_fa116_and1 = f_s_dadda_rca16_fa116_xor0 & f_s_dadda_rca16_fa113_or0;
  assign f_s_dadda_rca16_fa116_or0 = f_s_dadda_rca16_fa116_and0 | f_s_dadda_rca16_fa116_and1;
  assign f_s_dadda_rca16_fa117_xor0 = f_s_dadda_rca16_fa112_or0 ^ f_s_dadda_rca16_fa111_or0;
  assign f_s_dadda_rca16_fa117_and0 = f_s_dadda_rca16_fa112_or0 & f_s_dadda_rca16_fa111_or0;
  assign f_s_dadda_rca16_fa117_xor1 = f_s_dadda_rca16_fa117_xor0 ^ f_s_dadda_rca16_fa110_or0;
  assign f_s_dadda_rca16_fa117_and1 = f_s_dadda_rca16_fa117_xor0 & f_s_dadda_rca16_fa110_or0;
  assign f_s_dadda_rca16_fa117_or0 = f_s_dadda_rca16_fa117_and0 | f_s_dadda_rca16_fa117_and1;
  assign f_s_dadda_rca16_nand_15_6 = ~(a[15] & b[6]);
  assign f_s_dadda_rca16_fa118_xor0 = f_s_dadda_rca16_fa109_or0 ^ f_s_dadda_rca16_fa108_or0;
  assign f_s_dadda_rca16_fa118_and0 = f_s_dadda_rca16_fa109_or0 & f_s_dadda_rca16_fa108_or0;
  assign f_s_dadda_rca16_fa118_xor1 = f_s_dadda_rca16_fa118_xor0 ^ f_s_dadda_rca16_nand_15_6;
  assign f_s_dadda_rca16_fa118_and1 = f_s_dadda_rca16_fa118_xor0 & f_s_dadda_rca16_nand_15_6;
  assign f_s_dadda_rca16_fa118_or0 = f_s_dadda_rca16_fa118_and0 | f_s_dadda_rca16_fa118_and1;
  assign f_s_dadda_rca16_and_14_7 = a[14] & b[7];
  assign f_s_dadda_rca16_and_13_8 = a[13] & b[8];
  assign f_s_dadda_rca16_and_12_9 = a[12] & b[9];
  assign f_s_dadda_rca16_fa119_xor0 = f_s_dadda_rca16_and_14_7 ^ f_s_dadda_rca16_and_13_8;
  assign f_s_dadda_rca16_fa119_and0 = f_s_dadda_rca16_and_14_7 & f_s_dadda_rca16_and_13_8;
  assign f_s_dadda_rca16_fa119_xor1 = f_s_dadda_rca16_fa119_xor0 ^ f_s_dadda_rca16_and_12_9;
  assign f_s_dadda_rca16_fa119_and1 = f_s_dadda_rca16_fa119_xor0 & f_s_dadda_rca16_and_12_9;
  assign f_s_dadda_rca16_fa119_or0 = f_s_dadda_rca16_fa119_and0 | f_s_dadda_rca16_fa119_and1;
  assign f_s_dadda_rca16_and_11_10 = a[11] & b[10];
  assign f_s_dadda_rca16_and_10_11 = a[10] & b[11];
  assign f_s_dadda_rca16_and_9_12 = a[9] & b[12];
  assign f_s_dadda_rca16_fa120_xor0 = f_s_dadda_rca16_and_11_10 ^ f_s_dadda_rca16_and_10_11;
  assign f_s_dadda_rca16_fa120_and0 = f_s_dadda_rca16_and_11_10 & f_s_dadda_rca16_and_10_11;
  assign f_s_dadda_rca16_fa120_xor1 = f_s_dadda_rca16_fa120_xor0 ^ f_s_dadda_rca16_and_9_12;
  assign f_s_dadda_rca16_fa120_and1 = f_s_dadda_rca16_fa120_xor0 & f_s_dadda_rca16_and_9_12;
  assign f_s_dadda_rca16_fa120_or0 = f_s_dadda_rca16_fa120_and0 | f_s_dadda_rca16_fa120_and1;
  assign f_s_dadda_rca16_and_8_13 = a[8] & b[13];
  assign f_s_dadda_rca16_and_7_14 = a[7] & b[14];
  assign f_s_dadda_rca16_nand_6_15 = ~(a[6] & b[15]);
  assign f_s_dadda_rca16_fa121_xor0 = f_s_dadda_rca16_and_8_13 ^ f_s_dadda_rca16_and_7_14;
  assign f_s_dadda_rca16_fa121_and0 = f_s_dadda_rca16_and_8_13 & f_s_dadda_rca16_and_7_14;
  assign f_s_dadda_rca16_fa121_xor1 = f_s_dadda_rca16_fa121_xor0 ^ f_s_dadda_rca16_nand_6_15;
  assign f_s_dadda_rca16_fa121_and1 = f_s_dadda_rca16_fa121_xor0 & f_s_dadda_rca16_nand_6_15;
  assign f_s_dadda_rca16_fa121_or0 = f_s_dadda_rca16_fa121_and0 | f_s_dadda_rca16_fa121_and1;
  assign f_s_dadda_rca16_fa122_xor0 = f_s_dadda_rca16_fa116_xor1 ^ f_s_dadda_rca16_fa117_xor1;
  assign f_s_dadda_rca16_fa122_and0 = f_s_dadda_rca16_fa116_xor1 & f_s_dadda_rca16_fa117_xor1;
  assign f_s_dadda_rca16_fa122_xor1 = f_s_dadda_rca16_fa122_xor0 ^ f_s_dadda_rca16_fa118_xor1;
  assign f_s_dadda_rca16_fa122_and1 = f_s_dadda_rca16_fa122_xor0 & f_s_dadda_rca16_fa118_xor1;
  assign f_s_dadda_rca16_fa122_or0 = f_s_dadda_rca16_fa122_and0 | f_s_dadda_rca16_fa122_and1;
  assign f_s_dadda_rca16_fa123_xor0 = f_s_dadda_rca16_fa122_or0 ^ f_s_dadda_rca16_fa121_or0;
  assign f_s_dadda_rca16_fa123_and0 = f_s_dadda_rca16_fa122_or0 & f_s_dadda_rca16_fa121_or0;
  assign f_s_dadda_rca16_fa123_xor1 = f_s_dadda_rca16_fa123_xor0 ^ f_s_dadda_rca16_fa120_or0;
  assign f_s_dadda_rca16_fa123_and1 = f_s_dadda_rca16_fa123_xor0 & f_s_dadda_rca16_fa120_or0;
  assign f_s_dadda_rca16_fa123_or0 = f_s_dadda_rca16_fa123_and0 | f_s_dadda_rca16_fa123_and1;
  assign f_s_dadda_rca16_fa124_xor0 = f_s_dadda_rca16_fa119_or0 ^ f_s_dadda_rca16_fa118_or0;
  assign f_s_dadda_rca16_fa124_and0 = f_s_dadda_rca16_fa119_or0 & f_s_dadda_rca16_fa118_or0;
  assign f_s_dadda_rca16_fa124_xor1 = f_s_dadda_rca16_fa124_xor0 ^ f_s_dadda_rca16_fa117_or0;
  assign f_s_dadda_rca16_fa124_and1 = f_s_dadda_rca16_fa124_xor0 & f_s_dadda_rca16_fa117_or0;
  assign f_s_dadda_rca16_fa124_or0 = f_s_dadda_rca16_fa124_and0 | f_s_dadda_rca16_fa124_and1;
  assign f_s_dadda_rca16_nand_15_7 = ~(a[15] & b[7]);
  assign f_s_dadda_rca16_and_14_8 = a[14] & b[8];
  assign f_s_dadda_rca16_fa125_xor0 = f_s_dadda_rca16_fa116_or0 ^ f_s_dadda_rca16_nand_15_7;
  assign f_s_dadda_rca16_fa125_and0 = f_s_dadda_rca16_fa116_or0 & f_s_dadda_rca16_nand_15_7;
  assign f_s_dadda_rca16_fa125_xor1 = f_s_dadda_rca16_fa125_xor0 ^ f_s_dadda_rca16_and_14_8;
  assign f_s_dadda_rca16_fa125_and1 = f_s_dadda_rca16_fa125_xor0 & f_s_dadda_rca16_and_14_8;
  assign f_s_dadda_rca16_fa125_or0 = f_s_dadda_rca16_fa125_and0 | f_s_dadda_rca16_fa125_and1;
  assign f_s_dadda_rca16_and_13_9 = a[13] & b[9];
  assign f_s_dadda_rca16_and_12_10 = a[12] & b[10];
  assign f_s_dadda_rca16_and_11_11 = a[11] & b[11];
  assign f_s_dadda_rca16_fa126_xor0 = f_s_dadda_rca16_and_13_9 ^ f_s_dadda_rca16_and_12_10;
  assign f_s_dadda_rca16_fa126_and0 = f_s_dadda_rca16_and_13_9 & f_s_dadda_rca16_and_12_10;
  assign f_s_dadda_rca16_fa126_xor1 = f_s_dadda_rca16_fa126_xor0 ^ f_s_dadda_rca16_and_11_11;
  assign f_s_dadda_rca16_fa126_and1 = f_s_dadda_rca16_fa126_xor0 & f_s_dadda_rca16_and_11_11;
  assign f_s_dadda_rca16_fa126_or0 = f_s_dadda_rca16_fa126_and0 | f_s_dadda_rca16_fa126_and1;
  assign f_s_dadda_rca16_and_10_12 = a[10] & b[12];
  assign f_s_dadda_rca16_and_9_13 = a[9] & b[13];
  assign f_s_dadda_rca16_and_8_14 = a[8] & b[14];
  assign f_s_dadda_rca16_fa127_xor0 = f_s_dadda_rca16_and_10_12 ^ f_s_dadda_rca16_and_9_13;
  assign f_s_dadda_rca16_fa127_and0 = f_s_dadda_rca16_and_10_12 & f_s_dadda_rca16_and_9_13;
  assign f_s_dadda_rca16_fa127_xor1 = f_s_dadda_rca16_fa127_xor0 ^ f_s_dadda_rca16_and_8_14;
  assign f_s_dadda_rca16_fa127_and1 = f_s_dadda_rca16_fa127_xor0 & f_s_dadda_rca16_and_8_14;
  assign f_s_dadda_rca16_fa127_or0 = f_s_dadda_rca16_fa127_and0 | f_s_dadda_rca16_fa127_and1;
  assign f_s_dadda_rca16_nand_7_15 = ~(a[7] & b[15]);
  assign f_s_dadda_rca16_fa128_xor0 = f_s_dadda_rca16_nand_7_15 ^ f_s_dadda_rca16_fa123_xor1;
  assign f_s_dadda_rca16_fa128_and0 = f_s_dadda_rca16_nand_7_15 & f_s_dadda_rca16_fa123_xor1;
  assign f_s_dadda_rca16_fa128_xor1 = f_s_dadda_rca16_fa128_xor0 ^ f_s_dadda_rca16_fa124_xor1;
  assign f_s_dadda_rca16_fa128_and1 = f_s_dadda_rca16_fa128_xor0 & f_s_dadda_rca16_fa124_xor1;
  assign f_s_dadda_rca16_fa128_or0 = f_s_dadda_rca16_fa128_and0 | f_s_dadda_rca16_fa128_and1;
  assign f_s_dadda_rca16_fa129_xor0 = f_s_dadda_rca16_fa128_or0 ^ f_s_dadda_rca16_fa127_or0;
  assign f_s_dadda_rca16_fa129_and0 = f_s_dadda_rca16_fa128_or0 & f_s_dadda_rca16_fa127_or0;
  assign f_s_dadda_rca16_fa129_xor1 = f_s_dadda_rca16_fa129_xor0 ^ f_s_dadda_rca16_fa126_or0;
  assign f_s_dadda_rca16_fa129_and1 = f_s_dadda_rca16_fa129_xor0 & f_s_dadda_rca16_fa126_or0;
  assign f_s_dadda_rca16_fa129_or0 = f_s_dadda_rca16_fa129_and0 | f_s_dadda_rca16_fa129_and1;
  assign f_s_dadda_rca16_fa130_xor0 = f_s_dadda_rca16_fa125_or0 ^ f_s_dadda_rca16_fa124_or0;
  assign f_s_dadda_rca16_fa130_and0 = f_s_dadda_rca16_fa125_or0 & f_s_dadda_rca16_fa124_or0;
  assign f_s_dadda_rca16_fa130_xor1 = f_s_dadda_rca16_fa130_xor0 ^ f_s_dadda_rca16_fa123_or0;
  assign f_s_dadda_rca16_fa130_and1 = f_s_dadda_rca16_fa130_xor0 & f_s_dadda_rca16_fa123_or0;
  assign f_s_dadda_rca16_fa130_or0 = f_s_dadda_rca16_fa130_and0 | f_s_dadda_rca16_fa130_and1;
  assign f_s_dadda_rca16_nand_15_8 = ~(a[15] & b[8]);
  assign f_s_dadda_rca16_and_14_9 = a[14] & b[9];
  assign f_s_dadda_rca16_and_13_10 = a[13] & b[10];
  assign f_s_dadda_rca16_fa131_xor0 = f_s_dadda_rca16_nand_15_8 ^ f_s_dadda_rca16_and_14_9;
  assign f_s_dadda_rca16_fa131_and0 = f_s_dadda_rca16_nand_15_8 & f_s_dadda_rca16_and_14_9;
  assign f_s_dadda_rca16_fa131_xor1 = f_s_dadda_rca16_fa131_xor0 ^ f_s_dadda_rca16_and_13_10;
  assign f_s_dadda_rca16_fa131_and1 = f_s_dadda_rca16_fa131_xor0 & f_s_dadda_rca16_and_13_10;
  assign f_s_dadda_rca16_fa131_or0 = f_s_dadda_rca16_fa131_and0 | f_s_dadda_rca16_fa131_and1;
  assign f_s_dadda_rca16_and_12_11 = a[12] & b[11];
  assign f_s_dadda_rca16_and_11_12 = a[11] & b[12];
  assign f_s_dadda_rca16_and_10_13 = a[10] & b[13];
  assign f_s_dadda_rca16_fa132_xor0 = f_s_dadda_rca16_and_12_11 ^ f_s_dadda_rca16_and_11_12;
  assign f_s_dadda_rca16_fa132_and0 = f_s_dadda_rca16_and_12_11 & f_s_dadda_rca16_and_11_12;
  assign f_s_dadda_rca16_fa132_xor1 = f_s_dadda_rca16_fa132_xor0 ^ f_s_dadda_rca16_and_10_13;
  assign f_s_dadda_rca16_fa132_and1 = f_s_dadda_rca16_fa132_xor0 & f_s_dadda_rca16_and_10_13;
  assign f_s_dadda_rca16_fa132_or0 = f_s_dadda_rca16_fa132_and0 | f_s_dadda_rca16_fa132_and1;
  assign f_s_dadda_rca16_and_9_14 = a[9] & b[14];
  assign f_s_dadda_rca16_nand_8_15 = ~(a[8] & b[15]);
  assign f_s_dadda_rca16_fa133_xor0 = f_s_dadda_rca16_and_9_14 ^ f_s_dadda_rca16_nand_8_15;
  assign f_s_dadda_rca16_fa133_and0 = f_s_dadda_rca16_and_9_14 & f_s_dadda_rca16_nand_8_15;
  assign f_s_dadda_rca16_fa133_xor1 = f_s_dadda_rca16_fa133_xor0 ^ f_s_dadda_rca16_fa129_xor1;
  assign f_s_dadda_rca16_fa133_and1 = f_s_dadda_rca16_fa133_xor0 & f_s_dadda_rca16_fa129_xor1;
  assign f_s_dadda_rca16_fa133_or0 = f_s_dadda_rca16_fa133_and0 | f_s_dadda_rca16_fa133_and1;
  assign f_s_dadda_rca16_fa134_xor0 = f_s_dadda_rca16_fa133_or0 ^ f_s_dadda_rca16_fa132_or0;
  assign f_s_dadda_rca16_fa134_and0 = f_s_dadda_rca16_fa133_or0 & f_s_dadda_rca16_fa132_or0;
  assign f_s_dadda_rca16_fa134_xor1 = f_s_dadda_rca16_fa134_xor0 ^ f_s_dadda_rca16_fa131_or0;
  assign f_s_dadda_rca16_fa134_and1 = f_s_dadda_rca16_fa134_xor0 & f_s_dadda_rca16_fa131_or0;
  assign f_s_dadda_rca16_fa134_or0 = f_s_dadda_rca16_fa134_and0 | f_s_dadda_rca16_fa134_and1;
  assign f_s_dadda_rca16_nand_15_9 = ~(a[15] & b[9]);
  assign f_s_dadda_rca16_fa135_xor0 = f_s_dadda_rca16_fa130_or0 ^ f_s_dadda_rca16_fa129_or0;
  assign f_s_dadda_rca16_fa135_and0 = f_s_dadda_rca16_fa130_or0 & f_s_dadda_rca16_fa129_or0;
  assign f_s_dadda_rca16_fa135_xor1 = f_s_dadda_rca16_fa135_xor0 ^ f_s_dadda_rca16_nand_15_9;
  assign f_s_dadda_rca16_fa135_and1 = f_s_dadda_rca16_fa135_xor0 & f_s_dadda_rca16_nand_15_9;
  assign f_s_dadda_rca16_fa135_or0 = f_s_dadda_rca16_fa135_and0 | f_s_dadda_rca16_fa135_and1;
  assign f_s_dadda_rca16_and_14_10 = a[14] & b[10];
  assign f_s_dadda_rca16_and_13_11 = a[13] & b[11];
  assign f_s_dadda_rca16_and_12_12 = a[12] & b[12];
  assign f_s_dadda_rca16_fa136_xor0 = f_s_dadda_rca16_and_14_10 ^ f_s_dadda_rca16_and_13_11;
  assign f_s_dadda_rca16_fa136_and0 = f_s_dadda_rca16_and_14_10 & f_s_dadda_rca16_and_13_11;
  assign f_s_dadda_rca16_fa136_xor1 = f_s_dadda_rca16_fa136_xor0 ^ f_s_dadda_rca16_and_12_12;
  assign f_s_dadda_rca16_fa136_and1 = f_s_dadda_rca16_fa136_xor0 & f_s_dadda_rca16_and_12_12;
  assign f_s_dadda_rca16_fa136_or0 = f_s_dadda_rca16_fa136_and0 | f_s_dadda_rca16_fa136_and1;
  assign f_s_dadda_rca16_and_11_13 = a[11] & b[13];
  assign f_s_dadda_rca16_and_10_14 = a[10] & b[14];
  assign f_s_dadda_rca16_nand_9_15 = ~(a[9] & b[15]);
  assign f_s_dadda_rca16_fa137_xor0 = f_s_dadda_rca16_and_11_13 ^ f_s_dadda_rca16_and_10_14;
  assign f_s_dadda_rca16_fa137_and0 = f_s_dadda_rca16_and_11_13 & f_s_dadda_rca16_and_10_14;
  assign f_s_dadda_rca16_fa137_xor1 = f_s_dadda_rca16_fa137_xor0 ^ f_s_dadda_rca16_nand_9_15;
  assign f_s_dadda_rca16_fa137_and1 = f_s_dadda_rca16_fa137_xor0 & f_s_dadda_rca16_nand_9_15;
  assign f_s_dadda_rca16_fa137_or0 = f_s_dadda_rca16_fa137_and0 | f_s_dadda_rca16_fa137_and1;
  assign f_s_dadda_rca16_fa138_xor0 = f_s_dadda_rca16_fa137_or0 ^ f_s_dadda_rca16_fa136_or0;
  assign f_s_dadda_rca16_fa138_and0 = f_s_dadda_rca16_fa137_or0 & f_s_dadda_rca16_fa136_or0;
  assign f_s_dadda_rca16_fa138_xor1 = f_s_dadda_rca16_fa138_xor0 ^ f_s_dadda_rca16_fa135_or0;
  assign f_s_dadda_rca16_fa138_and1 = f_s_dadda_rca16_fa138_xor0 & f_s_dadda_rca16_fa135_or0;
  assign f_s_dadda_rca16_fa138_or0 = f_s_dadda_rca16_fa138_and0 | f_s_dadda_rca16_fa138_and1;
  assign f_s_dadda_rca16_nand_15_10 = ~(a[15] & b[10]);
  assign f_s_dadda_rca16_and_14_11 = a[14] & b[11];
  assign f_s_dadda_rca16_fa139_xor0 = f_s_dadda_rca16_fa134_or0 ^ f_s_dadda_rca16_nand_15_10;
  assign f_s_dadda_rca16_fa139_and0 = f_s_dadda_rca16_fa134_or0 & f_s_dadda_rca16_nand_15_10;
  assign f_s_dadda_rca16_fa139_xor1 = f_s_dadda_rca16_fa139_xor0 ^ f_s_dadda_rca16_and_14_11;
  assign f_s_dadda_rca16_fa139_and1 = f_s_dadda_rca16_fa139_xor0 & f_s_dadda_rca16_and_14_11;
  assign f_s_dadda_rca16_fa139_or0 = f_s_dadda_rca16_fa139_and0 | f_s_dadda_rca16_fa139_and1;
  assign f_s_dadda_rca16_and_13_12 = a[13] & b[12];
  assign f_s_dadda_rca16_and_12_13 = a[12] & b[13];
  assign f_s_dadda_rca16_and_11_14 = a[11] & b[14];
  assign f_s_dadda_rca16_fa140_xor0 = f_s_dadda_rca16_and_13_12 ^ f_s_dadda_rca16_and_12_13;
  assign f_s_dadda_rca16_fa140_and0 = f_s_dadda_rca16_and_13_12 & f_s_dadda_rca16_and_12_13;
  assign f_s_dadda_rca16_fa140_xor1 = f_s_dadda_rca16_fa140_xor0 ^ f_s_dadda_rca16_and_11_14;
  assign f_s_dadda_rca16_fa140_and1 = f_s_dadda_rca16_fa140_xor0 & f_s_dadda_rca16_and_11_14;
  assign f_s_dadda_rca16_fa140_or0 = f_s_dadda_rca16_fa140_and0 | f_s_dadda_rca16_fa140_and1;
  assign f_s_dadda_rca16_fa141_xor0 = f_s_dadda_rca16_fa140_or0 ^ f_s_dadda_rca16_fa139_or0;
  assign f_s_dadda_rca16_fa141_and0 = f_s_dadda_rca16_fa140_or0 & f_s_dadda_rca16_fa139_or0;
  assign f_s_dadda_rca16_fa141_xor1 = f_s_dadda_rca16_fa141_xor0 ^ f_s_dadda_rca16_fa138_or0;
  assign f_s_dadda_rca16_fa141_and1 = f_s_dadda_rca16_fa141_xor0 & f_s_dadda_rca16_fa138_or0;
  assign f_s_dadda_rca16_fa141_or0 = f_s_dadda_rca16_fa141_and0 | f_s_dadda_rca16_fa141_and1;
  assign f_s_dadda_rca16_nand_15_11 = ~(a[15] & b[11]);
  assign f_s_dadda_rca16_and_14_12 = a[14] & b[12];
  assign f_s_dadda_rca16_and_13_13 = a[13] & b[13];
  assign f_s_dadda_rca16_fa142_xor0 = f_s_dadda_rca16_nand_15_11 ^ f_s_dadda_rca16_and_14_12;
  assign f_s_dadda_rca16_fa142_and0 = f_s_dadda_rca16_nand_15_11 & f_s_dadda_rca16_and_14_12;
  assign f_s_dadda_rca16_fa142_xor1 = f_s_dadda_rca16_fa142_xor0 ^ f_s_dadda_rca16_and_13_13;
  assign f_s_dadda_rca16_fa142_and1 = f_s_dadda_rca16_fa142_xor0 & f_s_dadda_rca16_and_13_13;
  assign f_s_dadda_rca16_fa142_or0 = f_s_dadda_rca16_fa142_and0 | f_s_dadda_rca16_fa142_and1;
  assign f_s_dadda_rca16_nand_15_12 = ~(a[15] & b[12]);
  assign f_s_dadda_rca16_fa143_xor0 = f_s_dadda_rca16_fa142_or0 ^ f_s_dadda_rca16_fa141_or0;
  assign f_s_dadda_rca16_fa143_and0 = f_s_dadda_rca16_fa142_or0 & f_s_dadda_rca16_fa141_or0;
  assign f_s_dadda_rca16_fa143_xor1 = f_s_dadda_rca16_fa143_xor0 ^ f_s_dadda_rca16_nand_15_12;
  assign f_s_dadda_rca16_fa143_and1 = f_s_dadda_rca16_fa143_xor0 & f_s_dadda_rca16_nand_15_12;
  assign f_s_dadda_rca16_fa143_or0 = f_s_dadda_rca16_fa143_and0 | f_s_dadda_rca16_fa143_and1;
  assign f_s_dadda_rca16_and_3_0 = a[3] & b[0];
  assign f_s_dadda_rca16_and_2_1 = a[2] & b[1];
  assign f_s_dadda_rca16_ha12_xor0 = f_s_dadda_rca16_and_3_0 ^ f_s_dadda_rca16_and_2_1;
  assign f_s_dadda_rca16_ha12_and0 = f_s_dadda_rca16_and_3_0 & f_s_dadda_rca16_and_2_1;
  assign f_s_dadda_rca16_and_2_2 = a[2] & b[2];
  assign f_s_dadda_rca16_and_1_3 = a[1] & b[3];
  assign f_s_dadda_rca16_fa144_xor0 = f_s_dadda_rca16_ha12_and0 ^ f_s_dadda_rca16_and_2_2;
  assign f_s_dadda_rca16_fa144_and0 = f_s_dadda_rca16_ha12_and0 & f_s_dadda_rca16_and_2_2;
  assign f_s_dadda_rca16_fa144_xor1 = f_s_dadda_rca16_fa144_xor0 ^ f_s_dadda_rca16_and_1_3;
  assign f_s_dadda_rca16_fa144_and1 = f_s_dadda_rca16_fa144_xor0 & f_s_dadda_rca16_and_1_3;
  assign f_s_dadda_rca16_fa144_or0 = f_s_dadda_rca16_fa144_and0 | f_s_dadda_rca16_fa144_and1;
  assign f_s_dadda_rca16_and_1_4 = a[1] & b[4];
  assign f_s_dadda_rca16_and_0_5 = a[0] & b[5];
  assign f_s_dadda_rca16_fa145_xor0 = f_s_dadda_rca16_fa144_or0 ^ f_s_dadda_rca16_and_1_4;
  assign f_s_dadda_rca16_fa145_and0 = f_s_dadda_rca16_fa144_or0 & f_s_dadda_rca16_and_1_4;
  assign f_s_dadda_rca16_fa145_xor1 = f_s_dadda_rca16_fa145_xor0 ^ f_s_dadda_rca16_and_0_5;
  assign f_s_dadda_rca16_fa145_and1 = f_s_dadda_rca16_fa145_xor0 & f_s_dadda_rca16_and_0_5;
  assign f_s_dadda_rca16_fa145_or0 = f_s_dadda_rca16_fa145_and0 | f_s_dadda_rca16_fa145_and1;
  assign f_s_dadda_rca16_and_0_6 = a[0] & b[6];
  assign f_s_dadda_rca16_fa146_xor0 = f_s_dadda_rca16_fa145_or0 ^ f_s_dadda_rca16_and_0_6;
  assign f_s_dadda_rca16_fa146_and0 = f_s_dadda_rca16_fa145_or0 & f_s_dadda_rca16_and_0_6;
  assign f_s_dadda_rca16_fa146_xor1 = f_s_dadda_rca16_fa146_xor0 ^ f_s_dadda_rca16_fa10_xor1;
  assign f_s_dadda_rca16_fa146_and1 = f_s_dadda_rca16_fa146_xor0 & f_s_dadda_rca16_fa10_xor1;
  assign f_s_dadda_rca16_fa146_or0 = f_s_dadda_rca16_fa146_and0 | f_s_dadda_rca16_fa146_and1;
  assign f_s_dadda_rca16_fa147_xor0 = f_s_dadda_rca16_fa146_or0 ^ f_s_dadda_rca16_fa12_xor1;
  assign f_s_dadda_rca16_fa147_and0 = f_s_dadda_rca16_fa146_or0 & f_s_dadda_rca16_fa12_xor1;
  assign f_s_dadda_rca16_fa147_xor1 = f_s_dadda_rca16_fa147_xor0 ^ f_s_dadda_rca16_fa13_xor1;
  assign f_s_dadda_rca16_fa147_and1 = f_s_dadda_rca16_fa147_xor0 & f_s_dadda_rca16_fa13_xor1;
  assign f_s_dadda_rca16_fa147_or0 = f_s_dadda_rca16_fa147_and0 | f_s_dadda_rca16_fa147_and1;
  assign f_s_dadda_rca16_fa148_xor0 = f_s_dadda_rca16_fa147_or0 ^ f_s_dadda_rca16_fa16_xor1;
  assign f_s_dadda_rca16_fa148_and0 = f_s_dadda_rca16_fa147_or0 & f_s_dadda_rca16_fa16_xor1;
  assign f_s_dadda_rca16_fa148_xor1 = f_s_dadda_rca16_fa148_xor0 ^ f_s_dadda_rca16_fa17_xor1;
  assign f_s_dadda_rca16_fa148_and1 = f_s_dadda_rca16_fa148_xor0 & f_s_dadda_rca16_fa17_xor1;
  assign f_s_dadda_rca16_fa148_or0 = f_s_dadda_rca16_fa148_and0 | f_s_dadda_rca16_fa148_and1;
  assign f_s_dadda_rca16_fa149_xor0 = f_s_dadda_rca16_fa148_or0 ^ f_s_dadda_rca16_fa21_xor1;
  assign f_s_dadda_rca16_fa149_and0 = f_s_dadda_rca16_fa148_or0 & f_s_dadda_rca16_fa21_xor1;
  assign f_s_dadda_rca16_fa149_xor1 = f_s_dadda_rca16_fa149_xor0 ^ f_s_dadda_rca16_fa22_xor1;
  assign f_s_dadda_rca16_fa149_and1 = f_s_dadda_rca16_fa149_xor0 & f_s_dadda_rca16_fa22_xor1;
  assign f_s_dadda_rca16_fa149_or0 = f_s_dadda_rca16_fa149_and0 | f_s_dadda_rca16_fa149_and1;
  assign f_s_dadda_rca16_fa150_xor0 = f_s_dadda_rca16_fa149_or0 ^ f_s_dadda_rca16_fa27_xor1;
  assign f_s_dadda_rca16_fa150_and0 = f_s_dadda_rca16_fa149_or0 & f_s_dadda_rca16_fa27_xor1;
  assign f_s_dadda_rca16_fa150_xor1 = f_s_dadda_rca16_fa150_xor0 ^ f_s_dadda_rca16_fa28_xor1;
  assign f_s_dadda_rca16_fa150_and1 = f_s_dadda_rca16_fa150_xor0 & f_s_dadda_rca16_fa28_xor1;
  assign f_s_dadda_rca16_fa150_or0 = f_s_dadda_rca16_fa150_and0 | f_s_dadda_rca16_fa150_and1;
  assign f_s_dadda_rca16_fa151_xor0 = f_s_dadda_rca16_fa150_or0 ^ f_s_dadda_rca16_fa34_xor1;
  assign f_s_dadda_rca16_fa151_and0 = f_s_dadda_rca16_fa150_or0 & f_s_dadda_rca16_fa34_xor1;
  assign f_s_dadda_rca16_fa151_xor1 = f_s_dadda_rca16_fa151_xor0 ^ f_s_dadda_rca16_fa35_xor1;
  assign f_s_dadda_rca16_fa151_and1 = f_s_dadda_rca16_fa151_xor0 & f_s_dadda_rca16_fa35_xor1;
  assign f_s_dadda_rca16_fa151_or0 = f_s_dadda_rca16_fa151_and0 | f_s_dadda_rca16_fa151_and1;
  assign f_s_dadda_rca16_fa152_xor0 = f_s_dadda_rca16_fa151_or0 ^ f_s_dadda_rca16_fa42_xor1;
  assign f_s_dadda_rca16_fa152_and0 = f_s_dadda_rca16_fa151_or0 & f_s_dadda_rca16_fa42_xor1;
  assign f_s_dadda_rca16_fa152_xor1 = f_s_dadda_rca16_fa152_xor0 ^ f_s_dadda_rca16_fa43_xor1;
  assign f_s_dadda_rca16_fa152_and1 = f_s_dadda_rca16_fa152_xor0 & f_s_dadda_rca16_fa43_xor1;
  assign f_s_dadda_rca16_fa152_or0 = f_s_dadda_rca16_fa152_and0 | f_s_dadda_rca16_fa152_and1;
  assign f_s_dadda_rca16_fa153_xor0 = f_s_dadda_rca16_fa152_or0 ^ f_s_dadda_rca16_fa50_xor1;
  assign f_s_dadda_rca16_fa153_and0 = f_s_dadda_rca16_fa152_or0 & f_s_dadda_rca16_fa50_xor1;
  assign f_s_dadda_rca16_fa153_xor1 = f_s_dadda_rca16_fa153_xor0 ^ f_s_dadda_rca16_fa51_xor1;
  assign f_s_dadda_rca16_fa153_and1 = f_s_dadda_rca16_fa153_xor0 & f_s_dadda_rca16_fa51_xor1;
  assign f_s_dadda_rca16_fa153_or0 = f_s_dadda_rca16_fa153_and0 | f_s_dadda_rca16_fa153_and1;
  assign f_s_dadda_rca16_fa154_xor0 = f_s_dadda_rca16_fa153_or0 ^ f_s_dadda_rca16_fa59_xor1;
  assign f_s_dadda_rca16_fa154_and0 = f_s_dadda_rca16_fa153_or0 & f_s_dadda_rca16_fa59_xor1;
  assign f_s_dadda_rca16_fa154_xor1 = f_s_dadda_rca16_fa154_xor0 ^ f_s_dadda_rca16_fa60_xor1;
  assign f_s_dadda_rca16_fa154_and1 = f_s_dadda_rca16_fa154_xor0 & f_s_dadda_rca16_fa60_xor1;
  assign f_s_dadda_rca16_fa154_or0 = f_s_dadda_rca16_fa154_and0 | f_s_dadda_rca16_fa154_and1;
  assign f_s_dadda_rca16_fa155_xor0 = f_s_dadda_rca16_fa154_or0 ^ f_s_dadda_rca16_fa68_xor1;
  assign f_s_dadda_rca16_fa155_and0 = f_s_dadda_rca16_fa154_or0 & f_s_dadda_rca16_fa68_xor1;
  assign f_s_dadda_rca16_fa155_xor1 = f_s_dadda_rca16_fa155_xor0 ^ f_s_dadda_rca16_fa69_xor1;
  assign f_s_dadda_rca16_fa155_and1 = f_s_dadda_rca16_fa155_xor0 & f_s_dadda_rca16_fa69_xor1;
  assign f_s_dadda_rca16_fa155_or0 = f_s_dadda_rca16_fa155_and0 | f_s_dadda_rca16_fa155_and1;
  assign f_s_dadda_rca16_fa156_xor0 = f_s_dadda_rca16_fa155_or0 ^ f_s_dadda_rca16_fa77_xor1;
  assign f_s_dadda_rca16_fa156_and0 = f_s_dadda_rca16_fa155_or0 & f_s_dadda_rca16_fa77_xor1;
  assign f_s_dadda_rca16_fa156_xor1 = f_s_dadda_rca16_fa156_xor0 ^ f_s_dadda_rca16_fa78_xor1;
  assign f_s_dadda_rca16_fa156_and1 = f_s_dadda_rca16_fa156_xor0 & f_s_dadda_rca16_fa78_xor1;
  assign f_s_dadda_rca16_fa156_or0 = f_s_dadda_rca16_fa156_and0 | f_s_dadda_rca16_fa156_and1;
  assign f_s_dadda_rca16_fa157_xor0 = f_s_dadda_rca16_fa156_or0 ^ f_s_dadda_rca16_fa86_xor1;
  assign f_s_dadda_rca16_fa157_and0 = f_s_dadda_rca16_fa156_or0 & f_s_dadda_rca16_fa86_xor1;
  assign f_s_dadda_rca16_fa157_xor1 = f_s_dadda_rca16_fa157_xor0 ^ f_s_dadda_rca16_fa87_xor1;
  assign f_s_dadda_rca16_fa157_and1 = f_s_dadda_rca16_fa157_xor0 & f_s_dadda_rca16_fa87_xor1;
  assign f_s_dadda_rca16_fa157_or0 = f_s_dadda_rca16_fa157_and0 | f_s_dadda_rca16_fa157_and1;
  assign f_s_dadda_rca16_fa158_xor0 = f_s_dadda_rca16_fa157_or0 ^ f_s_dadda_rca16_fa95_xor1;
  assign f_s_dadda_rca16_fa158_and0 = f_s_dadda_rca16_fa157_or0 & f_s_dadda_rca16_fa95_xor1;
  assign f_s_dadda_rca16_fa158_xor1 = f_s_dadda_rca16_fa158_xor0 ^ f_s_dadda_rca16_fa96_xor1;
  assign f_s_dadda_rca16_fa158_and1 = f_s_dadda_rca16_fa158_xor0 & f_s_dadda_rca16_fa96_xor1;
  assign f_s_dadda_rca16_fa158_or0 = f_s_dadda_rca16_fa158_and0 | f_s_dadda_rca16_fa158_and1;
  assign f_s_dadda_rca16_fa159_xor0 = f_s_dadda_rca16_fa158_or0 ^ f_s_dadda_rca16_fa104_xor1;
  assign f_s_dadda_rca16_fa159_and0 = f_s_dadda_rca16_fa158_or0 & f_s_dadda_rca16_fa104_xor1;
  assign f_s_dadda_rca16_fa159_xor1 = f_s_dadda_rca16_fa159_xor0 ^ f_s_dadda_rca16_fa105_xor1;
  assign f_s_dadda_rca16_fa159_and1 = f_s_dadda_rca16_fa159_xor0 & f_s_dadda_rca16_fa105_xor1;
  assign f_s_dadda_rca16_fa159_or0 = f_s_dadda_rca16_fa159_and0 | f_s_dadda_rca16_fa159_and1;
  assign f_s_dadda_rca16_fa160_xor0 = f_s_dadda_rca16_fa159_or0 ^ f_s_dadda_rca16_fa112_xor1;
  assign f_s_dadda_rca16_fa160_and0 = f_s_dadda_rca16_fa159_or0 & f_s_dadda_rca16_fa112_xor1;
  assign f_s_dadda_rca16_fa160_xor1 = f_s_dadda_rca16_fa160_xor0 ^ f_s_dadda_rca16_fa113_xor1;
  assign f_s_dadda_rca16_fa160_and1 = f_s_dadda_rca16_fa160_xor0 & f_s_dadda_rca16_fa113_xor1;
  assign f_s_dadda_rca16_fa160_or0 = f_s_dadda_rca16_fa160_and0 | f_s_dadda_rca16_fa160_and1;
  assign f_s_dadda_rca16_fa161_xor0 = f_s_dadda_rca16_fa160_or0 ^ f_s_dadda_rca16_fa119_xor1;
  assign f_s_dadda_rca16_fa161_and0 = f_s_dadda_rca16_fa160_or0 & f_s_dadda_rca16_fa119_xor1;
  assign f_s_dadda_rca16_fa161_xor1 = f_s_dadda_rca16_fa161_xor0 ^ f_s_dadda_rca16_fa120_xor1;
  assign f_s_dadda_rca16_fa161_and1 = f_s_dadda_rca16_fa161_xor0 & f_s_dadda_rca16_fa120_xor1;
  assign f_s_dadda_rca16_fa161_or0 = f_s_dadda_rca16_fa161_and0 | f_s_dadda_rca16_fa161_and1;
  assign f_s_dadda_rca16_fa162_xor0 = f_s_dadda_rca16_fa161_or0 ^ f_s_dadda_rca16_fa125_xor1;
  assign f_s_dadda_rca16_fa162_and0 = f_s_dadda_rca16_fa161_or0 & f_s_dadda_rca16_fa125_xor1;
  assign f_s_dadda_rca16_fa162_xor1 = f_s_dadda_rca16_fa162_xor0 ^ f_s_dadda_rca16_fa126_xor1;
  assign f_s_dadda_rca16_fa162_and1 = f_s_dadda_rca16_fa162_xor0 & f_s_dadda_rca16_fa126_xor1;
  assign f_s_dadda_rca16_fa162_or0 = f_s_dadda_rca16_fa162_and0 | f_s_dadda_rca16_fa162_and1;
  assign f_s_dadda_rca16_fa163_xor0 = f_s_dadda_rca16_fa162_or0 ^ f_s_dadda_rca16_fa130_xor1;
  assign f_s_dadda_rca16_fa163_and0 = f_s_dadda_rca16_fa162_or0 & f_s_dadda_rca16_fa130_xor1;
  assign f_s_dadda_rca16_fa163_xor1 = f_s_dadda_rca16_fa163_xor0 ^ f_s_dadda_rca16_fa131_xor1;
  assign f_s_dadda_rca16_fa163_and1 = f_s_dadda_rca16_fa163_xor0 & f_s_dadda_rca16_fa131_xor1;
  assign f_s_dadda_rca16_fa163_or0 = f_s_dadda_rca16_fa163_and0 | f_s_dadda_rca16_fa163_and1;
  assign f_s_dadda_rca16_fa164_xor0 = f_s_dadda_rca16_fa163_or0 ^ f_s_dadda_rca16_fa134_xor1;
  assign f_s_dadda_rca16_fa164_and0 = f_s_dadda_rca16_fa163_or0 & f_s_dadda_rca16_fa134_xor1;
  assign f_s_dadda_rca16_fa164_xor1 = f_s_dadda_rca16_fa164_xor0 ^ f_s_dadda_rca16_fa135_xor1;
  assign f_s_dadda_rca16_fa164_and1 = f_s_dadda_rca16_fa164_xor0 & f_s_dadda_rca16_fa135_xor1;
  assign f_s_dadda_rca16_fa164_or0 = f_s_dadda_rca16_fa164_and0 | f_s_dadda_rca16_fa164_and1;
  assign f_s_dadda_rca16_nand_10_15 = ~(a[10] & b[15]);
  assign f_s_dadda_rca16_fa165_xor0 = f_s_dadda_rca16_fa164_or0 ^ f_s_dadda_rca16_nand_10_15;
  assign f_s_dadda_rca16_fa165_and0 = f_s_dadda_rca16_fa164_or0 & f_s_dadda_rca16_nand_10_15;
  assign f_s_dadda_rca16_fa165_xor1 = f_s_dadda_rca16_fa165_xor0 ^ f_s_dadda_rca16_fa138_xor1;
  assign f_s_dadda_rca16_fa165_and1 = f_s_dadda_rca16_fa165_xor0 & f_s_dadda_rca16_fa138_xor1;
  assign f_s_dadda_rca16_fa165_or0 = f_s_dadda_rca16_fa165_and0 | f_s_dadda_rca16_fa165_and1;
  assign f_s_dadda_rca16_and_12_14 = a[12] & b[14];
  assign f_s_dadda_rca16_nand_11_15 = ~(a[11] & b[15]);
  assign f_s_dadda_rca16_fa166_xor0 = f_s_dadda_rca16_fa165_or0 ^ f_s_dadda_rca16_and_12_14;
  assign f_s_dadda_rca16_fa166_and0 = f_s_dadda_rca16_fa165_or0 & f_s_dadda_rca16_and_12_14;
  assign f_s_dadda_rca16_fa166_xor1 = f_s_dadda_rca16_fa166_xor0 ^ f_s_dadda_rca16_nand_11_15;
  assign f_s_dadda_rca16_fa166_and1 = f_s_dadda_rca16_fa166_xor0 & f_s_dadda_rca16_nand_11_15;
  assign f_s_dadda_rca16_fa166_or0 = f_s_dadda_rca16_fa166_and0 | f_s_dadda_rca16_fa166_and1;
  assign f_s_dadda_rca16_and_14_13 = a[14] & b[13];
  assign f_s_dadda_rca16_and_13_14 = a[13] & b[14];
  assign f_s_dadda_rca16_fa167_xor0 = f_s_dadda_rca16_fa166_or0 ^ f_s_dadda_rca16_and_14_13;
  assign f_s_dadda_rca16_fa167_and0 = f_s_dadda_rca16_fa166_or0 & f_s_dadda_rca16_and_14_13;
  assign f_s_dadda_rca16_fa167_xor1 = f_s_dadda_rca16_fa167_xor0 ^ f_s_dadda_rca16_and_13_14;
  assign f_s_dadda_rca16_fa167_and1 = f_s_dadda_rca16_fa167_xor0 & f_s_dadda_rca16_and_13_14;
  assign f_s_dadda_rca16_fa167_or0 = f_s_dadda_rca16_fa167_and0 | f_s_dadda_rca16_fa167_and1;
  assign f_s_dadda_rca16_nand_15_13 = ~(a[15] & b[13]);
  assign f_s_dadda_rca16_fa168_xor0 = f_s_dadda_rca16_fa167_or0 ^ f_s_dadda_rca16_fa143_or0;
  assign f_s_dadda_rca16_fa168_and0 = f_s_dadda_rca16_fa167_or0 & f_s_dadda_rca16_fa143_or0;
  assign f_s_dadda_rca16_fa168_xor1 = f_s_dadda_rca16_fa168_xor0 ^ f_s_dadda_rca16_nand_15_13;
  assign f_s_dadda_rca16_fa168_and1 = f_s_dadda_rca16_fa168_xor0 & f_s_dadda_rca16_nand_15_13;
  assign f_s_dadda_rca16_fa168_or0 = f_s_dadda_rca16_fa168_and0 | f_s_dadda_rca16_fa168_and1;
  assign f_s_dadda_rca16_and_2_0 = a[2] & b[0];
  assign f_s_dadda_rca16_and_1_1 = a[1] & b[1];
  assign f_s_dadda_rca16_ha13_xor0 = f_s_dadda_rca16_and_2_0 ^ f_s_dadda_rca16_and_1_1;
  assign f_s_dadda_rca16_ha13_and0 = f_s_dadda_rca16_and_2_0 & f_s_dadda_rca16_and_1_1;
  assign f_s_dadda_rca16_and_1_2 = a[1] & b[2];
  assign f_s_dadda_rca16_and_0_3 = a[0] & b[3];
  assign f_s_dadda_rca16_fa169_xor0 = f_s_dadda_rca16_ha13_and0 ^ f_s_dadda_rca16_and_1_2;
  assign f_s_dadda_rca16_fa169_and0 = f_s_dadda_rca16_ha13_and0 & f_s_dadda_rca16_and_1_2;
  assign f_s_dadda_rca16_fa169_xor1 = f_s_dadda_rca16_fa169_xor0 ^ f_s_dadda_rca16_and_0_3;
  assign f_s_dadda_rca16_fa169_and1 = f_s_dadda_rca16_fa169_xor0 & f_s_dadda_rca16_and_0_3;
  assign f_s_dadda_rca16_fa169_or0 = f_s_dadda_rca16_fa169_and0 | f_s_dadda_rca16_fa169_and1;
  assign f_s_dadda_rca16_and_0_4 = a[0] & b[4];
  assign f_s_dadda_rca16_fa170_xor0 = f_s_dadda_rca16_fa169_or0 ^ f_s_dadda_rca16_and_0_4;
  assign f_s_dadda_rca16_fa170_and0 = f_s_dadda_rca16_fa169_or0 & f_s_dadda_rca16_and_0_4;
  assign f_s_dadda_rca16_fa170_xor1 = f_s_dadda_rca16_fa170_xor0 ^ f_s_dadda_rca16_ha3_xor0;
  assign f_s_dadda_rca16_fa170_and1 = f_s_dadda_rca16_fa170_xor0 & f_s_dadda_rca16_ha3_xor0;
  assign f_s_dadda_rca16_fa170_or0 = f_s_dadda_rca16_fa170_and0 | f_s_dadda_rca16_fa170_and1;
  assign f_s_dadda_rca16_fa171_xor0 = f_s_dadda_rca16_fa170_or0 ^ f_s_dadda_rca16_fa9_xor1;
  assign f_s_dadda_rca16_fa171_and0 = f_s_dadda_rca16_fa170_or0 & f_s_dadda_rca16_fa9_xor1;
  assign f_s_dadda_rca16_fa171_xor1 = f_s_dadda_rca16_fa171_xor0 ^ f_s_dadda_rca16_ha4_xor0;
  assign f_s_dadda_rca16_fa171_and1 = f_s_dadda_rca16_fa171_xor0 & f_s_dadda_rca16_ha4_xor0;
  assign f_s_dadda_rca16_fa171_or0 = f_s_dadda_rca16_fa171_and0 | f_s_dadda_rca16_fa171_and1;
  assign f_s_dadda_rca16_fa172_xor0 = f_s_dadda_rca16_fa171_or0 ^ f_s_dadda_rca16_fa11_xor1;
  assign f_s_dadda_rca16_fa172_and0 = f_s_dadda_rca16_fa171_or0 & f_s_dadda_rca16_fa11_xor1;
  assign f_s_dadda_rca16_fa172_xor1 = f_s_dadda_rca16_fa172_xor0 ^ f_s_dadda_rca16_ha5_xor0;
  assign f_s_dadda_rca16_fa172_and1 = f_s_dadda_rca16_fa172_xor0 & f_s_dadda_rca16_ha5_xor0;
  assign f_s_dadda_rca16_fa172_or0 = f_s_dadda_rca16_fa172_and0 | f_s_dadda_rca16_fa172_and1;
  assign f_s_dadda_rca16_fa173_xor0 = f_s_dadda_rca16_fa172_or0 ^ f_s_dadda_rca16_fa14_xor1;
  assign f_s_dadda_rca16_fa173_and0 = f_s_dadda_rca16_fa172_or0 & f_s_dadda_rca16_fa14_xor1;
  assign f_s_dadda_rca16_fa173_xor1 = f_s_dadda_rca16_fa173_xor0 ^ f_s_dadda_rca16_ha6_xor0;
  assign f_s_dadda_rca16_fa173_and1 = f_s_dadda_rca16_fa173_xor0 & f_s_dadda_rca16_ha6_xor0;
  assign f_s_dadda_rca16_fa173_or0 = f_s_dadda_rca16_fa173_and0 | f_s_dadda_rca16_fa173_and1;
  assign f_s_dadda_rca16_fa174_xor0 = f_s_dadda_rca16_fa173_or0 ^ f_s_dadda_rca16_fa18_xor1;
  assign f_s_dadda_rca16_fa174_and0 = f_s_dadda_rca16_fa173_or0 & f_s_dadda_rca16_fa18_xor1;
  assign f_s_dadda_rca16_fa174_xor1 = f_s_dadda_rca16_fa174_xor0 ^ f_s_dadda_rca16_ha7_xor0;
  assign f_s_dadda_rca16_fa174_and1 = f_s_dadda_rca16_fa174_xor0 & f_s_dadda_rca16_ha7_xor0;
  assign f_s_dadda_rca16_fa174_or0 = f_s_dadda_rca16_fa174_and0 | f_s_dadda_rca16_fa174_and1;
  assign f_s_dadda_rca16_fa175_xor0 = f_s_dadda_rca16_fa174_or0 ^ f_s_dadda_rca16_fa23_xor1;
  assign f_s_dadda_rca16_fa175_and0 = f_s_dadda_rca16_fa174_or0 & f_s_dadda_rca16_fa23_xor1;
  assign f_s_dadda_rca16_fa175_xor1 = f_s_dadda_rca16_fa175_xor0 ^ f_s_dadda_rca16_ha8_xor0;
  assign f_s_dadda_rca16_fa175_and1 = f_s_dadda_rca16_fa175_xor0 & f_s_dadda_rca16_ha8_xor0;
  assign f_s_dadda_rca16_fa175_or0 = f_s_dadda_rca16_fa175_and0 | f_s_dadda_rca16_fa175_and1;
  assign f_s_dadda_rca16_fa176_xor0 = f_s_dadda_rca16_fa175_or0 ^ f_s_dadda_rca16_fa29_xor1;
  assign f_s_dadda_rca16_fa176_and0 = f_s_dadda_rca16_fa175_or0 & f_s_dadda_rca16_fa29_xor1;
  assign f_s_dadda_rca16_fa176_xor1 = f_s_dadda_rca16_fa176_xor0 ^ f_s_dadda_rca16_ha9_xor0;
  assign f_s_dadda_rca16_fa176_and1 = f_s_dadda_rca16_fa176_xor0 & f_s_dadda_rca16_ha9_xor0;
  assign f_s_dadda_rca16_fa176_or0 = f_s_dadda_rca16_fa176_and0 | f_s_dadda_rca16_fa176_and1;
  assign f_s_dadda_rca16_fa177_xor0 = f_s_dadda_rca16_fa176_or0 ^ f_s_dadda_rca16_fa36_xor1;
  assign f_s_dadda_rca16_fa177_and0 = f_s_dadda_rca16_fa176_or0 & f_s_dadda_rca16_fa36_xor1;
  assign f_s_dadda_rca16_fa177_xor1 = f_s_dadda_rca16_fa177_xor0 ^ f_s_dadda_rca16_ha10_xor0;
  assign f_s_dadda_rca16_fa177_and1 = f_s_dadda_rca16_fa177_xor0 & f_s_dadda_rca16_ha10_xor0;
  assign f_s_dadda_rca16_fa177_or0 = f_s_dadda_rca16_fa177_and0 | f_s_dadda_rca16_fa177_and1;
  assign f_s_dadda_rca16_fa178_xor0 = f_s_dadda_rca16_fa177_or0 ^ f_s_dadda_rca16_fa44_xor1;
  assign f_s_dadda_rca16_fa178_and0 = f_s_dadda_rca16_fa177_or0 & f_s_dadda_rca16_fa44_xor1;
  assign f_s_dadda_rca16_fa178_xor1 = f_s_dadda_rca16_fa178_xor0 ^ f_s_dadda_rca16_ha11_xor0;
  assign f_s_dadda_rca16_fa178_and1 = f_s_dadda_rca16_fa178_xor0 & f_s_dadda_rca16_ha11_xor0;
  assign f_s_dadda_rca16_fa178_or0 = f_s_dadda_rca16_fa178_and0 | f_s_dadda_rca16_fa178_and1;
  assign f_s_dadda_rca16_fa179_xor0 = f_s_dadda_rca16_fa178_or0 ^ f_s_dadda_rca16_fa52_xor1;
  assign f_s_dadda_rca16_fa179_and0 = f_s_dadda_rca16_fa178_or0 & f_s_dadda_rca16_fa52_xor1;
  assign f_s_dadda_rca16_fa179_xor1 = f_s_dadda_rca16_fa179_xor0 ^ f_s_dadda_rca16_fa53_xor1;
  assign f_s_dadda_rca16_fa179_and1 = f_s_dadda_rca16_fa179_xor0 & f_s_dadda_rca16_fa53_xor1;
  assign f_s_dadda_rca16_fa179_or0 = f_s_dadda_rca16_fa179_and0 | f_s_dadda_rca16_fa179_and1;
  assign f_s_dadda_rca16_fa180_xor0 = f_s_dadda_rca16_fa179_or0 ^ f_s_dadda_rca16_fa61_xor1;
  assign f_s_dadda_rca16_fa180_and0 = f_s_dadda_rca16_fa179_or0 & f_s_dadda_rca16_fa61_xor1;
  assign f_s_dadda_rca16_fa180_xor1 = f_s_dadda_rca16_fa180_xor0 ^ f_s_dadda_rca16_fa62_xor1;
  assign f_s_dadda_rca16_fa180_and1 = f_s_dadda_rca16_fa180_xor0 & f_s_dadda_rca16_fa62_xor1;
  assign f_s_dadda_rca16_fa180_or0 = f_s_dadda_rca16_fa180_and0 | f_s_dadda_rca16_fa180_and1;
  assign f_s_dadda_rca16_fa181_xor0 = f_s_dadda_rca16_fa180_or0 ^ f_s_dadda_rca16_fa70_xor1;
  assign f_s_dadda_rca16_fa181_and0 = f_s_dadda_rca16_fa180_or0 & f_s_dadda_rca16_fa70_xor1;
  assign f_s_dadda_rca16_fa181_xor1 = f_s_dadda_rca16_fa181_xor0 ^ f_s_dadda_rca16_fa71_xor1;
  assign f_s_dadda_rca16_fa181_and1 = f_s_dadda_rca16_fa181_xor0 & f_s_dadda_rca16_fa71_xor1;
  assign f_s_dadda_rca16_fa181_or0 = f_s_dadda_rca16_fa181_and0 | f_s_dadda_rca16_fa181_and1;
  assign f_s_dadda_rca16_fa182_xor0 = f_s_dadda_rca16_fa181_or0 ^ f_s_dadda_rca16_fa79_xor1;
  assign f_s_dadda_rca16_fa182_and0 = f_s_dadda_rca16_fa181_or0 & f_s_dadda_rca16_fa79_xor1;
  assign f_s_dadda_rca16_fa182_xor1 = f_s_dadda_rca16_fa182_xor0 ^ f_s_dadda_rca16_fa80_xor1;
  assign f_s_dadda_rca16_fa182_and1 = f_s_dadda_rca16_fa182_xor0 & f_s_dadda_rca16_fa80_xor1;
  assign f_s_dadda_rca16_fa182_or0 = f_s_dadda_rca16_fa182_and0 | f_s_dadda_rca16_fa182_and1;
  assign f_s_dadda_rca16_fa183_xor0 = f_s_dadda_rca16_fa182_or0 ^ f_s_dadda_rca16_fa88_xor1;
  assign f_s_dadda_rca16_fa183_and0 = f_s_dadda_rca16_fa182_or0 & f_s_dadda_rca16_fa88_xor1;
  assign f_s_dadda_rca16_fa183_xor1 = f_s_dadda_rca16_fa183_xor0 ^ f_s_dadda_rca16_fa89_xor1;
  assign f_s_dadda_rca16_fa183_and1 = f_s_dadda_rca16_fa183_xor0 & f_s_dadda_rca16_fa89_xor1;
  assign f_s_dadda_rca16_fa183_or0 = f_s_dadda_rca16_fa183_and0 | f_s_dadda_rca16_fa183_and1;
  assign f_s_dadda_rca16_fa184_xor0 = f_s_dadda_rca16_fa183_or0 ^ f_s_dadda_rca16_fa97_xor1;
  assign f_s_dadda_rca16_fa184_and0 = f_s_dadda_rca16_fa183_or0 & f_s_dadda_rca16_fa97_xor1;
  assign f_s_dadda_rca16_fa184_xor1 = f_s_dadda_rca16_fa184_xor0 ^ f_s_dadda_rca16_fa98_xor1;
  assign f_s_dadda_rca16_fa184_and1 = f_s_dadda_rca16_fa184_xor0 & f_s_dadda_rca16_fa98_xor1;
  assign f_s_dadda_rca16_fa184_or0 = f_s_dadda_rca16_fa184_and0 | f_s_dadda_rca16_fa184_and1;
  assign f_s_dadda_rca16_fa185_xor0 = f_s_dadda_rca16_fa184_or0 ^ f_s_dadda_rca16_fa106_xor1;
  assign f_s_dadda_rca16_fa185_and0 = f_s_dadda_rca16_fa184_or0 & f_s_dadda_rca16_fa106_xor1;
  assign f_s_dadda_rca16_fa185_xor1 = f_s_dadda_rca16_fa185_xor0 ^ f_s_dadda_rca16_fa107_xor1;
  assign f_s_dadda_rca16_fa185_and1 = f_s_dadda_rca16_fa185_xor0 & f_s_dadda_rca16_fa107_xor1;
  assign f_s_dadda_rca16_fa185_or0 = f_s_dadda_rca16_fa185_and0 | f_s_dadda_rca16_fa185_and1;
  assign f_s_dadda_rca16_fa186_xor0 = f_s_dadda_rca16_fa185_or0 ^ f_s_dadda_rca16_fa114_xor1;
  assign f_s_dadda_rca16_fa186_and0 = f_s_dadda_rca16_fa185_or0 & f_s_dadda_rca16_fa114_xor1;
  assign f_s_dadda_rca16_fa186_xor1 = f_s_dadda_rca16_fa186_xor0 ^ f_s_dadda_rca16_fa115_xor1;
  assign f_s_dadda_rca16_fa186_and1 = f_s_dadda_rca16_fa186_xor0 & f_s_dadda_rca16_fa115_xor1;
  assign f_s_dadda_rca16_fa186_or0 = f_s_dadda_rca16_fa186_and0 | f_s_dadda_rca16_fa186_and1;
  assign f_s_dadda_rca16_fa187_xor0 = f_s_dadda_rca16_fa186_or0 ^ f_s_dadda_rca16_fa121_xor1;
  assign f_s_dadda_rca16_fa187_and0 = f_s_dadda_rca16_fa186_or0 & f_s_dadda_rca16_fa121_xor1;
  assign f_s_dadda_rca16_fa187_xor1 = f_s_dadda_rca16_fa187_xor0 ^ f_s_dadda_rca16_fa122_xor1;
  assign f_s_dadda_rca16_fa187_and1 = f_s_dadda_rca16_fa187_xor0 & f_s_dadda_rca16_fa122_xor1;
  assign f_s_dadda_rca16_fa187_or0 = f_s_dadda_rca16_fa187_and0 | f_s_dadda_rca16_fa187_and1;
  assign f_s_dadda_rca16_fa188_xor0 = f_s_dadda_rca16_fa187_or0 ^ f_s_dadda_rca16_fa127_xor1;
  assign f_s_dadda_rca16_fa188_and0 = f_s_dadda_rca16_fa187_or0 & f_s_dadda_rca16_fa127_xor1;
  assign f_s_dadda_rca16_fa188_xor1 = f_s_dadda_rca16_fa188_xor0 ^ f_s_dadda_rca16_fa128_xor1;
  assign f_s_dadda_rca16_fa188_and1 = f_s_dadda_rca16_fa188_xor0 & f_s_dadda_rca16_fa128_xor1;
  assign f_s_dadda_rca16_fa188_or0 = f_s_dadda_rca16_fa188_and0 | f_s_dadda_rca16_fa188_and1;
  assign f_s_dadda_rca16_fa189_xor0 = f_s_dadda_rca16_fa188_or0 ^ f_s_dadda_rca16_fa132_xor1;
  assign f_s_dadda_rca16_fa189_and0 = f_s_dadda_rca16_fa188_or0 & f_s_dadda_rca16_fa132_xor1;
  assign f_s_dadda_rca16_fa189_xor1 = f_s_dadda_rca16_fa189_xor0 ^ f_s_dadda_rca16_fa133_xor1;
  assign f_s_dadda_rca16_fa189_and1 = f_s_dadda_rca16_fa189_xor0 & f_s_dadda_rca16_fa133_xor1;
  assign f_s_dadda_rca16_fa189_or0 = f_s_dadda_rca16_fa189_and0 | f_s_dadda_rca16_fa189_and1;
  assign f_s_dadda_rca16_fa190_xor0 = f_s_dadda_rca16_fa189_or0 ^ f_s_dadda_rca16_fa136_xor1;
  assign f_s_dadda_rca16_fa190_and0 = f_s_dadda_rca16_fa189_or0 & f_s_dadda_rca16_fa136_xor1;
  assign f_s_dadda_rca16_fa190_xor1 = f_s_dadda_rca16_fa190_xor0 ^ f_s_dadda_rca16_fa137_xor1;
  assign f_s_dadda_rca16_fa190_and1 = f_s_dadda_rca16_fa190_xor0 & f_s_dadda_rca16_fa137_xor1;
  assign f_s_dadda_rca16_fa190_or0 = f_s_dadda_rca16_fa190_and0 | f_s_dadda_rca16_fa190_and1;
  assign f_s_dadda_rca16_fa191_xor0 = f_s_dadda_rca16_fa190_or0 ^ f_s_dadda_rca16_fa139_xor1;
  assign f_s_dadda_rca16_fa191_and0 = f_s_dadda_rca16_fa190_or0 & f_s_dadda_rca16_fa139_xor1;
  assign f_s_dadda_rca16_fa191_xor1 = f_s_dadda_rca16_fa191_xor0 ^ f_s_dadda_rca16_fa140_xor1;
  assign f_s_dadda_rca16_fa191_and1 = f_s_dadda_rca16_fa191_xor0 & f_s_dadda_rca16_fa140_xor1;
  assign f_s_dadda_rca16_fa191_or0 = f_s_dadda_rca16_fa191_and0 | f_s_dadda_rca16_fa191_and1;
  assign f_s_dadda_rca16_fa192_xor0 = f_s_dadda_rca16_fa191_or0 ^ f_s_dadda_rca16_fa141_xor1;
  assign f_s_dadda_rca16_fa192_and0 = f_s_dadda_rca16_fa191_or0 & f_s_dadda_rca16_fa141_xor1;
  assign f_s_dadda_rca16_fa192_xor1 = f_s_dadda_rca16_fa192_xor0 ^ f_s_dadda_rca16_fa142_xor1;
  assign f_s_dadda_rca16_fa192_and1 = f_s_dadda_rca16_fa192_xor0 & f_s_dadda_rca16_fa142_xor1;
  assign f_s_dadda_rca16_fa192_or0 = f_s_dadda_rca16_fa192_and0 | f_s_dadda_rca16_fa192_and1;
  assign f_s_dadda_rca16_nand_12_15 = ~(a[12] & b[15]);
  assign f_s_dadda_rca16_fa193_xor0 = f_s_dadda_rca16_fa192_or0 ^ f_s_dadda_rca16_nand_12_15;
  assign f_s_dadda_rca16_fa193_and0 = f_s_dadda_rca16_fa192_or0 & f_s_dadda_rca16_nand_12_15;
  assign f_s_dadda_rca16_fa193_xor1 = f_s_dadda_rca16_fa193_xor0 ^ f_s_dadda_rca16_fa143_xor1;
  assign f_s_dadda_rca16_fa193_and1 = f_s_dadda_rca16_fa193_xor0 & f_s_dadda_rca16_fa143_xor1;
  assign f_s_dadda_rca16_fa193_or0 = f_s_dadda_rca16_fa193_and0 | f_s_dadda_rca16_fa193_and1;
  assign f_s_dadda_rca16_and_14_14 = a[14] & b[14];
  assign f_s_dadda_rca16_nand_13_15 = ~(a[13] & b[15]);
  assign f_s_dadda_rca16_fa194_xor0 = f_s_dadda_rca16_fa193_or0 ^ f_s_dadda_rca16_and_14_14;
  assign f_s_dadda_rca16_fa194_and0 = f_s_dadda_rca16_fa193_or0 & f_s_dadda_rca16_and_14_14;
  assign f_s_dadda_rca16_fa194_xor1 = f_s_dadda_rca16_fa194_xor0 ^ f_s_dadda_rca16_nand_13_15;
  assign f_s_dadda_rca16_fa194_and1 = f_s_dadda_rca16_fa194_xor0 & f_s_dadda_rca16_nand_13_15;
  assign f_s_dadda_rca16_fa194_or0 = f_s_dadda_rca16_fa194_and0 | f_s_dadda_rca16_fa194_and1;
  assign f_s_dadda_rca16_nand_15_14 = ~(a[15] & b[14]);
  assign f_s_dadda_rca16_fa195_xor0 = f_s_dadda_rca16_fa194_or0 ^ f_s_dadda_rca16_fa168_or0;
  assign f_s_dadda_rca16_fa195_and0 = f_s_dadda_rca16_fa194_or0 & f_s_dadda_rca16_fa168_or0;
  assign f_s_dadda_rca16_fa195_xor1 = f_s_dadda_rca16_fa195_xor0 ^ f_s_dadda_rca16_nand_15_14;
  assign f_s_dadda_rca16_fa195_and1 = f_s_dadda_rca16_fa195_xor0 & f_s_dadda_rca16_nand_15_14;
  assign f_s_dadda_rca16_fa195_or0 = f_s_dadda_rca16_fa195_and0 | f_s_dadda_rca16_fa195_and1;
  assign f_s_dadda_rca16_and_0_0 = a[0] & b[0];
  assign f_s_dadda_rca16_and_1_0 = a[1] & b[0];
  assign f_s_dadda_rca16_and_0_2 = a[0] & b[2];
  assign f_s_dadda_rca16_nand_14_15 = ~(a[14] & b[15]);
  assign f_s_dadda_rca16_and_0_1 = a[0] & b[1];
  assign f_s_dadda_rca16_and_15_15 = a[15] & b[15];
  assign f_s_dadda_rca16_u_rca30_ha_xor0 = f_s_dadda_rca16_and_1_0 ^ f_s_dadda_rca16_and_0_1;
  assign f_s_dadda_rca16_u_rca30_ha_and0 = f_s_dadda_rca16_and_1_0 & f_s_dadda_rca16_and_0_1;
  assign f_s_dadda_rca16_u_rca30_fa1_xor0 = f_s_dadda_rca16_and_0_2 ^ f_s_dadda_rca16_ha13_xor0;
  assign f_s_dadda_rca16_u_rca30_fa1_and0 = f_s_dadda_rca16_and_0_2 & f_s_dadda_rca16_ha13_xor0;
  assign f_s_dadda_rca16_u_rca30_fa1_xor1 = f_s_dadda_rca16_u_rca30_fa1_xor0 ^ f_s_dadda_rca16_u_rca30_ha_and0;
  assign f_s_dadda_rca16_u_rca30_fa1_and1 = f_s_dadda_rca16_u_rca30_fa1_xor0 & f_s_dadda_rca16_u_rca30_ha_and0;
  assign f_s_dadda_rca16_u_rca30_fa1_or0 = f_s_dadda_rca16_u_rca30_fa1_and0 | f_s_dadda_rca16_u_rca30_fa1_and1;
  assign f_s_dadda_rca16_u_rca30_fa2_xor0 = f_s_dadda_rca16_ha12_xor0 ^ f_s_dadda_rca16_fa169_xor1;
  assign f_s_dadda_rca16_u_rca30_fa2_and0 = f_s_dadda_rca16_ha12_xor0 & f_s_dadda_rca16_fa169_xor1;
  assign f_s_dadda_rca16_u_rca30_fa2_xor1 = f_s_dadda_rca16_u_rca30_fa2_xor0 ^ f_s_dadda_rca16_u_rca30_fa1_or0;
  assign f_s_dadda_rca16_u_rca30_fa2_and1 = f_s_dadda_rca16_u_rca30_fa2_xor0 & f_s_dadda_rca16_u_rca30_fa1_or0;
  assign f_s_dadda_rca16_u_rca30_fa2_or0 = f_s_dadda_rca16_u_rca30_fa2_and0 | f_s_dadda_rca16_u_rca30_fa2_and1;
  assign f_s_dadda_rca16_u_rca30_fa3_xor0 = f_s_dadda_rca16_fa144_xor1 ^ f_s_dadda_rca16_fa170_xor1;
  assign f_s_dadda_rca16_u_rca30_fa3_and0 = f_s_dadda_rca16_fa144_xor1 & f_s_dadda_rca16_fa170_xor1;
  assign f_s_dadda_rca16_u_rca30_fa3_xor1 = f_s_dadda_rca16_u_rca30_fa3_xor0 ^ f_s_dadda_rca16_u_rca30_fa2_or0;
  assign f_s_dadda_rca16_u_rca30_fa3_and1 = f_s_dadda_rca16_u_rca30_fa3_xor0 & f_s_dadda_rca16_u_rca30_fa2_or0;
  assign f_s_dadda_rca16_u_rca30_fa3_or0 = f_s_dadda_rca16_u_rca30_fa3_and0 | f_s_dadda_rca16_u_rca30_fa3_and1;
  assign f_s_dadda_rca16_u_rca30_fa4_xor0 = f_s_dadda_rca16_fa145_xor1 ^ f_s_dadda_rca16_fa171_xor1;
  assign f_s_dadda_rca16_u_rca30_fa4_and0 = f_s_dadda_rca16_fa145_xor1 & f_s_dadda_rca16_fa171_xor1;
  assign f_s_dadda_rca16_u_rca30_fa4_xor1 = f_s_dadda_rca16_u_rca30_fa4_xor0 ^ f_s_dadda_rca16_u_rca30_fa3_or0;
  assign f_s_dadda_rca16_u_rca30_fa4_and1 = f_s_dadda_rca16_u_rca30_fa4_xor0 & f_s_dadda_rca16_u_rca30_fa3_or0;
  assign f_s_dadda_rca16_u_rca30_fa4_or0 = f_s_dadda_rca16_u_rca30_fa4_and0 | f_s_dadda_rca16_u_rca30_fa4_and1;
  assign f_s_dadda_rca16_u_rca30_fa5_xor0 = f_s_dadda_rca16_fa146_xor1 ^ f_s_dadda_rca16_fa172_xor1;
  assign f_s_dadda_rca16_u_rca30_fa5_and0 = f_s_dadda_rca16_fa146_xor1 & f_s_dadda_rca16_fa172_xor1;
  assign f_s_dadda_rca16_u_rca30_fa5_xor1 = f_s_dadda_rca16_u_rca30_fa5_xor0 ^ f_s_dadda_rca16_u_rca30_fa4_or0;
  assign f_s_dadda_rca16_u_rca30_fa5_and1 = f_s_dadda_rca16_u_rca30_fa5_xor0 & f_s_dadda_rca16_u_rca30_fa4_or0;
  assign f_s_dadda_rca16_u_rca30_fa5_or0 = f_s_dadda_rca16_u_rca30_fa5_and0 | f_s_dadda_rca16_u_rca30_fa5_and1;
  assign f_s_dadda_rca16_u_rca30_fa6_xor0 = f_s_dadda_rca16_fa147_xor1 ^ f_s_dadda_rca16_fa173_xor1;
  assign f_s_dadda_rca16_u_rca30_fa6_and0 = f_s_dadda_rca16_fa147_xor1 & f_s_dadda_rca16_fa173_xor1;
  assign f_s_dadda_rca16_u_rca30_fa6_xor1 = f_s_dadda_rca16_u_rca30_fa6_xor0 ^ f_s_dadda_rca16_u_rca30_fa5_or0;
  assign f_s_dadda_rca16_u_rca30_fa6_and1 = f_s_dadda_rca16_u_rca30_fa6_xor0 & f_s_dadda_rca16_u_rca30_fa5_or0;
  assign f_s_dadda_rca16_u_rca30_fa6_or0 = f_s_dadda_rca16_u_rca30_fa6_and0 | f_s_dadda_rca16_u_rca30_fa6_and1;
  assign f_s_dadda_rca16_u_rca30_fa7_xor0 = f_s_dadda_rca16_fa148_xor1 ^ f_s_dadda_rca16_fa174_xor1;
  assign f_s_dadda_rca16_u_rca30_fa7_and0 = f_s_dadda_rca16_fa148_xor1 & f_s_dadda_rca16_fa174_xor1;
  assign f_s_dadda_rca16_u_rca30_fa7_xor1 = f_s_dadda_rca16_u_rca30_fa7_xor0 ^ f_s_dadda_rca16_u_rca30_fa6_or0;
  assign f_s_dadda_rca16_u_rca30_fa7_and1 = f_s_dadda_rca16_u_rca30_fa7_xor0 & f_s_dadda_rca16_u_rca30_fa6_or0;
  assign f_s_dadda_rca16_u_rca30_fa7_or0 = f_s_dadda_rca16_u_rca30_fa7_and0 | f_s_dadda_rca16_u_rca30_fa7_and1;
  assign f_s_dadda_rca16_u_rca30_fa8_xor0 = f_s_dadda_rca16_fa149_xor1 ^ f_s_dadda_rca16_fa175_xor1;
  assign f_s_dadda_rca16_u_rca30_fa8_and0 = f_s_dadda_rca16_fa149_xor1 & f_s_dadda_rca16_fa175_xor1;
  assign f_s_dadda_rca16_u_rca30_fa8_xor1 = f_s_dadda_rca16_u_rca30_fa8_xor0 ^ f_s_dadda_rca16_u_rca30_fa7_or0;
  assign f_s_dadda_rca16_u_rca30_fa8_and1 = f_s_dadda_rca16_u_rca30_fa8_xor0 & f_s_dadda_rca16_u_rca30_fa7_or0;
  assign f_s_dadda_rca16_u_rca30_fa8_or0 = f_s_dadda_rca16_u_rca30_fa8_and0 | f_s_dadda_rca16_u_rca30_fa8_and1;
  assign f_s_dadda_rca16_u_rca30_fa9_xor0 = f_s_dadda_rca16_fa150_xor1 ^ f_s_dadda_rca16_fa176_xor1;
  assign f_s_dadda_rca16_u_rca30_fa9_and0 = f_s_dadda_rca16_fa150_xor1 & f_s_dadda_rca16_fa176_xor1;
  assign f_s_dadda_rca16_u_rca30_fa9_xor1 = f_s_dadda_rca16_u_rca30_fa9_xor0 ^ f_s_dadda_rca16_u_rca30_fa8_or0;
  assign f_s_dadda_rca16_u_rca30_fa9_and1 = f_s_dadda_rca16_u_rca30_fa9_xor0 & f_s_dadda_rca16_u_rca30_fa8_or0;
  assign f_s_dadda_rca16_u_rca30_fa9_or0 = f_s_dadda_rca16_u_rca30_fa9_and0 | f_s_dadda_rca16_u_rca30_fa9_and1;
  assign f_s_dadda_rca16_u_rca30_fa10_xor0 = f_s_dadda_rca16_fa151_xor1 ^ f_s_dadda_rca16_fa177_xor1;
  assign f_s_dadda_rca16_u_rca30_fa10_and0 = f_s_dadda_rca16_fa151_xor1 & f_s_dadda_rca16_fa177_xor1;
  assign f_s_dadda_rca16_u_rca30_fa10_xor1 = f_s_dadda_rca16_u_rca30_fa10_xor0 ^ f_s_dadda_rca16_u_rca30_fa9_or0;
  assign f_s_dadda_rca16_u_rca30_fa10_and1 = f_s_dadda_rca16_u_rca30_fa10_xor0 & f_s_dadda_rca16_u_rca30_fa9_or0;
  assign f_s_dadda_rca16_u_rca30_fa10_or0 = f_s_dadda_rca16_u_rca30_fa10_and0 | f_s_dadda_rca16_u_rca30_fa10_and1;
  assign f_s_dadda_rca16_u_rca30_fa11_xor0 = f_s_dadda_rca16_fa152_xor1 ^ f_s_dadda_rca16_fa178_xor1;
  assign f_s_dadda_rca16_u_rca30_fa11_and0 = f_s_dadda_rca16_fa152_xor1 & f_s_dadda_rca16_fa178_xor1;
  assign f_s_dadda_rca16_u_rca30_fa11_xor1 = f_s_dadda_rca16_u_rca30_fa11_xor0 ^ f_s_dadda_rca16_u_rca30_fa10_or0;
  assign f_s_dadda_rca16_u_rca30_fa11_and1 = f_s_dadda_rca16_u_rca30_fa11_xor0 & f_s_dadda_rca16_u_rca30_fa10_or0;
  assign f_s_dadda_rca16_u_rca30_fa11_or0 = f_s_dadda_rca16_u_rca30_fa11_and0 | f_s_dadda_rca16_u_rca30_fa11_and1;
  assign f_s_dadda_rca16_u_rca30_fa12_xor0 = f_s_dadda_rca16_fa153_xor1 ^ f_s_dadda_rca16_fa179_xor1;
  assign f_s_dadda_rca16_u_rca30_fa12_and0 = f_s_dadda_rca16_fa153_xor1 & f_s_dadda_rca16_fa179_xor1;
  assign f_s_dadda_rca16_u_rca30_fa12_xor1 = f_s_dadda_rca16_u_rca30_fa12_xor0 ^ f_s_dadda_rca16_u_rca30_fa11_or0;
  assign f_s_dadda_rca16_u_rca30_fa12_and1 = f_s_dadda_rca16_u_rca30_fa12_xor0 & f_s_dadda_rca16_u_rca30_fa11_or0;
  assign f_s_dadda_rca16_u_rca30_fa12_or0 = f_s_dadda_rca16_u_rca30_fa12_and0 | f_s_dadda_rca16_u_rca30_fa12_and1;
  assign f_s_dadda_rca16_u_rca30_fa13_xor0 = f_s_dadda_rca16_fa154_xor1 ^ f_s_dadda_rca16_fa180_xor1;
  assign f_s_dadda_rca16_u_rca30_fa13_and0 = f_s_dadda_rca16_fa154_xor1 & f_s_dadda_rca16_fa180_xor1;
  assign f_s_dadda_rca16_u_rca30_fa13_xor1 = f_s_dadda_rca16_u_rca30_fa13_xor0 ^ f_s_dadda_rca16_u_rca30_fa12_or0;
  assign f_s_dadda_rca16_u_rca30_fa13_and1 = f_s_dadda_rca16_u_rca30_fa13_xor0 & f_s_dadda_rca16_u_rca30_fa12_or0;
  assign f_s_dadda_rca16_u_rca30_fa13_or0 = f_s_dadda_rca16_u_rca30_fa13_and0 | f_s_dadda_rca16_u_rca30_fa13_and1;
  assign f_s_dadda_rca16_u_rca30_fa14_xor0 = f_s_dadda_rca16_fa155_xor1 ^ f_s_dadda_rca16_fa181_xor1;
  assign f_s_dadda_rca16_u_rca30_fa14_and0 = f_s_dadda_rca16_fa155_xor1 & f_s_dadda_rca16_fa181_xor1;
  assign f_s_dadda_rca16_u_rca30_fa14_xor1 = f_s_dadda_rca16_u_rca30_fa14_xor0 ^ f_s_dadda_rca16_u_rca30_fa13_or0;
  assign f_s_dadda_rca16_u_rca30_fa14_and1 = f_s_dadda_rca16_u_rca30_fa14_xor0 & f_s_dadda_rca16_u_rca30_fa13_or0;
  assign f_s_dadda_rca16_u_rca30_fa14_or0 = f_s_dadda_rca16_u_rca30_fa14_and0 | f_s_dadda_rca16_u_rca30_fa14_and1;
  assign f_s_dadda_rca16_u_rca30_fa15_xor0 = f_s_dadda_rca16_fa156_xor1 ^ f_s_dadda_rca16_fa182_xor1;
  assign f_s_dadda_rca16_u_rca30_fa15_and0 = f_s_dadda_rca16_fa156_xor1 & f_s_dadda_rca16_fa182_xor1;
  assign f_s_dadda_rca16_u_rca30_fa15_xor1 = f_s_dadda_rca16_u_rca30_fa15_xor0 ^ f_s_dadda_rca16_u_rca30_fa14_or0;
  assign f_s_dadda_rca16_u_rca30_fa15_and1 = f_s_dadda_rca16_u_rca30_fa15_xor0 & f_s_dadda_rca16_u_rca30_fa14_or0;
  assign f_s_dadda_rca16_u_rca30_fa15_or0 = f_s_dadda_rca16_u_rca30_fa15_and0 | f_s_dadda_rca16_u_rca30_fa15_and1;
  assign f_s_dadda_rca16_u_rca30_fa16_xor0 = f_s_dadda_rca16_fa157_xor1 ^ f_s_dadda_rca16_fa183_xor1;
  assign f_s_dadda_rca16_u_rca30_fa16_and0 = f_s_dadda_rca16_fa157_xor1 & f_s_dadda_rca16_fa183_xor1;
  assign f_s_dadda_rca16_u_rca30_fa16_xor1 = f_s_dadda_rca16_u_rca30_fa16_xor0 ^ f_s_dadda_rca16_u_rca30_fa15_or0;
  assign f_s_dadda_rca16_u_rca30_fa16_and1 = f_s_dadda_rca16_u_rca30_fa16_xor0 & f_s_dadda_rca16_u_rca30_fa15_or0;
  assign f_s_dadda_rca16_u_rca30_fa16_or0 = f_s_dadda_rca16_u_rca30_fa16_and0 | f_s_dadda_rca16_u_rca30_fa16_and1;
  assign f_s_dadda_rca16_u_rca30_fa17_xor0 = f_s_dadda_rca16_fa158_xor1 ^ f_s_dadda_rca16_fa184_xor1;
  assign f_s_dadda_rca16_u_rca30_fa17_and0 = f_s_dadda_rca16_fa158_xor1 & f_s_dadda_rca16_fa184_xor1;
  assign f_s_dadda_rca16_u_rca30_fa17_xor1 = f_s_dadda_rca16_u_rca30_fa17_xor0 ^ f_s_dadda_rca16_u_rca30_fa16_or0;
  assign f_s_dadda_rca16_u_rca30_fa17_and1 = f_s_dadda_rca16_u_rca30_fa17_xor0 & f_s_dadda_rca16_u_rca30_fa16_or0;
  assign f_s_dadda_rca16_u_rca30_fa17_or0 = f_s_dadda_rca16_u_rca30_fa17_and0 | f_s_dadda_rca16_u_rca30_fa17_and1;
  assign f_s_dadda_rca16_u_rca30_fa18_xor0 = f_s_dadda_rca16_fa159_xor1 ^ f_s_dadda_rca16_fa185_xor1;
  assign f_s_dadda_rca16_u_rca30_fa18_and0 = f_s_dadda_rca16_fa159_xor1 & f_s_dadda_rca16_fa185_xor1;
  assign f_s_dadda_rca16_u_rca30_fa18_xor1 = f_s_dadda_rca16_u_rca30_fa18_xor0 ^ f_s_dadda_rca16_u_rca30_fa17_or0;
  assign f_s_dadda_rca16_u_rca30_fa18_and1 = f_s_dadda_rca16_u_rca30_fa18_xor0 & f_s_dadda_rca16_u_rca30_fa17_or0;
  assign f_s_dadda_rca16_u_rca30_fa18_or0 = f_s_dadda_rca16_u_rca30_fa18_and0 | f_s_dadda_rca16_u_rca30_fa18_and1;
  assign f_s_dadda_rca16_u_rca30_fa19_xor0 = f_s_dadda_rca16_fa160_xor1 ^ f_s_dadda_rca16_fa186_xor1;
  assign f_s_dadda_rca16_u_rca30_fa19_and0 = f_s_dadda_rca16_fa160_xor1 & f_s_dadda_rca16_fa186_xor1;
  assign f_s_dadda_rca16_u_rca30_fa19_xor1 = f_s_dadda_rca16_u_rca30_fa19_xor0 ^ f_s_dadda_rca16_u_rca30_fa18_or0;
  assign f_s_dadda_rca16_u_rca30_fa19_and1 = f_s_dadda_rca16_u_rca30_fa19_xor0 & f_s_dadda_rca16_u_rca30_fa18_or0;
  assign f_s_dadda_rca16_u_rca30_fa19_or0 = f_s_dadda_rca16_u_rca30_fa19_and0 | f_s_dadda_rca16_u_rca30_fa19_and1;
  assign f_s_dadda_rca16_u_rca30_fa20_xor0 = f_s_dadda_rca16_fa161_xor1 ^ f_s_dadda_rca16_fa187_xor1;
  assign f_s_dadda_rca16_u_rca30_fa20_and0 = f_s_dadda_rca16_fa161_xor1 & f_s_dadda_rca16_fa187_xor1;
  assign f_s_dadda_rca16_u_rca30_fa20_xor1 = f_s_dadda_rca16_u_rca30_fa20_xor0 ^ f_s_dadda_rca16_u_rca30_fa19_or0;
  assign f_s_dadda_rca16_u_rca30_fa20_and1 = f_s_dadda_rca16_u_rca30_fa20_xor0 & f_s_dadda_rca16_u_rca30_fa19_or0;
  assign f_s_dadda_rca16_u_rca30_fa20_or0 = f_s_dadda_rca16_u_rca30_fa20_and0 | f_s_dadda_rca16_u_rca30_fa20_and1;
  assign f_s_dadda_rca16_u_rca30_fa21_xor0 = f_s_dadda_rca16_fa162_xor1 ^ f_s_dadda_rca16_fa188_xor1;
  assign f_s_dadda_rca16_u_rca30_fa21_and0 = f_s_dadda_rca16_fa162_xor1 & f_s_dadda_rca16_fa188_xor1;
  assign f_s_dadda_rca16_u_rca30_fa21_xor1 = f_s_dadda_rca16_u_rca30_fa21_xor0 ^ f_s_dadda_rca16_u_rca30_fa20_or0;
  assign f_s_dadda_rca16_u_rca30_fa21_and1 = f_s_dadda_rca16_u_rca30_fa21_xor0 & f_s_dadda_rca16_u_rca30_fa20_or0;
  assign f_s_dadda_rca16_u_rca30_fa21_or0 = f_s_dadda_rca16_u_rca30_fa21_and0 | f_s_dadda_rca16_u_rca30_fa21_and1;
  assign f_s_dadda_rca16_u_rca30_fa22_xor0 = f_s_dadda_rca16_fa163_xor1 ^ f_s_dadda_rca16_fa189_xor1;
  assign f_s_dadda_rca16_u_rca30_fa22_and0 = f_s_dadda_rca16_fa163_xor1 & f_s_dadda_rca16_fa189_xor1;
  assign f_s_dadda_rca16_u_rca30_fa22_xor1 = f_s_dadda_rca16_u_rca30_fa22_xor0 ^ f_s_dadda_rca16_u_rca30_fa21_or0;
  assign f_s_dadda_rca16_u_rca30_fa22_and1 = f_s_dadda_rca16_u_rca30_fa22_xor0 & f_s_dadda_rca16_u_rca30_fa21_or0;
  assign f_s_dadda_rca16_u_rca30_fa22_or0 = f_s_dadda_rca16_u_rca30_fa22_and0 | f_s_dadda_rca16_u_rca30_fa22_and1;
  assign f_s_dadda_rca16_u_rca30_fa23_xor0 = f_s_dadda_rca16_fa164_xor1 ^ f_s_dadda_rca16_fa190_xor1;
  assign f_s_dadda_rca16_u_rca30_fa23_and0 = f_s_dadda_rca16_fa164_xor1 & f_s_dadda_rca16_fa190_xor1;
  assign f_s_dadda_rca16_u_rca30_fa23_xor1 = f_s_dadda_rca16_u_rca30_fa23_xor0 ^ f_s_dadda_rca16_u_rca30_fa22_or0;
  assign f_s_dadda_rca16_u_rca30_fa23_and1 = f_s_dadda_rca16_u_rca30_fa23_xor0 & f_s_dadda_rca16_u_rca30_fa22_or0;
  assign f_s_dadda_rca16_u_rca30_fa23_or0 = f_s_dadda_rca16_u_rca30_fa23_and0 | f_s_dadda_rca16_u_rca30_fa23_and1;
  assign f_s_dadda_rca16_u_rca30_fa24_xor0 = f_s_dadda_rca16_fa165_xor1 ^ f_s_dadda_rca16_fa191_xor1;
  assign f_s_dadda_rca16_u_rca30_fa24_and0 = f_s_dadda_rca16_fa165_xor1 & f_s_dadda_rca16_fa191_xor1;
  assign f_s_dadda_rca16_u_rca30_fa24_xor1 = f_s_dadda_rca16_u_rca30_fa24_xor0 ^ f_s_dadda_rca16_u_rca30_fa23_or0;
  assign f_s_dadda_rca16_u_rca30_fa24_and1 = f_s_dadda_rca16_u_rca30_fa24_xor0 & f_s_dadda_rca16_u_rca30_fa23_or0;
  assign f_s_dadda_rca16_u_rca30_fa24_or0 = f_s_dadda_rca16_u_rca30_fa24_and0 | f_s_dadda_rca16_u_rca30_fa24_and1;
  assign f_s_dadda_rca16_u_rca30_fa25_xor0 = f_s_dadda_rca16_fa166_xor1 ^ f_s_dadda_rca16_fa192_xor1;
  assign f_s_dadda_rca16_u_rca30_fa25_and0 = f_s_dadda_rca16_fa166_xor1 & f_s_dadda_rca16_fa192_xor1;
  assign f_s_dadda_rca16_u_rca30_fa25_xor1 = f_s_dadda_rca16_u_rca30_fa25_xor0 ^ f_s_dadda_rca16_u_rca30_fa24_or0;
  assign f_s_dadda_rca16_u_rca30_fa25_and1 = f_s_dadda_rca16_u_rca30_fa25_xor0 & f_s_dadda_rca16_u_rca30_fa24_or0;
  assign f_s_dadda_rca16_u_rca30_fa25_or0 = f_s_dadda_rca16_u_rca30_fa25_and0 | f_s_dadda_rca16_u_rca30_fa25_and1;
  assign f_s_dadda_rca16_u_rca30_fa26_xor0 = f_s_dadda_rca16_fa167_xor1 ^ f_s_dadda_rca16_fa193_xor1;
  assign f_s_dadda_rca16_u_rca30_fa26_and0 = f_s_dadda_rca16_fa167_xor1 & f_s_dadda_rca16_fa193_xor1;
  assign f_s_dadda_rca16_u_rca30_fa26_xor1 = f_s_dadda_rca16_u_rca30_fa26_xor0 ^ f_s_dadda_rca16_u_rca30_fa25_or0;
  assign f_s_dadda_rca16_u_rca30_fa26_and1 = f_s_dadda_rca16_u_rca30_fa26_xor0 & f_s_dadda_rca16_u_rca30_fa25_or0;
  assign f_s_dadda_rca16_u_rca30_fa26_or0 = f_s_dadda_rca16_u_rca30_fa26_and0 | f_s_dadda_rca16_u_rca30_fa26_and1;
  assign f_s_dadda_rca16_u_rca30_fa27_xor0 = f_s_dadda_rca16_fa168_xor1 ^ f_s_dadda_rca16_fa194_xor1;
  assign f_s_dadda_rca16_u_rca30_fa27_and0 = f_s_dadda_rca16_fa168_xor1 & f_s_dadda_rca16_fa194_xor1;
  assign f_s_dadda_rca16_u_rca30_fa27_xor1 = f_s_dadda_rca16_u_rca30_fa27_xor0 ^ f_s_dadda_rca16_u_rca30_fa26_or0;
  assign f_s_dadda_rca16_u_rca30_fa27_and1 = f_s_dadda_rca16_u_rca30_fa27_xor0 & f_s_dadda_rca16_u_rca30_fa26_or0;
  assign f_s_dadda_rca16_u_rca30_fa27_or0 = f_s_dadda_rca16_u_rca30_fa27_and0 | f_s_dadda_rca16_u_rca30_fa27_and1;
  assign f_s_dadda_rca16_u_rca30_fa28_xor0 = f_s_dadda_rca16_nand_14_15 ^ f_s_dadda_rca16_fa195_xor1;
  assign f_s_dadda_rca16_u_rca30_fa28_and0 = f_s_dadda_rca16_nand_14_15 & f_s_dadda_rca16_fa195_xor1;
  assign f_s_dadda_rca16_u_rca30_fa28_xor1 = f_s_dadda_rca16_u_rca30_fa28_xor0 ^ f_s_dadda_rca16_u_rca30_fa27_or0;
  assign f_s_dadda_rca16_u_rca30_fa28_and1 = f_s_dadda_rca16_u_rca30_fa28_xor0 & f_s_dadda_rca16_u_rca30_fa27_or0;
  assign f_s_dadda_rca16_u_rca30_fa28_or0 = f_s_dadda_rca16_u_rca30_fa28_and0 | f_s_dadda_rca16_u_rca30_fa28_and1;
  assign f_s_dadda_rca16_u_rca30_fa29_xor0 = f_s_dadda_rca16_fa195_or0 ^ f_s_dadda_rca16_and_15_15;
  assign f_s_dadda_rca16_u_rca30_fa29_and0 = f_s_dadda_rca16_fa195_or0 & f_s_dadda_rca16_and_15_15;
  assign f_s_dadda_rca16_u_rca30_fa29_xor1 = f_s_dadda_rca16_u_rca30_fa29_xor0 ^ f_s_dadda_rca16_u_rca30_fa28_or0;
  assign f_s_dadda_rca16_u_rca30_fa29_and1 = f_s_dadda_rca16_u_rca30_fa29_xor0 & f_s_dadda_rca16_u_rca30_fa28_or0;
  assign f_s_dadda_rca16_u_rca30_fa29_or0 = f_s_dadda_rca16_u_rca30_fa29_and0 | f_s_dadda_rca16_u_rca30_fa29_and1;
  assign f_s_dadda_rca16_xor0 = ~f_s_dadda_rca16_u_rca30_fa29_or0;

  assign f_s_dadda_rca16_out[0] = f_s_dadda_rca16_and_0_0;
  assign f_s_dadda_rca16_out[1] = f_s_dadda_rca16_u_rca30_ha_xor0;
  assign f_s_dadda_rca16_out[2] = f_s_dadda_rca16_u_rca30_fa1_xor1;
  assign f_s_dadda_rca16_out[3] = f_s_dadda_rca16_u_rca30_fa2_xor1;
  assign f_s_dadda_rca16_out[4] = f_s_dadda_rca16_u_rca30_fa3_xor1;
  assign f_s_dadda_rca16_out[5] = f_s_dadda_rca16_u_rca30_fa4_xor1;
  assign f_s_dadda_rca16_out[6] = f_s_dadda_rca16_u_rca30_fa5_xor1;
  assign f_s_dadda_rca16_out[7] = f_s_dadda_rca16_u_rca30_fa6_xor1;
  assign f_s_dadda_rca16_out[8] = f_s_dadda_rca16_u_rca30_fa7_xor1;
  assign f_s_dadda_rca16_out[9] = f_s_dadda_rca16_u_rca30_fa8_xor1;
  assign f_s_dadda_rca16_out[10] = f_s_dadda_rca16_u_rca30_fa9_xor1;
  assign f_s_dadda_rca16_out[11] = f_s_dadda_rca16_u_rca30_fa10_xor1;
  assign f_s_dadda_rca16_out[12] = f_s_dadda_rca16_u_rca30_fa11_xor1;
  assign f_s_dadda_rca16_out[13] = f_s_dadda_rca16_u_rca30_fa12_xor1;
  assign f_s_dadda_rca16_out[14] = f_s_dadda_rca16_u_rca30_fa13_xor1;
  assign f_s_dadda_rca16_out[15] = f_s_dadda_rca16_u_rca30_fa14_xor1;
  assign f_s_dadda_rca16_out[16] = f_s_dadda_rca16_u_rca30_fa15_xor1;
  assign f_s_dadda_rca16_out[17] = f_s_dadda_rca16_u_rca30_fa16_xor1;
  assign f_s_dadda_rca16_out[18] = f_s_dadda_rca16_u_rca30_fa17_xor1;
  assign f_s_dadda_rca16_out[19] = f_s_dadda_rca16_u_rca30_fa18_xor1;
  assign f_s_dadda_rca16_out[20] = f_s_dadda_rca16_u_rca30_fa19_xor1;
  assign f_s_dadda_rca16_out[21] = f_s_dadda_rca16_u_rca30_fa20_xor1;
  assign f_s_dadda_rca16_out[22] = f_s_dadda_rca16_u_rca30_fa21_xor1;
  assign f_s_dadda_rca16_out[23] = f_s_dadda_rca16_u_rca30_fa22_xor1;
  assign f_s_dadda_rca16_out[24] = f_s_dadda_rca16_u_rca30_fa23_xor1;
  assign f_s_dadda_rca16_out[25] = f_s_dadda_rca16_u_rca30_fa24_xor1;
  assign f_s_dadda_rca16_out[26] = f_s_dadda_rca16_u_rca30_fa25_xor1;
  assign f_s_dadda_rca16_out[27] = f_s_dadda_rca16_u_rca30_fa26_xor1;
  assign f_s_dadda_rca16_out[28] = f_s_dadda_rca16_u_rca30_fa27_xor1;
  assign f_s_dadda_rca16_out[29] = f_s_dadda_rca16_u_rca30_fa28_xor1;
  assign f_s_dadda_rca16_out[30] = f_s_dadda_rca16_u_rca30_fa29_xor1;
  assign f_s_dadda_rca16_out[31] = f_s_dadda_rca16_xor0;
endmodule