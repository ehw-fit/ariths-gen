module f_u_arrmul12(input [11:0] a, input [11:0] b, output [23:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire f_u_arrmul12_and0_0_a_0;
  wire f_u_arrmul12_and0_0_b_0;
  wire f_u_arrmul12_and0_0_y0;
  wire f_u_arrmul12_and1_0_a_1;
  wire f_u_arrmul12_and1_0_b_0;
  wire f_u_arrmul12_and1_0_y0;
  wire f_u_arrmul12_and2_0_a_2;
  wire f_u_arrmul12_and2_0_b_0;
  wire f_u_arrmul12_and2_0_y0;
  wire f_u_arrmul12_and3_0_a_3;
  wire f_u_arrmul12_and3_0_b_0;
  wire f_u_arrmul12_and3_0_y0;
  wire f_u_arrmul12_and4_0_a_4;
  wire f_u_arrmul12_and4_0_b_0;
  wire f_u_arrmul12_and4_0_y0;
  wire f_u_arrmul12_and5_0_a_5;
  wire f_u_arrmul12_and5_0_b_0;
  wire f_u_arrmul12_and5_0_y0;
  wire f_u_arrmul12_and6_0_a_6;
  wire f_u_arrmul12_and6_0_b_0;
  wire f_u_arrmul12_and6_0_y0;
  wire f_u_arrmul12_and7_0_a_7;
  wire f_u_arrmul12_and7_0_b_0;
  wire f_u_arrmul12_and7_0_y0;
  wire f_u_arrmul12_and8_0_a_8;
  wire f_u_arrmul12_and8_0_b_0;
  wire f_u_arrmul12_and8_0_y0;
  wire f_u_arrmul12_and9_0_a_9;
  wire f_u_arrmul12_and9_0_b_0;
  wire f_u_arrmul12_and9_0_y0;
  wire f_u_arrmul12_and10_0_a_10;
  wire f_u_arrmul12_and10_0_b_0;
  wire f_u_arrmul12_and10_0_y0;
  wire f_u_arrmul12_and11_0_a_11;
  wire f_u_arrmul12_and11_0_b_0;
  wire f_u_arrmul12_and11_0_y0;
  wire f_u_arrmul12_and0_1_a_0;
  wire f_u_arrmul12_and0_1_b_1;
  wire f_u_arrmul12_and0_1_y0;
  wire f_u_arrmul12_ha0_1_f_u_arrmul12_and0_1_y0;
  wire f_u_arrmul12_ha0_1_f_u_arrmul12_and1_0_y0;
  wire f_u_arrmul12_ha0_1_y0;
  wire f_u_arrmul12_ha0_1_y1;
  wire f_u_arrmul12_and1_1_a_1;
  wire f_u_arrmul12_and1_1_b_1;
  wire f_u_arrmul12_and1_1_y0;
  wire f_u_arrmul12_fa1_1_f_u_arrmul12_and1_1_y0;
  wire f_u_arrmul12_fa1_1_f_u_arrmul12_and2_0_y0;
  wire f_u_arrmul12_fa1_1_y0;
  wire f_u_arrmul12_fa1_1_y1;
  wire f_u_arrmul12_fa1_1_f_u_arrmul12_ha0_1_y1;
  wire f_u_arrmul12_fa1_1_y2;
  wire f_u_arrmul12_fa1_1_y3;
  wire f_u_arrmul12_fa1_1_y4;
  wire f_u_arrmul12_and2_1_a_2;
  wire f_u_arrmul12_and2_1_b_1;
  wire f_u_arrmul12_and2_1_y0;
  wire f_u_arrmul12_fa2_1_f_u_arrmul12_and2_1_y0;
  wire f_u_arrmul12_fa2_1_f_u_arrmul12_and3_0_y0;
  wire f_u_arrmul12_fa2_1_y0;
  wire f_u_arrmul12_fa2_1_y1;
  wire f_u_arrmul12_fa2_1_f_u_arrmul12_fa1_1_y4;
  wire f_u_arrmul12_fa2_1_y2;
  wire f_u_arrmul12_fa2_1_y3;
  wire f_u_arrmul12_fa2_1_y4;
  wire f_u_arrmul12_and3_1_a_3;
  wire f_u_arrmul12_and3_1_b_1;
  wire f_u_arrmul12_and3_1_y0;
  wire f_u_arrmul12_fa3_1_f_u_arrmul12_and3_1_y0;
  wire f_u_arrmul12_fa3_1_f_u_arrmul12_and4_0_y0;
  wire f_u_arrmul12_fa3_1_y0;
  wire f_u_arrmul12_fa3_1_y1;
  wire f_u_arrmul12_fa3_1_f_u_arrmul12_fa2_1_y4;
  wire f_u_arrmul12_fa3_1_y2;
  wire f_u_arrmul12_fa3_1_y3;
  wire f_u_arrmul12_fa3_1_y4;
  wire f_u_arrmul12_and4_1_a_4;
  wire f_u_arrmul12_and4_1_b_1;
  wire f_u_arrmul12_and4_1_y0;
  wire f_u_arrmul12_fa4_1_f_u_arrmul12_and4_1_y0;
  wire f_u_arrmul12_fa4_1_f_u_arrmul12_and5_0_y0;
  wire f_u_arrmul12_fa4_1_y0;
  wire f_u_arrmul12_fa4_1_y1;
  wire f_u_arrmul12_fa4_1_f_u_arrmul12_fa3_1_y4;
  wire f_u_arrmul12_fa4_1_y2;
  wire f_u_arrmul12_fa4_1_y3;
  wire f_u_arrmul12_fa4_1_y4;
  wire f_u_arrmul12_and5_1_a_5;
  wire f_u_arrmul12_and5_1_b_1;
  wire f_u_arrmul12_and5_1_y0;
  wire f_u_arrmul12_fa5_1_f_u_arrmul12_and5_1_y0;
  wire f_u_arrmul12_fa5_1_f_u_arrmul12_and6_0_y0;
  wire f_u_arrmul12_fa5_1_y0;
  wire f_u_arrmul12_fa5_1_y1;
  wire f_u_arrmul12_fa5_1_f_u_arrmul12_fa4_1_y4;
  wire f_u_arrmul12_fa5_1_y2;
  wire f_u_arrmul12_fa5_1_y3;
  wire f_u_arrmul12_fa5_1_y4;
  wire f_u_arrmul12_and6_1_a_6;
  wire f_u_arrmul12_and6_1_b_1;
  wire f_u_arrmul12_and6_1_y0;
  wire f_u_arrmul12_fa6_1_f_u_arrmul12_and6_1_y0;
  wire f_u_arrmul12_fa6_1_f_u_arrmul12_and7_0_y0;
  wire f_u_arrmul12_fa6_1_y0;
  wire f_u_arrmul12_fa6_1_y1;
  wire f_u_arrmul12_fa6_1_f_u_arrmul12_fa5_1_y4;
  wire f_u_arrmul12_fa6_1_y2;
  wire f_u_arrmul12_fa6_1_y3;
  wire f_u_arrmul12_fa6_1_y4;
  wire f_u_arrmul12_and7_1_a_7;
  wire f_u_arrmul12_and7_1_b_1;
  wire f_u_arrmul12_and7_1_y0;
  wire f_u_arrmul12_fa7_1_f_u_arrmul12_and7_1_y0;
  wire f_u_arrmul12_fa7_1_f_u_arrmul12_and8_0_y0;
  wire f_u_arrmul12_fa7_1_y0;
  wire f_u_arrmul12_fa7_1_y1;
  wire f_u_arrmul12_fa7_1_f_u_arrmul12_fa6_1_y4;
  wire f_u_arrmul12_fa7_1_y2;
  wire f_u_arrmul12_fa7_1_y3;
  wire f_u_arrmul12_fa7_1_y4;
  wire f_u_arrmul12_and8_1_a_8;
  wire f_u_arrmul12_and8_1_b_1;
  wire f_u_arrmul12_and8_1_y0;
  wire f_u_arrmul12_fa8_1_f_u_arrmul12_and8_1_y0;
  wire f_u_arrmul12_fa8_1_f_u_arrmul12_and9_0_y0;
  wire f_u_arrmul12_fa8_1_y0;
  wire f_u_arrmul12_fa8_1_y1;
  wire f_u_arrmul12_fa8_1_f_u_arrmul12_fa7_1_y4;
  wire f_u_arrmul12_fa8_1_y2;
  wire f_u_arrmul12_fa8_1_y3;
  wire f_u_arrmul12_fa8_1_y4;
  wire f_u_arrmul12_and9_1_a_9;
  wire f_u_arrmul12_and9_1_b_1;
  wire f_u_arrmul12_and9_1_y0;
  wire f_u_arrmul12_fa9_1_f_u_arrmul12_and9_1_y0;
  wire f_u_arrmul12_fa9_1_f_u_arrmul12_and10_0_y0;
  wire f_u_arrmul12_fa9_1_y0;
  wire f_u_arrmul12_fa9_1_y1;
  wire f_u_arrmul12_fa9_1_f_u_arrmul12_fa8_1_y4;
  wire f_u_arrmul12_fa9_1_y2;
  wire f_u_arrmul12_fa9_1_y3;
  wire f_u_arrmul12_fa9_1_y4;
  wire f_u_arrmul12_and10_1_a_10;
  wire f_u_arrmul12_and10_1_b_1;
  wire f_u_arrmul12_and10_1_y0;
  wire f_u_arrmul12_fa10_1_f_u_arrmul12_and10_1_y0;
  wire f_u_arrmul12_fa10_1_f_u_arrmul12_and11_0_y0;
  wire f_u_arrmul12_fa10_1_y0;
  wire f_u_arrmul12_fa10_1_y1;
  wire f_u_arrmul12_fa10_1_f_u_arrmul12_fa9_1_y4;
  wire f_u_arrmul12_fa10_1_y2;
  wire f_u_arrmul12_fa10_1_y3;
  wire f_u_arrmul12_fa10_1_y4;
  wire f_u_arrmul12_and11_1_a_11;
  wire f_u_arrmul12_and11_1_b_1;
  wire f_u_arrmul12_and11_1_y0;
  wire f_u_arrmul12_ha11_1_f_u_arrmul12_and11_1_y0;
  wire f_u_arrmul12_ha11_1_f_u_arrmul12_fa10_1_y4;
  wire f_u_arrmul12_ha11_1_y0;
  wire f_u_arrmul12_ha11_1_y1;
  wire f_u_arrmul12_and0_2_a_0;
  wire f_u_arrmul12_and0_2_b_2;
  wire f_u_arrmul12_and0_2_y0;
  wire f_u_arrmul12_ha0_2_f_u_arrmul12_and0_2_y0;
  wire f_u_arrmul12_ha0_2_f_u_arrmul12_fa1_1_y2;
  wire f_u_arrmul12_ha0_2_y0;
  wire f_u_arrmul12_ha0_2_y1;
  wire f_u_arrmul12_and1_2_a_1;
  wire f_u_arrmul12_and1_2_b_2;
  wire f_u_arrmul12_and1_2_y0;
  wire f_u_arrmul12_fa1_2_f_u_arrmul12_and1_2_y0;
  wire f_u_arrmul12_fa1_2_f_u_arrmul12_fa2_1_y2;
  wire f_u_arrmul12_fa1_2_y0;
  wire f_u_arrmul12_fa1_2_y1;
  wire f_u_arrmul12_fa1_2_f_u_arrmul12_ha0_2_y1;
  wire f_u_arrmul12_fa1_2_y2;
  wire f_u_arrmul12_fa1_2_y3;
  wire f_u_arrmul12_fa1_2_y4;
  wire f_u_arrmul12_and2_2_a_2;
  wire f_u_arrmul12_and2_2_b_2;
  wire f_u_arrmul12_and2_2_y0;
  wire f_u_arrmul12_fa2_2_f_u_arrmul12_and2_2_y0;
  wire f_u_arrmul12_fa2_2_f_u_arrmul12_fa3_1_y2;
  wire f_u_arrmul12_fa2_2_y0;
  wire f_u_arrmul12_fa2_2_y1;
  wire f_u_arrmul12_fa2_2_f_u_arrmul12_fa1_2_y4;
  wire f_u_arrmul12_fa2_2_y2;
  wire f_u_arrmul12_fa2_2_y3;
  wire f_u_arrmul12_fa2_2_y4;
  wire f_u_arrmul12_and3_2_a_3;
  wire f_u_arrmul12_and3_2_b_2;
  wire f_u_arrmul12_and3_2_y0;
  wire f_u_arrmul12_fa3_2_f_u_arrmul12_and3_2_y0;
  wire f_u_arrmul12_fa3_2_f_u_arrmul12_fa4_1_y2;
  wire f_u_arrmul12_fa3_2_y0;
  wire f_u_arrmul12_fa3_2_y1;
  wire f_u_arrmul12_fa3_2_f_u_arrmul12_fa2_2_y4;
  wire f_u_arrmul12_fa3_2_y2;
  wire f_u_arrmul12_fa3_2_y3;
  wire f_u_arrmul12_fa3_2_y4;
  wire f_u_arrmul12_and4_2_a_4;
  wire f_u_arrmul12_and4_2_b_2;
  wire f_u_arrmul12_and4_2_y0;
  wire f_u_arrmul12_fa4_2_f_u_arrmul12_and4_2_y0;
  wire f_u_arrmul12_fa4_2_f_u_arrmul12_fa5_1_y2;
  wire f_u_arrmul12_fa4_2_y0;
  wire f_u_arrmul12_fa4_2_y1;
  wire f_u_arrmul12_fa4_2_f_u_arrmul12_fa3_2_y4;
  wire f_u_arrmul12_fa4_2_y2;
  wire f_u_arrmul12_fa4_2_y3;
  wire f_u_arrmul12_fa4_2_y4;
  wire f_u_arrmul12_and5_2_a_5;
  wire f_u_arrmul12_and5_2_b_2;
  wire f_u_arrmul12_and5_2_y0;
  wire f_u_arrmul12_fa5_2_f_u_arrmul12_and5_2_y0;
  wire f_u_arrmul12_fa5_2_f_u_arrmul12_fa6_1_y2;
  wire f_u_arrmul12_fa5_2_y0;
  wire f_u_arrmul12_fa5_2_y1;
  wire f_u_arrmul12_fa5_2_f_u_arrmul12_fa4_2_y4;
  wire f_u_arrmul12_fa5_2_y2;
  wire f_u_arrmul12_fa5_2_y3;
  wire f_u_arrmul12_fa5_2_y4;
  wire f_u_arrmul12_and6_2_a_6;
  wire f_u_arrmul12_and6_2_b_2;
  wire f_u_arrmul12_and6_2_y0;
  wire f_u_arrmul12_fa6_2_f_u_arrmul12_and6_2_y0;
  wire f_u_arrmul12_fa6_2_f_u_arrmul12_fa7_1_y2;
  wire f_u_arrmul12_fa6_2_y0;
  wire f_u_arrmul12_fa6_2_y1;
  wire f_u_arrmul12_fa6_2_f_u_arrmul12_fa5_2_y4;
  wire f_u_arrmul12_fa6_2_y2;
  wire f_u_arrmul12_fa6_2_y3;
  wire f_u_arrmul12_fa6_2_y4;
  wire f_u_arrmul12_and7_2_a_7;
  wire f_u_arrmul12_and7_2_b_2;
  wire f_u_arrmul12_and7_2_y0;
  wire f_u_arrmul12_fa7_2_f_u_arrmul12_and7_2_y0;
  wire f_u_arrmul12_fa7_2_f_u_arrmul12_fa8_1_y2;
  wire f_u_arrmul12_fa7_2_y0;
  wire f_u_arrmul12_fa7_2_y1;
  wire f_u_arrmul12_fa7_2_f_u_arrmul12_fa6_2_y4;
  wire f_u_arrmul12_fa7_2_y2;
  wire f_u_arrmul12_fa7_2_y3;
  wire f_u_arrmul12_fa7_2_y4;
  wire f_u_arrmul12_and8_2_a_8;
  wire f_u_arrmul12_and8_2_b_2;
  wire f_u_arrmul12_and8_2_y0;
  wire f_u_arrmul12_fa8_2_f_u_arrmul12_and8_2_y0;
  wire f_u_arrmul12_fa8_2_f_u_arrmul12_fa9_1_y2;
  wire f_u_arrmul12_fa8_2_y0;
  wire f_u_arrmul12_fa8_2_y1;
  wire f_u_arrmul12_fa8_2_f_u_arrmul12_fa7_2_y4;
  wire f_u_arrmul12_fa8_2_y2;
  wire f_u_arrmul12_fa8_2_y3;
  wire f_u_arrmul12_fa8_2_y4;
  wire f_u_arrmul12_and9_2_a_9;
  wire f_u_arrmul12_and9_2_b_2;
  wire f_u_arrmul12_and9_2_y0;
  wire f_u_arrmul12_fa9_2_f_u_arrmul12_and9_2_y0;
  wire f_u_arrmul12_fa9_2_f_u_arrmul12_fa10_1_y2;
  wire f_u_arrmul12_fa9_2_y0;
  wire f_u_arrmul12_fa9_2_y1;
  wire f_u_arrmul12_fa9_2_f_u_arrmul12_fa8_2_y4;
  wire f_u_arrmul12_fa9_2_y2;
  wire f_u_arrmul12_fa9_2_y3;
  wire f_u_arrmul12_fa9_2_y4;
  wire f_u_arrmul12_and10_2_a_10;
  wire f_u_arrmul12_and10_2_b_2;
  wire f_u_arrmul12_and10_2_y0;
  wire f_u_arrmul12_fa10_2_f_u_arrmul12_and10_2_y0;
  wire f_u_arrmul12_fa10_2_f_u_arrmul12_ha11_1_y0;
  wire f_u_arrmul12_fa10_2_y0;
  wire f_u_arrmul12_fa10_2_y1;
  wire f_u_arrmul12_fa10_2_f_u_arrmul12_fa9_2_y4;
  wire f_u_arrmul12_fa10_2_y2;
  wire f_u_arrmul12_fa10_2_y3;
  wire f_u_arrmul12_fa10_2_y4;
  wire f_u_arrmul12_and11_2_a_11;
  wire f_u_arrmul12_and11_2_b_2;
  wire f_u_arrmul12_and11_2_y0;
  wire f_u_arrmul12_fa11_2_f_u_arrmul12_and11_2_y0;
  wire f_u_arrmul12_fa11_2_f_u_arrmul12_ha11_1_y1;
  wire f_u_arrmul12_fa11_2_y0;
  wire f_u_arrmul12_fa11_2_y1;
  wire f_u_arrmul12_fa11_2_f_u_arrmul12_fa10_2_y4;
  wire f_u_arrmul12_fa11_2_y2;
  wire f_u_arrmul12_fa11_2_y3;
  wire f_u_arrmul12_fa11_2_y4;
  wire f_u_arrmul12_and0_3_a_0;
  wire f_u_arrmul12_and0_3_b_3;
  wire f_u_arrmul12_and0_3_y0;
  wire f_u_arrmul12_ha0_3_f_u_arrmul12_and0_3_y0;
  wire f_u_arrmul12_ha0_3_f_u_arrmul12_fa1_2_y2;
  wire f_u_arrmul12_ha0_3_y0;
  wire f_u_arrmul12_ha0_3_y1;
  wire f_u_arrmul12_and1_3_a_1;
  wire f_u_arrmul12_and1_3_b_3;
  wire f_u_arrmul12_and1_3_y0;
  wire f_u_arrmul12_fa1_3_f_u_arrmul12_and1_3_y0;
  wire f_u_arrmul12_fa1_3_f_u_arrmul12_fa2_2_y2;
  wire f_u_arrmul12_fa1_3_y0;
  wire f_u_arrmul12_fa1_3_y1;
  wire f_u_arrmul12_fa1_3_f_u_arrmul12_ha0_3_y1;
  wire f_u_arrmul12_fa1_3_y2;
  wire f_u_arrmul12_fa1_3_y3;
  wire f_u_arrmul12_fa1_3_y4;
  wire f_u_arrmul12_and2_3_a_2;
  wire f_u_arrmul12_and2_3_b_3;
  wire f_u_arrmul12_and2_3_y0;
  wire f_u_arrmul12_fa2_3_f_u_arrmul12_and2_3_y0;
  wire f_u_arrmul12_fa2_3_f_u_arrmul12_fa3_2_y2;
  wire f_u_arrmul12_fa2_3_y0;
  wire f_u_arrmul12_fa2_3_y1;
  wire f_u_arrmul12_fa2_3_f_u_arrmul12_fa1_3_y4;
  wire f_u_arrmul12_fa2_3_y2;
  wire f_u_arrmul12_fa2_3_y3;
  wire f_u_arrmul12_fa2_3_y4;
  wire f_u_arrmul12_and3_3_a_3;
  wire f_u_arrmul12_and3_3_b_3;
  wire f_u_arrmul12_and3_3_y0;
  wire f_u_arrmul12_fa3_3_f_u_arrmul12_and3_3_y0;
  wire f_u_arrmul12_fa3_3_f_u_arrmul12_fa4_2_y2;
  wire f_u_arrmul12_fa3_3_y0;
  wire f_u_arrmul12_fa3_3_y1;
  wire f_u_arrmul12_fa3_3_f_u_arrmul12_fa2_3_y4;
  wire f_u_arrmul12_fa3_3_y2;
  wire f_u_arrmul12_fa3_3_y3;
  wire f_u_arrmul12_fa3_3_y4;
  wire f_u_arrmul12_and4_3_a_4;
  wire f_u_arrmul12_and4_3_b_3;
  wire f_u_arrmul12_and4_3_y0;
  wire f_u_arrmul12_fa4_3_f_u_arrmul12_and4_3_y0;
  wire f_u_arrmul12_fa4_3_f_u_arrmul12_fa5_2_y2;
  wire f_u_arrmul12_fa4_3_y0;
  wire f_u_arrmul12_fa4_3_y1;
  wire f_u_arrmul12_fa4_3_f_u_arrmul12_fa3_3_y4;
  wire f_u_arrmul12_fa4_3_y2;
  wire f_u_arrmul12_fa4_3_y3;
  wire f_u_arrmul12_fa4_3_y4;
  wire f_u_arrmul12_and5_3_a_5;
  wire f_u_arrmul12_and5_3_b_3;
  wire f_u_arrmul12_and5_3_y0;
  wire f_u_arrmul12_fa5_3_f_u_arrmul12_and5_3_y0;
  wire f_u_arrmul12_fa5_3_f_u_arrmul12_fa6_2_y2;
  wire f_u_arrmul12_fa5_3_y0;
  wire f_u_arrmul12_fa5_3_y1;
  wire f_u_arrmul12_fa5_3_f_u_arrmul12_fa4_3_y4;
  wire f_u_arrmul12_fa5_3_y2;
  wire f_u_arrmul12_fa5_3_y3;
  wire f_u_arrmul12_fa5_3_y4;
  wire f_u_arrmul12_and6_3_a_6;
  wire f_u_arrmul12_and6_3_b_3;
  wire f_u_arrmul12_and6_3_y0;
  wire f_u_arrmul12_fa6_3_f_u_arrmul12_and6_3_y0;
  wire f_u_arrmul12_fa6_3_f_u_arrmul12_fa7_2_y2;
  wire f_u_arrmul12_fa6_3_y0;
  wire f_u_arrmul12_fa6_3_y1;
  wire f_u_arrmul12_fa6_3_f_u_arrmul12_fa5_3_y4;
  wire f_u_arrmul12_fa6_3_y2;
  wire f_u_arrmul12_fa6_3_y3;
  wire f_u_arrmul12_fa6_3_y4;
  wire f_u_arrmul12_and7_3_a_7;
  wire f_u_arrmul12_and7_3_b_3;
  wire f_u_arrmul12_and7_3_y0;
  wire f_u_arrmul12_fa7_3_f_u_arrmul12_and7_3_y0;
  wire f_u_arrmul12_fa7_3_f_u_arrmul12_fa8_2_y2;
  wire f_u_arrmul12_fa7_3_y0;
  wire f_u_arrmul12_fa7_3_y1;
  wire f_u_arrmul12_fa7_3_f_u_arrmul12_fa6_3_y4;
  wire f_u_arrmul12_fa7_3_y2;
  wire f_u_arrmul12_fa7_3_y3;
  wire f_u_arrmul12_fa7_3_y4;
  wire f_u_arrmul12_and8_3_a_8;
  wire f_u_arrmul12_and8_3_b_3;
  wire f_u_arrmul12_and8_3_y0;
  wire f_u_arrmul12_fa8_3_f_u_arrmul12_and8_3_y0;
  wire f_u_arrmul12_fa8_3_f_u_arrmul12_fa9_2_y2;
  wire f_u_arrmul12_fa8_3_y0;
  wire f_u_arrmul12_fa8_3_y1;
  wire f_u_arrmul12_fa8_3_f_u_arrmul12_fa7_3_y4;
  wire f_u_arrmul12_fa8_3_y2;
  wire f_u_arrmul12_fa8_3_y3;
  wire f_u_arrmul12_fa8_3_y4;
  wire f_u_arrmul12_and9_3_a_9;
  wire f_u_arrmul12_and9_3_b_3;
  wire f_u_arrmul12_and9_3_y0;
  wire f_u_arrmul12_fa9_3_f_u_arrmul12_and9_3_y0;
  wire f_u_arrmul12_fa9_3_f_u_arrmul12_fa10_2_y2;
  wire f_u_arrmul12_fa9_3_y0;
  wire f_u_arrmul12_fa9_3_y1;
  wire f_u_arrmul12_fa9_3_f_u_arrmul12_fa8_3_y4;
  wire f_u_arrmul12_fa9_3_y2;
  wire f_u_arrmul12_fa9_3_y3;
  wire f_u_arrmul12_fa9_3_y4;
  wire f_u_arrmul12_and10_3_a_10;
  wire f_u_arrmul12_and10_3_b_3;
  wire f_u_arrmul12_and10_3_y0;
  wire f_u_arrmul12_fa10_3_f_u_arrmul12_and10_3_y0;
  wire f_u_arrmul12_fa10_3_f_u_arrmul12_fa11_2_y2;
  wire f_u_arrmul12_fa10_3_y0;
  wire f_u_arrmul12_fa10_3_y1;
  wire f_u_arrmul12_fa10_3_f_u_arrmul12_fa9_3_y4;
  wire f_u_arrmul12_fa10_3_y2;
  wire f_u_arrmul12_fa10_3_y3;
  wire f_u_arrmul12_fa10_3_y4;
  wire f_u_arrmul12_and11_3_a_11;
  wire f_u_arrmul12_and11_3_b_3;
  wire f_u_arrmul12_and11_3_y0;
  wire f_u_arrmul12_fa11_3_f_u_arrmul12_and11_3_y0;
  wire f_u_arrmul12_fa11_3_f_u_arrmul12_fa11_2_y4;
  wire f_u_arrmul12_fa11_3_y0;
  wire f_u_arrmul12_fa11_3_y1;
  wire f_u_arrmul12_fa11_3_f_u_arrmul12_fa10_3_y4;
  wire f_u_arrmul12_fa11_3_y2;
  wire f_u_arrmul12_fa11_3_y3;
  wire f_u_arrmul12_fa11_3_y4;
  wire f_u_arrmul12_and0_4_a_0;
  wire f_u_arrmul12_and0_4_b_4;
  wire f_u_arrmul12_and0_4_y0;
  wire f_u_arrmul12_ha0_4_f_u_arrmul12_and0_4_y0;
  wire f_u_arrmul12_ha0_4_f_u_arrmul12_fa1_3_y2;
  wire f_u_arrmul12_ha0_4_y0;
  wire f_u_arrmul12_ha0_4_y1;
  wire f_u_arrmul12_and1_4_a_1;
  wire f_u_arrmul12_and1_4_b_4;
  wire f_u_arrmul12_and1_4_y0;
  wire f_u_arrmul12_fa1_4_f_u_arrmul12_and1_4_y0;
  wire f_u_arrmul12_fa1_4_f_u_arrmul12_fa2_3_y2;
  wire f_u_arrmul12_fa1_4_y0;
  wire f_u_arrmul12_fa1_4_y1;
  wire f_u_arrmul12_fa1_4_f_u_arrmul12_ha0_4_y1;
  wire f_u_arrmul12_fa1_4_y2;
  wire f_u_arrmul12_fa1_4_y3;
  wire f_u_arrmul12_fa1_4_y4;
  wire f_u_arrmul12_and2_4_a_2;
  wire f_u_arrmul12_and2_4_b_4;
  wire f_u_arrmul12_and2_4_y0;
  wire f_u_arrmul12_fa2_4_f_u_arrmul12_and2_4_y0;
  wire f_u_arrmul12_fa2_4_f_u_arrmul12_fa3_3_y2;
  wire f_u_arrmul12_fa2_4_y0;
  wire f_u_arrmul12_fa2_4_y1;
  wire f_u_arrmul12_fa2_4_f_u_arrmul12_fa1_4_y4;
  wire f_u_arrmul12_fa2_4_y2;
  wire f_u_arrmul12_fa2_4_y3;
  wire f_u_arrmul12_fa2_4_y4;
  wire f_u_arrmul12_and3_4_a_3;
  wire f_u_arrmul12_and3_4_b_4;
  wire f_u_arrmul12_and3_4_y0;
  wire f_u_arrmul12_fa3_4_f_u_arrmul12_and3_4_y0;
  wire f_u_arrmul12_fa3_4_f_u_arrmul12_fa4_3_y2;
  wire f_u_arrmul12_fa3_4_y0;
  wire f_u_arrmul12_fa3_4_y1;
  wire f_u_arrmul12_fa3_4_f_u_arrmul12_fa2_4_y4;
  wire f_u_arrmul12_fa3_4_y2;
  wire f_u_arrmul12_fa3_4_y3;
  wire f_u_arrmul12_fa3_4_y4;
  wire f_u_arrmul12_and4_4_a_4;
  wire f_u_arrmul12_and4_4_b_4;
  wire f_u_arrmul12_and4_4_y0;
  wire f_u_arrmul12_fa4_4_f_u_arrmul12_and4_4_y0;
  wire f_u_arrmul12_fa4_4_f_u_arrmul12_fa5_3_y2;
  wire f_u_arrmul12_fa4_4_y0;
  wire f_u_arrmul12_fa4_4_y1;
  wire f_u_arrmul12_fa4_4_f_u_arrmul12_fa3_4_y4;
  wire f_u_arrmul12_fa4_4_y2;
  wire f_u_arrmul12_fa4_4_y3;
  wire f_u_arrmul12_fa4_4_y4;
  wire f_u_arrmul12_and5_4_a_5;
  wire f_u_arrmul12_and5_4_b_4;
  wire f_u_arrmul12_and5_4_y0;
  wire f_u_arrmul12_fa5_4_f_u_arrmul12_and5_4_y0;
  wire f_u_arrmul12_fa5_4_f_u_arrmul12_fa6_3_y2;
  wire f_u_arrmul12_fa5_4_y0;
  wire f_u_arrmul12_fa5_4_y1;
  wire f_u_arrmul12_fa5_4_f_u_arrmul12_fa4_4_y4;
  wire f_u_arrmul12_fa5_4_y2;
  wire f_u_arrmul12_fa5_4_y3;
  wire f_u_arrmul12_fa5_4_y4;
  wire f_u_arrmul12_and6_4_a_6;
  wire f_u_arrmul12_and6_4_b_4;
  wire f_u_arrmul12_and6_4_y0;
  wire f_u_arrmul12_fa6_4_f_u_arrmul12_and6_4_y0;
  wire f_u_arrmul12_fa6_4_f_u_arrmul12_fa7_3_y2;
  wire f_u_arrmul12_fa6_4_y0;
  wire f_u_arrmul12_fa6_4_y1;
  wire f_u_arrmul12_fa6_4_f_u_arrmul12_fa5_4_y4;
  wire f_u_arrmul12_fa6_4_y2;
  wire f_u_arrmul12_fa6_4_y3;
  wire f_u_arrmul12_fa6_4_y4;
  wire f_u_arrmul12_and7_4_a_7;
  wire f_u_arrmul12_and7_4_b_4;
  wire f_u_arrmul12_and7_4_y0;
  wire f_u_arrmul12_fa7_4_f_u_arrmul12_and7_4_y0;
  wire f_u_arrmul12_fa7_4_f_u_arrmul12_fa8_3_y2;
  wire f_u_arrmul12_fa7_4_y0;
  wire f_u_arrmul12_fa7_4_y1;
  wire f_u_arrmul12_fa7_4_f_u_arrmul12_fa6_4_y4;
  wire f_u_arrmul12_fa7_4_y2;
  wire f_u_arrmul12_fa7_4_y3;
  wire f_u_arrmul12_fa7_4_y4;
  wire f_u_arrmul12_and8_4_a_8;
  wire f_u_arrmul12_and8_4_b_4;
  wire f_u_arrmul12_and8_4_y0;
  wire f_u_arrmul12_fa8_4_f_u_arrmul12_and8_4_y0;
  wire f_u_arrmul12_fa8_4_f_u_arrmul12_fa9_3_y2;
  wire f_u_arrmul12_fa8_4_y0;
  wire f_u_arrmul12_fa8_4_y1;
  wire f_u_arrmul12_fa8_4_f_u_arrmul12_fa7_4_y4;
  wire f_u_arrmul12_fa8_4_y2;
  wire f_u_arrmul12_fa8_4_y3;
  wire f_u_arrmul12_fa8_4_y4;
  wire f_u_arrmul12_and9_4_a_9;
  wire f_u_arrmul12_and9_4_b_4;
  wire f_u_arrmul12_and9_4_y0;
  wire f_u_arrmul12_fa9_4_f_u_arrmul12_and9_4_y0;
  wire f_u_arrmul12_fa9_4_f_u_arrmul12_fa10_3_y2;
  wire f_u_arrmul12_fa9_4_y0;
  wire f_u_arrmul12_fa9_4_y1;
  wire f_u_arrmul12_fa9_4_f_u_arrmul12_fa8_4_y4;
  wire f_u_arrmul12_fa9_4_y2;
  wire f_u_arrmul12_fa9_4_y3;
  wire f_u_arrmul12_fa9_4_y4;
  wire f_u_arrmul12_and10_4_a_10;
  wire f_u_arrmul12_and10_4_b_4;
  wire f_u_arrmul12_and10_4_y0;
  wire f_u_arrmul12_fa10_4_f_u_arrmul12_and10_4_y0;
  wire f_u_arrmul12_fa10_4_f_u_arrmul12_fa11_3_y2;
  wire f_u_arrmul12_fa10_4_y0;
  wire f_u_arrmul12_fa10_4_y1;
  wire f_u_arrmul12_fa10_4_f_u_arrmul12_fa9_4_y4;
  wire f_u_arrmul12_fa10_4_y2;
  wire f_u_arrmul12_fa10_4_y3;
  wire f_u_arrmul12_fa10_4_y4;
  wire f_u_arrmul12_and11_4_a_11;
  wire f_u_arrmul12_and11_4_b_4;
  wire f_u_arrmul12_and11_4_y0;
  wire f_u_arrmul12_fa11_4_f_u_arrmul12_and11_4_y0;
  wire f_u_arrmul12_fa11_4_f_u_arrmul12_fa11_3_y4;
  wire f_u_arrmul12_fa11_4_y0;
  wire f_u_arrmul12_fa11_4_y1;
  wire f_u_arrmul12_fa11_4_f_u_arrmul12_fa10_4_y4;
  wire f_u_arrmul12_fa11_4_y2;
  wire f_u_arrmul12_fa11_4_y3;
  wire f_u_arrmul12_fa11_4_y4;
  wire f_u_arrmul12_and0_5_a_0;
  wire f_u_arrmul12_and0_5_b_5;
  wire f_u_arrmul12_and0_5_y0;
  wire f_u_arrmul12_ha0_5_f_u_arrmul12_and0_5_y0;
  wire f_u_arrmul12_ha0_5_f_u_arrmul12_fa1_4_y2;
  wire f_u_arrmul12_ha0_5_y0;
  wire f_u_arrmul12_ha0_5_y1;
  wire f_u_arrmul12_and1_5_a_1;
  wire f_u_arrmul12_and1_5_b_5;
  wire f_u_arrmul12_and1_5_y0;
  wire f_u_arrmul12_fa1_5_f_u_arrmul12_and1_5_y0;
  wire f_u_arrmul12_fa1_5_f_u_arrmul12_fa2_4_y2;
  wire f_u_arrmul12_fa1_5_y0;
  wire f_u_arrmul12_fa1_5_y1;
  wire f_u_arrmul12_fa1_5_f_u_arrmul12_ha0_5_y1;
  wire f_u_arrmul12_fa1_5_y2;
  wire f_u_arrmul12_fa1_5_y3;
  wire f_u_arrmul12_fa1_5_y4;
  wire f_u_arrmul12_and2_5_a_2;
  wire f_u_arrmul12_and2_5_b_5;
  wire f_u_arrmul12_and2_5_y0;
  wire f_u_arrmul12_fa2_5_f_u_arrmul12_and2_5_y0;
  wire f_u_arrmul12_fa2_5_f_u_arrmul12_fa3_4_y2;
  wire f_u_arrmul12_fa2_5_y0;
  wire f_u_arrmul12_fa2_5_y1;
  wire f_u_arrmul12_fa2_5_f_u_arrmul12_fa1_5_y4;
  wire f_u_arrmul12_fa2_5_y2;
  wire f_u_arrmul12_fa2_5_y3;
  wire f_u_arrmul12_fa2_5_y4;
  wire f_u_arrmul12_and3_5_a_3;
  wire f_u_arrmul12_and3_5_b_5;
  wire f_u_arrmul12_and3_5_y0;
  wire f_u_arrmul12_fa3_5_f_u_arrmul12_and3_5_y0;
  wire f_u_arrmul12_fa3_5_f_u_arrmul12_fa4_4_y2;
  wire f_u_arrmul12_fa3_5_y0;
  wire f_u_arrmul12_fa3_5_y1;
  wire f_u_arrmul12_fa3_5_f_u_arrmul12_fa2_5_y4;
  wire f_u_arrmul12_fa3_5_y2;
  wire f_u_arrmul12_fa3_5_y3;
  wire f_u_arrmul12_fa3_5_y4;
  wire f_u_arrmul12_and4_5_a_4;
  wire f_u_arrmul12_and4_5_b_5;
  wire f_u_arrmul12_and4_5_y0;
  wire f_u_arrmul12_fa4_5_f_u_arrmul12_and4_5_y0;
  wire f_u_arrmul12_fa4_5_f_u_arrmul12_fa5_4_y2;
  wire f_u_arrmul12_fa4_5_y0;
  wire f_u_arrmul12_fa4_5_y1;
  wire f_u_arrmul12_fa4_5_f_u_arrmul12_fa3_5_y4;
  wire f_u_arrmul12_fa4_5_y2;
  wire f_u_arrmul12_fa4_5_y3;
  wire f_u_arrmul12_fa4_5_y4;
  wire f_u_arrmul12_and5_5_a_5;
  wire f_u_arrmul12_and5_5_b_5;
  wire f_u_arrmul12_and5_5_y0;
  wire f_u_arrmul12_fa5_5_f_u_arrmul12_and5_5_y0;
  wire f_u_arrmul12_fa5_5_f_u_arrmul12_fa6_4_y2;
  wire f_u_arrmul12_fa5_5_y0;
  wire f_u_arrmul12_fa5_5_y1;
  wire f_u_arrmul12_fa5_5_f_u_arrmul12_fa4_5_y4;
  wire f_u_arrmul12_fa5_5_y2;
  wire f_u_arrmul12_fa5_5_y3;
  wire f_u_arrmul12_fa5_5_y4;
  wire f_u_arrmul12_and6_5_a_6;
  wire f_u_arrmul12_and6_5_b_5;
  wire f_u_arrmul12_and6_5_y0;
  wire f_u_arrmul12_fa6_5_f_u_arrmul12_and6_5_y0;
  wire f_u_arrmul12_fa6_5_f_u_arrmul12_fa7_4_y2;
  wire f_u_arrmul12_fa6_5_y0;
  wire f_u_arrmul12_fa6_5_y1;
  wire f_u_arrmul12_fa6_5_f_u_arrmul12_fa5_5_y4;
  wire f_u_arrmul12_fa6_5_y2;
  wire f_u_arrmul12_fa6_5_y3;
  wire f_u_arrmul12_fa6_5_y4;
  wire f_u_arrmul12_and7_5_a_7;
  wire f_u_arrmul12_and7_5_b_5;
  wire f_u_arrmul12_and7_5_y0;
  wire f_u_arrmul12_fa7_5_f_u_arrmul12_and7_5_y0;
  wire f_u_arrmul12_fa7_5_f_u_arrmul12_fa8_4_y2;
  wire f_u_arrmul12_fa7_5_y0;
  wire f_u_arrmul12_fa7_5_y1;
  wire f_u_arrmul12_fa7_5_f_u_arrmul12_fa6_5_y4;
  wire f_u_arrmul12_fa7_5_y2;
  wire f_u_arrmul12_fa7_5_y3;
  wire f_u_arrmul12_fa7_5_y4;
  wire f_u_arrmul12_and8_5_a_8;
  wire f_u_arrmul12_and8_5_b_5;
  wire f_u_arrmul12_and8_5_y0;
  wire f_u_arrmul12_fa8_5_f_u_arrmul12_and8_5_y0;
  wire f_u_arrmul12_fa8_5_f_u_arrmul12_fa9_4_y2;
  wire f_u_arrmul12_fa8_5_y0;
  wire f_u_arrmul12_fa8_5_y1;
  wire f_u_arrmul12_fa8_5_f_u_arrmul12_fa7_5_y4;
  wire f_u_arrmul12_fa8_5_y2;
  wire f_u_arrmul12_fa8_5_y3;
  wire f_u_arrmul12_fa8_5_y4;
  wire f_u_arrmul12_and9_5_a_9;
  wire f_u_arrmul12_and9_5_b_5;
  wire f_u_arrmul12_and9_5_y0;
  wire f_u_arrmul12_fa9_5_f_u_arrmul12_and9_5_y0;
  wire f_u_arrmul12_fa9_5_f_u_arrmul12_fa10_4_y2;
  wire f_u_arrmul12_fa9_5_y0;
  wire f_u_arrmul12_fa9_5_y1;
  wire f_u_arrmul12_fa9_5_f_u_arrmul12_fa8_5_y4;
  wire f_u_arrmul12_fa9_5_y2;
  wire f_u_arrmul12_fa9_5_y3;
  wire f_u_arrmul12_fa9_5_y4;
  wire f_u_arrmul12_and10_5_a_10;
  wire f_u_arrmul12_and10_5_b_5;
  wire f_u_arrmul12_and10_5_y0;
  wire f_u_arrmul12_fa10_5_f_u_arrmul12_and10_5_y0;
  wire f_u_arrmul12_fa10_5_f_u_arrmul12_fa11_4_y2;
  wire f_u_arrmul12_fa10_5_y0;
  wire f_u_arrmul12_fa10_5_y1;
  wire f_u_arrmul12_fa10_5_f_u_arrmul12_fa9_5_y4;
  wire f_u_arrmul12_fa10_5_y2;
  wire f_u_arrmul12_fa10_5_y3;
  wire f_u_arrmul12_fa10_5_y4;
  wire f_u_arrmul12_and11_5_a_11;
  wire f_u_arrmul12_and11_5_b_5;
  wire f_u_arrmul12_and11_5_y0;
  wire f_u_arrmul12_fa11_5_f_u_arrmul12_and11_5_y0;
  wire f_u_arrmul12_fa11_5_f_u_arrmul12_fa11_4_y4;
  wire f_u_arrmul12_fa11_5_y0;
  wire f_u_arrmul12_fa11_5_y1;
  wire f_u_arrmul12_fa11_5_f_u_arrmul12_fa10_5_y4;
  wire f_u_arrmul12_fa11_5_y2;
  wire f_u_arrmul12_fa11_5_y3;
  wire f_u_arrmul12_fa11_5_y4;
  wire f_u_arrmul12_and0_6_a_0;
  wire f_u_arrmul12_and0_6_b_6;
  wire f_u_arrmul12_and0_6_y0;
  wire f_u_arrmul12_ha0_6_f_u_arrmul12_and0_6_y0;
  wire f_u_arrmul12_ha0_6_f_u_arrmul12_fa1_5_y2;
  wire f_u_arrmul12_ha0_6_y0;
  wire f_u_arrmul12_ha0_6_y1;
  wire f_u_arrmul12_and1_6_a_1;
  wire f_u_arrmul12_and1_6_b_6;
  wire f_u_arrmul12_and1_6_y0;
  wire f_u_arrmul12_fa1_6_f_u_arrmul12_and1_6_y0;
  wire f_u_arrmul12_fa1_6_f_u_arrmul12_fa2_5_y2;
  wire f_u_arrmul12_fa1_6_y0;
  wire f_u_arrmul12_fa1_6_y1;
  wire f_u_arrmul12_fa1_6_f_u_arrmul12_ha0_6_y1;
  wire f_u_arrmul12_fa1_6_y2;
  wire f_u_arrmul12_fa1_6_y3;
  wire f_u_arrmul12_fa1_6_y4;
  wire f_u_arrmul12_and2_6_a_2;
  wire f_u_arrmul12_and2_6_b_6;
  wire f_u_arrmul12_and2_6_y0;
  wire f_u_arrmul12_fa2_6_f_u_arrmul12_and2_6_y0;
  wire f_u_arrmul12_fa2_6_f_u_arrmul12_fa3_5_y2;
  wire f_u_arrmul12_fa2_6_y0;
  wire f_u_arrmul12_fa2_6_y1;
  wire f_u_arrmul12_fa2_6_f_u_arrmul12_fa1_6_y4;
  wire f_u_arrmul12_fa2_6_y2;
  wire f_u_arrmul12_fa2_6_y3;
  wire f_u_arrmul12_fa2_6_y4;
  wire f_u_arrmul12_and3_6_a_3;
  wire f_u_arrmul12_and3_6_b_6;
  wire f_u_arrmul12_and3_6_y0;
  wire f_u_arrmul12_fa3_6_f_u_arrmul12_and3_6_y0;
  wire f_u_arrmul12_fa3_6_f_u_arrmul12_fa4_5_y2;
  wire f_u_arrmul12_fa3_6_y0;
  wire f_u_arrmul12_fa3_6_y1;
  wire f_u_arrmul12_fa3_6_f_u_arrmul12_fa2_6_y4;
  wire f_u_arrmul12_fa3_6_y2;
  wire f_u_arrmul12_fa3_6_y3;
  wire f_u_arrmul12_fa3_6_y4;
  wire f_u_arrmul12_and4_6_a_4;
  wire f_u_arrmul12_and4_6_b_6;
  wire f_u_arrmul12_and4_6_y0;
  wire f_u_arrmul12_fa4_6_f_u_arrmul12_and4_6_y0;
  wire f_u_arrmul12_fa4_6_f_u_arrmul12_fa5_5_y2;
  wire f_u_arrmul12_fa4_6_y0;
  wire f_u_arrmul12_fa4_6_y1;
  wire f_u_arrmul12_fa4_6_f_u_arrmul12_fa3_6_y4;
  wire f_u_arrmul12_fa4_6_y2;
  wire f_u_arrmul12_fa4_6_y3;
  wire f_u_arrmul12_fa4_6_y4;
  wire f_u_arrmul12_and5_6_a_5;
  wire f_u_arrmul12_and5_6_b_6;
  wire f_u_arrmul12_and5_6_y0;
  wire f_u_arrmul12_fa5_6_f_u_arrmul12_and5_6_y0;
  wire f_u_arrmul12_fa5_6_f_u_arrmul12_fa6_5_y2;
  wire f_u_arrmul12_fa5_6_y0;
  wire f_u_arrmul12_fa5_6_y1;
  wire f_u_arrmul12_fa5_6_f_u_arrmul12_fa4_6_y4;
  wire f_u_arrmul12_fa5_6_y2;
  wire f_u_arrmul12_fa5_6_y3;
  wire f_u_arrmul12_fa5_6_y4;
  wire f_u_arrmul12_and6_6_a_6;
  wire f_u_arrmul12_and6_6_b_6;
  wire f_u_arrmul12_and6_6_y0;
  wire f_u_arrmul12_fa6_6_f_u_arrmul12_and6_6_y0;
  wire f_u_arrmul12_fa6_6_f_u_arrmul12_fa7_5_y2;
  wire f_u_arrmul12_fa6_6_y0;
  wire f_u_arrmul12_fa6_6_y1;
  wire f_u_arrmul12_fa6_6_f_u_arrmul12_fa5_6_y4;
  wire f_u_arrmul12_fa6_6_y2;
  wire f_u_arrmul12_fa6_6_y3;
  wire f_u_arrmul12_fa6_6_y4;
  wire f_u_arrmul12_and7_6_a_7;
  wire f_u_arrmul12_and7_6_b_6;
  wire f_u_arrmul12_and7_6_y0;
  wire f_u_arrmul12_fa7_6_f_u_arrmul12_and7_6_y0;
  wire f_u_arrmul12_fa7_6_f_u_arrmul12_fa8_5_y2;
  wire f_u_arrmul12_fa7_6_y0;
  wire f_u_arrmul12_fa7_6_y1;
  wire f_u_arrmul12_fa7_6_f_u_arrmul12_fa6_6_y4;
  wire f_u_arrmul12_fa7_6_y2;
  wire f_u_arrmul12_fa7_6_y3;
  wire f_u_arrmul12_fa7_6_y4;
  wire f_u_arrmul12_and8_6_a_8;
  wire f_u_arrmul12_and8_6_b_6;
  wire f_u_arrmul12_and8_6_y0;
  wire f_u_arrmul12_fa8_6_f_u_arrmul12_and8_6_y0;
  wire f_u_arrmul12_fa8_6_f_u_arrmul12_fa9_5_y2;
  wire f_u_arrmul12_fa8_6_y0;
  wire f_u_arrmul12_fa8_6_y1;
  wire f_u_arrmul12_fa8_6_f_u_arrmul12_fa7_6_y4;
  wire f_u_arrmul12_fa8_6_y2;
  wire f_u_arrmul12_fa8_6_y3;
  wire f_u_arrmul12_fa8_6_y4;
  wire f_u_arrmul12_and9_6_a_9;
  wire f_u_arrmul12_and9_6_b_6;
  wire f_u_arrmul12_and9_6_y0;
  wire f_u_arrmul12_fa9_6_f_u_arrmul12_and9_6_y0;
  wire f_u_arrmul12_fa9_6_f_u_arrmul12_fa10_5_y2;
  wire f_u_arrmul12_fa9_6_y0;
  wire f_u_arrmul12_fa9_6_y1;
  wire f_u_arrmul12_fa9_6_f_u_arrmul12_fa8_6_y4;
  wire f_u_arrmul12_fa9_6_y2;
  wire f_u_arrmul12_fa9_6_y3;
  wire f_u_arrmul12_fa9_6_y4;
  wire f_u_arrmul12_and10_6_a_10;
  wire f_u_arrmul12_and10_6_b_6;
  wire f_u_arrmul12_and10_6_y0;
  wire f_u_arrmul12_fa10_6_f_u_arrmul12_and10_6_y0;
  wire f_u_arrmul12_fa10_6_f_u_arrmul12_fa11_5_y2;
  wire f_u_arrmul12_fa10_6_y0;
  wire f_u_arrmul12_fa10_6_y1;
  wire f_u_arrmul12_fa10_6_f_u_arrmul12_fa9_6_y4;
  wire f_u_arrmul12_fa10_6_y2;
  wire f_u_arrmul12_fa10_6_y3;
  wire f_u_arrmul12_fa10_6_y4;
  wire f_u_arrmul12_and11_6_a_11;
  wire f_u_arrmul12_and11_6_b_6;
  wire f_u_arrmul12_and11_6_y0;
  wire f_u_arrmul12_fa11_6_f_u_arrmul12_and11_6_y0;
  wire f_u_arrmul12_fa11_6_f_u_arrmul12_fa11_5_y4;
  wire f_u_arrmul12_fa11_6_y0;
  wire f_u_arrmul12_fa11_6_y1;
  wire f_u_arrmul12_fa11_6_f_u_arrmul12_fa10_6_y4;
  wire f_u_arrmul12_fa11_6_y2;
  wire f_u_arrmul12_fa11_6_y3;
  wire f_u_arrmul12_fa11_6_y4;
  wire f_u_arrmul12_and0_7_a_0;
  wire f_u_arrmul12_and0_7_b_7;
  wire f_u_arrmul12_and0_7_y0;
  wire f_u_arrmul12_ha0_7_f_u_arrmul12_and0_7_y0;
  wire f_u_arrmul12_ha0_7_f_u_arrmul12_fa1_6_y2;
  wire f_u_arrmul12_ha0_7_y0;
  wire f_u_arrmul12_ha0_7_y1;
  wire f_u_arrmul12_and1_7_a_1;
  wire f_u_arrmul12_and1_7_b_7;
  wire f_u_arrmul12_and1_7_y0;
  wire f_u_arrmul12_fa1_7_f_u_arrmul12_and1_7_y0;
  wire f_u_arrmul12_fa1_7_f_u_arrmul12_fa2_6_y2;
  wire f_u_arrmul12_fa1_7_y0;
  wire f_u_arrmul12_fa1_7_y1;
  wire f_u_arrmul12_fa1_7_f_u_arrmul12_ha0_7_y1;
  wire f_u_arrmul12_fa1_7_y2;
  wire f_u_arrmul12_fa1_7_y3;
  wire f_u_arrmul12_fa1_7_y4;
  wire f_u_arrmul12_and2_7_a_2;
  wire f_u_arrmul12_and2_7_b_7;
  wire f_u_arrmul12_and2_7_y0;
  wire f_u_arrmul12_fa2_7_f_u_arrmul12_and2_7_y0;
  wire f_u_arrmul12_fa2_7_f_u_arrmul12_fa3_6_y2;
  wire f_u_arrmul12_fa2_7_y0;
  wire f_u_arrmul12_fa2_7_y1;
  wire f_u_arrmul12_fa2_7_f_u_arrmul12_fa1_7_y4;
  wire f_u_arrmul12_fa2_7_y2;
  wire f_u_arrmul12_fa2_7_y3;
  wire f_u_arrmul12_fa2_7_y4;
  wire f_u_arrmul12_and3_7_a_3;
  wire f_u_arrmul12_and3_7_b_7;
  wire f_u_arrmul12_and3_7_y0;
  wire f_u_arrmul12_fa3_7_f_u_arrmul12_and3_7_y0;
  wire f_u_arrmul12_fa3_7_f_u_arrmul12_fa4_6_y2;
  wire f_u_arrmul12_fa3_7_y0;
  wire f_u_arrmul12_fa3_7_y1;
  wire f_u_arrmul12_fa3_7_f_u_arrmul12_fa2_7_y4;
  wire f_u_arrmul12_fa3_7_y2;
  wire f_u_arrmul12_fa3_7_y3;
  wire f_u_arrmul12_fa3_7_y4;
  wire f_u_arrmul12_and4_7_a_4;
  wire f_u_arrmul12_and4_7_b_7;
  wire f_u_arrmul12_and4_7_y0;
  wire f_u_arrmul12_fa4_7_f_u_arrmul12_and4_7_y0;
  wire f_u_arrmul12_fa4_7_f_u_arrmul12_fa5_6_y2;
  wire f_u_arrmul12_fa4_7_y0;
  wire f_u_arrmul12_fa4_7_y1;
  wire f_u_arrmul12_fa4_7_f_u_arrmul12_fa3_7_y4;
  wire f_u_arrmul12_fa4_7_y2;
  wire f_u_arrmul12_fa4_7_y3;
  wire f_u_arrmul12_fa4_7_y4;
  wire f_u_arrmul12_and5_7_a_5;
  wire f_u_arrmul12_and5_7_b_7;
  wire f_u_arrmul12_and5_7_y0;
  wire f_u_arrmul12_fa5_7_f_u_arrmul12_and5_7_y0;
  wire f_u_arrmul12_fa5_7_f_u_arrmul12_fa6_6_y2;
  wire f_u_arrmul12_fa5_7_y0;
  wire f_u_arrmul12_fa5_7_y1;
  wire f_u_arrmul12_fa5_7_f_u_arrmul12_fa4_7_y4;
  wire f_u_arrmul12_fa5_7_y2;
  wire f_u_arrmul12_fa5_7_y3;
  wire f_u_arrmul12_fa5_7_y4;
  wire f_u_arrmul12_and6_7_a_6;
  wire f_u_arrmul12_and6_7_b_7;
  wire f_u_arrmul12_and6_7_y0;
  wire f_u_arrmul12_fa6_7_f_u_arrmul12_and6_7_y0;
  wire f_u_arrmul12_fa6_7_f_u_arrmul12_fa7_6_y2;
  wire f_u_arrmul12_fa6_7_y0;
  wire f_u_arrmul12_fa6_7_y1;
  wire f_u_arrmul12_fa6_7_f_u_arrmul12_fa5_7_y4;
  wire f_u_arrmul12_fa6_7_y2;
  wire f_u_arrmul12_fa6_7_y3;
  wire f_u_arrmul12_fa6_7_y4;
  wire f_u_arrmul12_and7_7_a_7;
  wire f_u_arrmul12_and7_7_b_7;
  wire f_u_arrmul12_and7_7_y0;
  wire f_u_arrmul12_fa7_7_f_u_arrmul12_and7_7_y0;
  wire f_u_arrmul12_fa7_7_f_u_arrmul12_fa8_6_y2;
  wire f_u_arrmul12_fa7_7_y0;
  wire f_u_arrmul12_fa7_7_y1;
  wire f_u_arrmul12_fa7_7_f_u_arrmul12_fa6_7_y4;
  wire f_u_arrmul12_fa7_7_y2;
  wire f_u_arrmul12_fa7_7_y3;
  wire f_u_arrmul12_fa7_7_y4;
  wire f_u_arrmul12_and8_7_a_8;
  wire f_u_arrmul12_and8_7_b_7;
  wire f_u_arrmul12_and8_7_y0;
  wire f_u_arrmul12_fa8_7_f_u_arrmul12_and8_7_y0;
  wire f_u_arrmul12_fa8_7_f_u_arrmul12_fa9_6_y2;
  wire f_u_arrmul12_fa8_7_y0;
  wire f_u_arrmul12_fa8_7_y1;
  wire f_u_arrmul12_fa8_7_f_u_arrmul12_fa7_7_y4;
  wire f_u_arrmul12_fa8_7_y2;
  wire f_u_arrmul12_fa8_7_y3;
  wire f_u_arrmul12_fa8_7_y4;
  wire f_u_arrmul12_and9_7_a_9;
  wire f_u_arrmul12_and9_7_b_7;
  wire f_u_arrmul12_and9_7_y0;
  wire f_u_arrmul12_fa9_7_f_u_arrmul12_and9_7_y0;
  wire f_u_arrmul12_fa9_7_f_u_arrmul12_fa10_6_y2;
  wire f_u_arrmul12_fa9_7_y0;
  wire f_u_arrmul12_fa9_7_y1;
  wire f_u_arrmul12_fa9_7_f_u_arrmul12_fa8_7_y4;
  wire f_u_arrmul12_fa9_7_y2;
  wire f_u_arrmul12_fa9_7_y3;
  wire f_u_arrmul12_fa9_7_y4;
  wire f_u_arrmul12_and10_7_a_10;
  wire f_u_arrmul12_and10_7_b_7;
  wire f_u_arrmul12_and10_7_y0;
  wire f_u_arrmul12_fa10_7_f_u_arrmul12_and10_7_y0;
  wire f_u_arrmul12_fa10_7_f_u_arrmul12_fa11_6_y2;
  wire f_u_arrmul12_fa10_7_y0;
  wire f_u_arrmul12_fa10_7_y1;
  wire f_u_arrmul12_fa10_7_f_u_arrmul12_fa9_7_y4;
  wire f_u_arrmul12_fa10_7_y2;
  wire f_u_arrmul12_fa10_7_y3;
  wire f_u_arrmul12_fa10_7_y4;
  wire f_u_arrmul12_and11_7_a_11;
  wire f_u_arrmul12_and11_7_b_7;
  wire f_u_arrmul12_and11_7_y0;
  wire f_u_arrmul12_fa11_7_f_u_arrmul12_and11_7_y0;
  wire f_u_arrmul12_fa11_7_f_u_arrmul12_fa11_6_y4;
  wire f_u_arrmul12_fa11_7_y0;
  wire f_u_arrmul12_fa11_7_y1;
  wire f_u_arrmul12_fa11_7_f_u_arrmul12_fa10_7_y4;
  wire f_u_arrmul12_fa11_7_y2;
  wire f_u_arrmul12_fa11_7_y3;
  wire f_u_arrmul12_fa11_7_y4;
  wire f_u_arrmul12_and0_8_a_0;
  wire f_u_arrmul12_and0_8_b_8;
  wire f_u_arrmul12_and0_8_y0;
  wire f_u_arrmul12_ha0_8_f_u_arrmul12_and0_8_y0;
  wire f_u_arrmul12_ha0_8_f_u_arrmul12_fa1_7_y2;
  wire f_u_arrmul12_ha0_8_y0;
  wire f_u_arrmul12_ha0_8_y1;
  wire f_u_arrmul12_and1_8_a_1;
  wire f_u_arrmul12_and1_8_b_8;
  wire f_u_arrmul12_and1_8_y0;
  wire f_u_arrmul12_fa1_8_f_u_arrmul12_and1_8_y0;
  wire f_u_arrmul12_fa1_8_f_u_arrmul12_fa2_7_y2;
  wire f_u_arrmul12_fa1_8_y0;
  wire f_u_arrmul12_fa1_8_y1;
  wire f_u_arrmul12_fa1_8_f_u_arrmul12_ha0_8_y1;
  wire f_u_arrmul12_fa1_8_y2;
  wire f_u_arrmul12_fa1_8_y3;
  wire f_u_arrmul12_fa1_8_y4;
  wire f_u_arrmul12_and2_8_a_2;
  wire f_u_arrmul12_and2_8_b_8;
  wire f_u_arrmul12_and2_8_y0;
  wire f_u_arrmul12_fa2_8_f_u_arrmul12_and2_8_y0;
  wire f_u_arrmul12_fa2_8_f_u_arrmul12_fa3_7_y2;
  wire f_u_arrmul12_fa2_8_y0;
  wire f_u_arrmul12_fa2_8_y1;
  wire f_u_arrmul12_fa2_8_f_u_arrmul12_fa1_8_y4;
  wire f_u_arrmul12_fa2_8_y2;
  wire f_u_arrmul12_fa2_8_y3;
  wire f_u_arrmul12_fa2_8_y4;
  wire f_u_arrmul12_and3_8_a_3;
  wire f_u_arrmul12_and3_8_b_8;
  wire f_u_arrmul12_and3_8_y0;
  wire f_u_arrmul12_fa3_8_f_u_arrmul12_and3_8_y0;
  wire f_u_arrmul12_fa3_8_f_u_arrmul12_fa4_7_y2;
  wire f_u_arrmul12_fa3_8_y0;
  wire f_u_arrmul12_fa3_8_y1;
  wire f_u_arrmul12_fa3_8_f_u_arrmul12_fa2_8_y4;
  wire f_u_arrmul12_fa3_8_y2;
  wire f_u_arrmul12_fa3_8_y3;
  wire f_u_arrmul12_fa3_8_y4;
  wire f_u_arrmul12_and4_8_a_4;
  wire f_u_arrmul12_and4_8_b_8;
  wire f_u_arrmul12_and4_8_y0;
  wire f_u_arrmul12_fa4_8_f_u_arrmul12_and4_8_y0;
  wire f_u_arrmul12_fa4_8_f_u_arrmul12_fa5_7_y2;
  wire f_u_arrmul12_fa4_8_y0;
  wire f_u_arrmul12_fa4_8_y1;
  wire f_u_arrmul12_fa4_8_f_u_arrmul12_fa3_8_y4;
  wire f_u_arrmul12_fa4_8_y2;
  wire f_u_arrmul12_fa4_8_y3;
  wire f_u_arrmul12_fa4_8_y4;
  wire f_u_arrmul12_and5_8_a_5;
  wire f_u_arrmul12_and5_8_b_8;
  wire f_u_arrmul12_and5_8_y0;
  wire f_u_arrmul12_fa5_8_f_u_arrmul12_and5_8_y0;
  wire f_u_arrmul12_fa5_8_f_u_arrmul12_fa6_7_y2;
  wire f_u_arrmul12_fa5_8_y0;
  wire f_u_arrmul12_fa5_8_y1;
  wire f_u_arrmul12_fa5_8_f_u_arrmul12_fa4_8_y4;
  wire f_u_arrmul12_fa5_8_y2;
  wire f_u_arrmul12_fa5_8_y3;
  wire f_u_arrmul12_fa5_8_y4;
  wire f_u_arrmul12_and6_8_a_6;
  wire f_u_arrmul12_and6_8_b_8;
  wire f_u_arrmul12_and6_8_y0;
  wire f_u_arrmul12_fa6_8_f_u_arrmul12_and6_8_y0;
  wire f_u_arrmul12_fa6_8_f_u_arrmul12_fa7_7_y2;
  wire f_u_arrmul12_fa6_8_y0;
  wire f_u_arrmul12_fa6_8_y1;
  wire f_u_arrmul12_fa6_8_f_u_arrmul12_fa5_8_y4;
  wire f_u_arrmul12_fa6_8_y2;
  wire f_u_arrmul12_fa6_8_y3;
  wire f_u_arrmul12_fa6_8_y4;
  wire f_u_arrmul12_and7_8_a_7;
  wire f_u_arrmul12_and7_8_b_8;
  wire f_u_arrmul12_and7_8_y0;
  wire f_u_arrmul12_fa7_8_f_u_arrmul12_and7_8_y0;
  wire f_u_arrmul12_fa7_8_f_u_arrmul12_fa8_7_y2;
  wire f_u_arrmul12_fa7_8_y0;
  wire f_u_arrmul12_fa7_8_y1;
  wire f_u_arrmul12_fa7_8_f_u_arrmul12_fa6_8_y4;
  wire f_u_arrmul12_fa7_8_y2;
  wire f_u_arrmul12_fa7_8_y3;
  wire f_u_arrmul12_fa7_8_y4;
  wire f_u_arrmul12_and8_8_a_8;
  wire f_u_arrmul12_and8_8_b_8;
  wire f_u_arrmul12_and8_8_y0;
  wire f_u_arrmul12_fa8_8_f_u_arrmul12_and8_8_y0;
  wire f_u_arrmul12_fa8_8_f_u_arrmul12_fa9_7_y2;
  wire f_u_arrmul12_fa8_8_y0;
  wire f_u_arrmul12_fa8_8_y1;
  wire f_u_arrmul12_fa8_8_f_u_arrmul12_fa7_8_y4;
  wire f_u_arrmul12_fa8_8_y2;
  wire f_u_arrmul12_fa8_8_y3;
  wire f_u_arrmul12_fa8_8_y4;
  wire f_u_arrmul12_and9_8_a_9;
  wire f_u_arrmul12_and9_8_b_8;
  wire f_u_arrmul12_and9_8_y0;
  wire f_u_arrmul12_fa9_8_f_u_arrmul12_and9_8_y0;
  wire f_u_arrmul12_fa9_8_f_u_arrmul12_fa10_7_y2;
  wire f_u_arrmul12_fa9_8_y0;
  wire f_u_arrmul12_fa9_8_y1;
  wire f_u_arrmul12_fa9_8_f_u_arrmul12_fa8_8_y4;
  wire f_u_arrmul12_fa9_8_y2;
  wire f_u_arrmul12_fa9_8_y3;
  wire f_u_arrmul12_fa9_8_y4;
  wire f_u_arrmul12_and10_8_a_10;
  wire f_u_arrmul12_and10_8_b_8;
  wire f_u_arrmul12_and10_8_y0;
  wire f_u_arrmul12_fa10_8_f_u_arrmul12_and10_8_y0;
  wire f_u_arrmul12_fa10_8_f_u_arrmul12_fa11_7_y2;
  wire f_u_arrmul12_fa10_8_y0;
  wire f_u_arrmul12_fa10_8_y1;
  wire f_u_arrmul12_fa10_8_f_u_arrmul12_fa9_8_y4;
  wire f_u_arrmul12_fa10_8_y2;
  wire f_u_arrmul12_fa10_8_y3;
  wire f_u_arrmul12_fa10_8_y4;
  wire f_u_arrmul12_and11_8_a_11;
  wire f_u_arrmul12_and11_8_b_8;
  wire f_u_arrmul12_and11_8_y0;
  wire f_u_arrmul12_fa11_8_f_u_arrmul12_and11_8_y0;
  wire f_u_arrmul12_fa11_8_f_u_arrmul12_fa11_7_y4;
  wire f_u_arrmul12_fa11_8_y0;
  wire f_u_arrmul12_fa11_8_y1;
  wire f_u_arrmul12_fa11_8_f_u_arrmul12_fa10_8_y4;
  wire f_u_arrmul12_fa11_8_y2;
  wire f_u_arrmul12_fa11_8_y3;
  wire f_u_arrmul12_fa11_8_y4;
  wire f_u_arrmul12_and0_9_a_0;
  wire f_u_arrmul12_and0_9_b_9;
  wire f_u_arrmul12_and0_9_y0;
  wire f_u_arrmul12_ha0_9_f_u_arrmul12_and0_9_y0;
  wire f_u_arrmul12_ha0_9_f_u_arrmul12_fa1_8_y2;
  wire f_u_arrmul12_ha0_9_y0;
  wire f_u_arrmul12_ha0_9_y1;
  wire f_u_arrmul12_and1_9_a_1;
  wire f_u_arrmul12_and1_9_b_9;
  wire f_u_arrmul12_and1_9_y0;
  wire f_u_arrmul12_fa1_9_f_u_arrmul12_and1_9_y0;
  wire f_u_arrmul12_fa1_9_f_u_arrmul12_fa2_8_y2;
  wire f_u_arrmul12_fa1_9_y0;
  wire f_u_arrmul12_fa1_9_y1;
  wire f_u_arrmul12_fa1_9_f_u_arrmul12_ha0_9_y1;
  wire f_u_arrmul12_fa1_9_y2;
  wire f_u_arrmul12_fa1_9_y3;
  wire f_u_arrmul12_fa1_9_y4;
  wire f_u_arrmul12_and2_9_a_2;
  wire f_u_arrmul12_and2_9_b_9;
  wire f_u_arrmul12_and2_9_y0;
  wire f_u_arrmul12_fa2_9_f_u_arrmul12_and2_9_y0;
  wire f_u_arrmul12_fa2_9_f_u_arrmul12_fa3_8_y2;
  wire f_u_arrmul12_fa2_9_y0;
  wire f_u_arrmul12_fa2_9_y1;
  wire f_u_arrmul12_fa2_9_f_u_arrmul12_fa1_9_y4;
  wire f_u_arrmul12_fa2_9_y2;
  wire f_u_arrmul12_fa2_9_y3;
  wire f_u_arrmul12_fa2_9_y4;
  wire f_u_arrmul12_and3_9_a_3;
  wire f_u_arrmul12_and3_9_b_9;
  wire f_u_arrmul12_and3_9_y0;
  wire f_u_arrmul12_fa3_9_f_u_arrmul12_and3_9_y0;
  wire f_u_arrmul12_fa3_9_f_u_arrmul12_fa4_8_y2;
  wire f_u_arrmul12_fa3_9_y0;
  wire f_u_arrmul12_fa3_9_y1;
  wire f_u_arrmul12_fa3_9_f_u_arrmul12_fa2_9_y4;
  wire f_u_arrmul12_fa3_9_y2;
  wire f_u_arrmul12_fa3_9_y3;
  wire f_u_arrmul12_fa3_9_y4;
  wire f_u_arrmul12_and4_9_a_4;
  wire f_u_arrmul12_and4_9_b_9;
  wire f_u_arrmul12_and4_9_y0;
  wire f_u_arrmul12_fa4_9_f_u_arrmul12_and4_9_y0;
  wire f_u_arrmul12_fa4_9_f_u_arrmul12_fa5_8_y2;
  wire f_u_arrmul12_fa4_9_y0;
  wire f_u_arrmul12_fa4_9_y1;
  wire f_u_arrmul12_fa4_9_f_u_arrmul12_fa3_9_y4;
  wire f_u_arrmul12_fa4_9_y2;
  wire f_u_arrmul12_fa4_9_y3;
  wire f_u_arrmul12_fa4_9_y4;
  wire f_u_arrmul12_and5_9_a_5;
  wire f_u_arrmul12_and5_9_b_9;
  wire f_u_arrmul12_and5_9_y0;
  wire f_u_arrmul12_fa5_9_f_u_arrmul12_and5_9_y0;
  wire f_u_arrmul12_fa5_9_f_u_arrmul12_fa6_8_y2;
  wire f_u_arrmul12_fa5_9_y0;
  wire f_u_arrmul12_fa5_9_y1;
  wire f_u_arrmul12_fa5_9_f_u_arrmul12_fa4_9_y4;
  wire f_u_arrmul12_fa5_9_y2;
  wire f_u_arrmul12_fa5_9_y3;
  wire f_u_arrmul12_fa5_9_y4;
  wire f_u_arrmul12_and6_9_a_6;
  wire f_u_arrmul12_and6_9_b_9;
  wire f_u_arrmul12_and6_9_y0;
  wire f_u_arrmul12_fa6_9_f_u_arrmul12_and6_9_y0;
  wire f_u_arrmul12_fa6_9_f_u_arrmul12_fa7_8_y2;
  wire f_u_arrmul12_fa6_9_y0;
  wire f_u_arrmul12_fa6_9_y1;
  wire f_u_arrmul12_fa6_9_f_u_arrmul12_fa5_9_y4;
  wire f_u_arrmul12_fa6_9_y2;
  wire f_u_arrmul12_fa6_9_y3;
  wire f_u_arrmul12_fa6_9_y4;
  wire f_u_arrmul12_and7_9_a_7;
  wire f_u_arrmul12_and7_9_b_9;
  wire f_u_arrmul12_and7_9_y0;
  wire f_u_arrmul12_fa7_9_f_u_arrmul12_and7_9_y0;
  wire f_u_arrmul12_fa7_9_f_u_arrmul12_fa8_8_y2;
  wire f_u_arrmul12_fa7_9_y0;
  wire f_u_arrmul12_fa7_9_y1;
  wire f_u_arrmul12_fa7_9_f_u_arrmul12_fa6_9_y4;
  wire f_u_arrmul12_fa7_9_y2;
  wire f_u_arrmul12_fa7_9_y3;
  wire f_u_arrmul12_fa7_9_y4;
  wire f_u_arrmul12_and8_9_a_8;
  wire f_u_arrmul12_and8_9_b_9;
  wire f_u_arrmul12_and8_9_y0;
  wire f_u_arrmul12_fa8_9_f_u_arrmul12_and8_9_y0;
  wire f_u_arrmul12_fa8_9_f_u_arrmul12_fa9_8_y2;
  wire f_u_arrmul12_fa8_9_y0;
  wire f_u_arrmul12_fa8_9_y1;
  wire f_u_arrmul12_fa8_9_f_u_arrmul12_fa7_9_y4;
  wire f_u_arrmul12_fa8_9_y2;
  wire f_u_arrmul12_fa8_9_y3;
  wire f_u_arrmul12_fa8_9_y4;
  wire f_u_arrmul12_and9_9_a_9;
  wire f_u_arrmul12_and9_9_b_9;
  wire f_u_arrmul12_and9_9_y0;
  wire f_u_arrmul12_fa9_9_f_u_arrmul12_and9_9_y0;
  wire f_u_arrmul12_fa9_9_f_u_arrmul12_fa10_8_y2;
  wire f_u_arrmul12_fa9_9_y0;
  wire f_u_arrmul12_fa9_9_y1;
  wire f_u_arrmul12_fa9_9_f_u_arrmul12_fa8_9_y4;
  wire f_u_arrmul12_fa9_9_y2;
  wire f_u_arrmul12_fa9_9_y3;
  wire f_u_arrmul12_fa9_9_y4;
  wire f_u_arrmul12_and10_9_a_10;
  wire f_u_arrmul12_and10_9_b_9;
  wire f_u_arrmul12_and10_9_y0;
  wire f_u_arrmul12_fa10_9_f_u_arrmul12_and10_9_y0;
  wire f_u_arrmul12_fa10_9_f_u_arrmul12_fa11_8_y2;
  wire f_u_arrmul12_fa10_9_y0;
  wire f_u_arrmul12_fa10_9_y1;
  wire f_u_arrmul12_fa10_9_f_u_arrmul12_fa9_9_y4;
  wire f_u_arrmul12_fa10_9_y2;
  wire f_u_arrmul12_fa10_9_y3;
  wire f_u_arrmul12_fa10_9_y4;
  wire f_u_arrmul12_and11_9_a_11;
  wire f_u_arrmul12_and11_9_b_9;
  wire f_u_arrmul12_and11_9_y0;
  wire f_u_arrmul12_fa11_9_f_u_arrmul12_and11_9_y0;
  wire f_u_arrmul12_fa11_9_f_u_arrmul12_fa11_8_y4;
  wire f_u_arrmul12_fa11_9_y0;
  wire f_u_arrmul12_fa11_9_y1;
  wire f_u_arrmul12_fa11_9_f_u_arrmul12_fa10_9_y4;
  wire f_u_arrmul12_fa11_9_y2;
  wire f_u_arrmul12_fa11_9_y3;
  wire f_u_arrmul12_fa11_9_y4;
  wire f_u_arrmul12_and0_10_a_0;
  wire f_u_arrmul12_and0_10_b_10;
  wire f_u_arrmul12_and0_10_y0;
  wire f_u_arrmul12_ha0_10_f_u_arrmul12_and0_10_y0;
  wire f_u_arrmul12_ha0_10_f_u_arrmul12_fa1_9_y2;
  wire f_u_arrmul12_ha0_10_y0;
  wire f_u_arrmul12_ha0_10_y1;
  wire f_u_arrmul12_and1_10_a_1;
  wire f_u_arrmul12_and1_10_b_10;
  wire f_u_arrmul12_and1_10_y0;
  wire f_u_arrmul12_fa1_10_f_u_arrmul12_and1_10_y0;
  wire f_u_arrmul12_fa1_10_f_u_arrmul12_fa2_9_y2;
  wire f_u_arrmul12_fa1_10_y0;
  wire f_u_arrmul12_fa1_10_y1;
  wire f_u_arrmul12_fa1_10_f_u_arrmul12_ha0_10_y1;
  wire f_u_arrmul12_fa1_10_y2;
  wire f_u_arrmul12_fa1_10_y3;
  wire f_u_arrmul12_fa1_10_y4;
  wire f_u_arrmul12_and2_10_a_2;
  wire f_u_arrmul12_and2_10_b_10;
  wire f_u_arrmul12_and2_10_y0;
  wire f_u_arrmul12_fa2_10_f_u_arrmul12_and2_10_y0;
  wire f_u_arrmul12_fa2_10_f_u_arrmul12_fa3_9_y2;
  wire f_u_arrmul12_fa2_10_y0;
  wire f_u_arrmul12_fa2_10_y1;
  wire f_u_arrmul12_fa2_10_f_u_arrmul12_fa1_10_y4;
  wire f_u_arrmul12_fa2_10_y2;
  wire f_u_arrmul12_fa2_10_y3;
  wire f_u_arrmul12_fa2_10_y4;
  wire f_u_arrmul12_and3_10_a_3;
  wire f_u_arrmul12_and3_10_b_10;
  wire f_u_arrmul12_and3_10_y0;
  wire f_u_arrmul12_fa3_10_f_u_arrmul12_and3_10_y0;
  wire f_u_arrmul12_fa3_10_f_u_arrmul12_fa4_9_y2;
  wire f_u_arrmul12_fa3_10_y0;
  wire f_u_arrmul12_fa3_10_y1;
  wire f_u_arrmul12_fa3_10_f_u_arrmul12_fa2_10_y4;
  wire f_u_arrmul12_fa3_10_y2;
  wire f_u_arrmul12_fa3_10_y3;
  wire f_u_arrmul12_fa3_10_y4;
  wire f_u_arrmul12_and4_10_a_4;
  wire f_u_arrmul12_and4_10_b_10;
  wire f_u_arrmul12_and4_10_y0;
  wire f_u_arrmul12_fa4_10_f_u_arrmul12_and4_10_y0;
  wire f_u_arrmul12_fa4_10_f_u_arrmul12_fa5_9_y2;
  wire f_u_arrmul12_fa4_10_y0;
  wire f_u_arrmul12_fa4_10_y1;
  wire f_u_arrmul12_fa4_10_f_u_arrmul12_fa3_10_y4;
  wire f_u_arrmul12_fa4_10_y2;
  wire f_u_arrmul12_fa4_10_y3;
  wire f_u_arrmul12_fa4_10_y4;
  wire f_u_arrmul12_and5_10_a_5;
  wire f_u_arrmul12_and5_10_b_10;
  wire f_u_arrmul12_and5_10_y0;
  wire f_u_arrmul12_fa5_10_f_u_arrmul12_and5_10_y0;
  wire f_u_arrmul12_fa5_10_f_u_arrmul12_fa6_9_y2;
  wire f_u_arrmul12_fa5_10_y0;
  wire f_u_arrmul12_fa5_10_y1;
  wire f_u_arrmul12_fa5_10_f_u_arrmul12_fa4_10_y4;
  wire f_u_arrmul12_fa5_10_y2;
  wire f_u_arrmul12_fa5_10_y3;
  wire f_u_arrmul12_fa5_10_y4;
  wire f_u_arrmul12_and6_10_a_6;
  wire f_u_arrmul12_and6_10_b_10;
  wire f_u_arrmul12_and6_10_y0;
  wire f_u_arrmul12_fa6_10_f_u_arrmul12_and6_10_y0;
  wire f_u_arrmul12_fa6_10_f_u_arrmul12_fa7_9_y2;
  wire f_u_arrmul12_fa6_10_y0;
  wire f_u_arrmul12_fa6_10_y1;
  wire f_u_arrmul12_fa6_10_f_u_arrmul12_fa5_10_y4;
  wire f_u_arrmul12_fa6_10_y2;
  wire f_u_arrmul12_fa6_10_y3;
  wire f_u_arrmul12_fa6_10_y4;
  wire f_u_arrmul12_and7_10_a_7;
  wire f_u_arrmul12_and7_10_b_10;
  wire f_u_arrmul12_and7_10_y0;
  wire f_u_arrmul12_fa7_10_f_u_arrmul12_and7_10_y0;
  wire f_u_arrmul12_fa7_10_f_u_arrmul12_fa8_9_y2;
  wire f_u_arrmul12_fa7_10_y0;
  wire f_u_arrmul12_fa7_10_y1;
  wire f_u_arrmul12_fa7_10_f_u_arrmul12_fa6_10_y4;
  wire f_u_arrmul12_fa7_10_y2;
  wire f_u_arrmul12_fa7_10_y3;
  wire f_u_arrmul12_fa7_10_y4;
  wire f_u_arrmul12_and8_10_a_8;
  wire f_u_arrmul12_and8_10_b_10;
  wire f_u_arrmul12_and8_10_y0;
  wire f_u_arrmul12_fa8_10_f_u_arrmul12_and8_10_y0;
  wire f_u_arrmul12_fa8_10_f_u_arrmul12_fa9_9_y2;
  wire f_u_arrmul12_fa8_10_y0;
  wire f_u_arrmul12_fa8_10_y1;
  wire f_u_arrmul12_fa8_10_f_u_arrmul12_fa7_10_y4;
  wire f_u_arrmul12_fa8_10_y2;
  wire f_u_arrmul12_fa8_10_y3;
  wire f_u_arrmul12_fa8_10_y4;
  wire f_u_arrmul12_and9_10_a_9;
  wire f_u_arrmul12_and9_10_b_10;
  wire f_u_arrmul12_and9_10_y0;
  wire f_u_arrmul12_fa9_10_f_u_arrmul12_and9_10_y0;
  wire f_u_arrmul12_fa9_10_f_u_arrmul12_fa10_9_y2;
  wire f_u_arrmul12_fa9_10_y0;
  wire f_u_arrmul12_fa9_10_y1;
  wire f_u_arrmul12_fa9_10_f_u_arrmul12_fa8_10_y4;
  wire f_u_arrmul12_fa9_10_y2;
  wire f_u_arrmul12_fa9_10_y3;
  wire f_u_arrmul12_fa9_10_y4;
  wire f_u_arrmul12_and10_10_a_10;
  wire f_u_arrmul12_and10_10_b_10;
  wire f_u_arrmul12_and10_10_y0;
  wire f_u_arrmul12_fa10_10_f_u_arrmul12_and10_10_y0;
  wire f_u_arrmul12_fa10_10_f_u_arrmul12_fa11_9_y2;
  wire f_u_arrmul12_fa10_10_y0;
  wire f_u_arrmul12_fa10_10_y1;
  wire f_u_arrmul12_fa10_10_f_u_arrmul12_fa9_10_y4;
  wire f_u_arrmul12_fa10_10_y2;
  wire f_u_arrmul12_fa10_10_y3;
  wire f_u_arrmul12_fa10_10_y4;
  wire f_u_arrmul12_and11_10_a_11;
  wire f_u_arrmul12_and11_10_b_10;
  wire f_u_arrmul12_and11_10_y0;
  wire f_u_arrmul12_fa11_10_f_u_arrmul12_and11_10_y0;
  wire f_u_arrmul12_fa11_10_f_u_arrmul12_fa11_9_y4;
  wire f_u_arrmul12_fa11_10_y0;
  wire f_u_arrmul12_fa11_10_y1;
  wire f_u_arrmul12_fa11_10_f_u_arrmul12_fa10_10_y4;
  wire f_u_arrmul12_fa11_10_y2;
  wire f_u_arrmul12_fa11_10_y3;
  wire f_u_arrmul12_fa11_10_y4;
  wire f_u_arrmul12_and0_11_a_0;
  wire f_u_arrmul12_and0_11_b_11;
  wire f_u_arrmul12_and0_11_y0;
  wire f_u_arrmul12_ha0_11_f_u_arrmul12_and0_11_y0;
  wire f_u_arrmul12_ha0_11_f_u_arrmul12_fa1_10_y2;
  wire f_u_arrmul12_ha0_11_y0;
  wire f_u_arrmul12_ha0_11_y1;
  wire f_u_arrmul12_and1_11_a_1;
  wire f_u_arrmul12_and1_11_b_11;
  wire f_u_arrmul12_and1_11_y0;
  wire f_u_arrmul12_fa1_11_f_u_arrmul12_and1_11_y0;
  wire f_u_arrmul12_fa1_11_f_u_arrmul12_fa2_10_y2;
  wire f_u_arrmul12_fa1_11_y0;
  wire f_u_arrmul12_fa1_11_y1;
  wire f_u_arrmul12_fa1_11_f_u_arrmul12_ha0_11_y1;
  wire f_u_arrmul12_fa1_11_y2;
  wire f_u_arrmul12_fa1_11_y3;
  wire f_u_arrmul12_fa1_11_y4;
  wire f_u_arrmul12_and2_11_a_2;
  wire f_u_arrmul12_and2_11_b_11;
  wire f_u_arrmul12_and2_11_y0;
  wire f_u_arrmul12_fa2_11_f_u_arrmul12_and2_11_y0;
  wire f_u_arrmul12_fa2_11_f_u_arrmul12_fa3_10_y2;
  wire f_u_arrmul12_fa2_11_y0;
  wire f_u_arrmul12_fa2_11_y1;
  wire f_u_arrmul12_fa2_11_f_u_arrmul12_fa1_11_y4;
  wire f_u_arrmul12_fa2_11_y2;
  wire f_u_arrmul12_fa2_11_y3;
  wire f_u_arrmul12_fa2_11_y4;
  wire f_u_arrmul12_and3_11_a_3;
  wire f_u_arrmul12_and3_11_b_11;
  wire f_u_arrmul12_and3_11_y0;
  wire f_u_arrmul12_fa3_11_f_u_arrmul12_and3_11_y0;
  wire f_u_arrmul12_fa3_11_f_u_arrmul12_fa4_10_y2;
  wire f_u_arrmul12_fa3_11_y0;
  wire f_u_arrmul12_fa3_11_y1;
  wire f_u_arrmul12_fa3_11_f_u_arrmul12_fa2_11_y4;
  wire f_u_arrmul12_fa3_11_y2;
  wire f_u_arrmul12_fa3_11_y3;
  wire f_u_arrmul12_fa3_11_y4;
  wire f_u_arrmul12_and4_11_a_4;
  wire f_u_arrmul12_and4_11_b_11;
  wire f_u_arrmul12_and4_11_y0;
  wire f_u_arrmul12_fa4_11_f_u_arrmul12_and4_11_y0;
  wire f_u_arrmul12_fa4_11_f_u_arrmul12_fa5_10_y2;
  wire f_u_arrmul12_fa4_11_y0;
  wire f_u_arrmul12_fa4_11_y1;
  wire f_u_arrmul12_fa4_11_f_u_arrmul12_fa3_11_y4;
  wire f_u_arrmul12_fa4_11_y2;
  wire f_u_arrmul12_fa4_11_y3;
  wire f_u_arrmul12_fa4_11_y4;
  wire f_u_arrmul12_and5_11_a_5;
  wire f_u_arrmul12_and5_11_b_11;
  wire f_u_arrmul12_and5_11_y0;
  wire f_u_arrmul12_fa5_11_f_u_arrmul12_and5_11_y0;
  wire f_u_arrmul12_fa5_11_f_u_arrmul12_fa6_10_y2;
  wire f_u_arrmul12_fa5_11_y0;
  wire f_u_arrmul12_fa5_11_y1;
  wire f_u_arrmul12_fa5_11_f_u_arrmul12_fa4_11_y4;
  wire f_u_arrmul12_fa5_11_y2;
  wire f_u_arrmul12_fa5_11_y3;
  wire f_u_arrmul12_fa5_11_y4;
  wire f_u_arrmul12_and6_11_a_6;
  wire f_u_arrmul12_and6_11_b_11;
  wire f_u_arrmul12_and6_11_y0;
  wire f_u_arrmul12_fa6_11_f_u_arrmul12_and6_11_y0;
  wire f_u_arrmul12_fa6_11_f_u_arrmul12_fa7_10_y2;
  wire f_u_arrmul12_fa6_11_y0;
  wire f_u_arrmul12_fa6_11_y1;
  wire f_u_arrmul12_fa6_11_f_u_arrmul12_fa5_11_y4;
  wire f_u_arrmul12_fa6_11_y2;
  wire f_u_arrmul12_fa6_11_y3;
  wire f_u_arrmul12_fa6_11_y4;
  wire f_u_arrmul12_and7_11_a_7;
  wire f_u_arrmul12_and7_11_b_11;
  wire f_u_arrmul12_and7_11_y0;
  wire f_u_arrmul12_fa7_11_f_u_arrmul12_and7_11_y0;
  wire f_u_arrmul12_fa7_11_f_u_arrmul12_fa8_10_y2;
  wire f_u_arrmul12_fa7_11_y0;
  wire f_u_arrmul12_fa7_11_y1;
  wire f_u_arrmul12_fa7_11_f_u_arrmul12_fa6_11_y4;
  wire f_u_arrmul12_fa7_11_y2;
  wire f_u_arrmul12_fa7_11_y3;
  wire f_u_arrmul12_fa7_11_y4;
  wire f_u_arrmul12_and8_11_a_8;
  wire f_u_arrmul12_and8_11_b_11;
  wire f_u_arrmul12_and8_11_y0;
  wire f_u_arrmul12_fa8_11_f_u_arrmul12_and8_11_y0;
  wire f_u_arrmul12_fa8_11_f_u_arrmul12_fa9_10_y2;
  wire f_u_arrmul12_fa8_11_y0;
  wire f_u_arrmul12_fa8_11_y1;
  wire f_u_arrmul12_fa8_11_f_u_arrmul12_fa7_11_y4;
  wire f_u_arrmul12_fa8_11_y2;
  wire f_u_arrmul12_fa8_11_y3;
  wire f_u_arrmul12_fa8_11_y4;
  wire f_u_arrmul12_and9_11_a_9;
  wire f_u_arrmul12_and9_11_b_11;
  wire f_u_arrmul12_and9_11_y0;
  wire f_u_arrmul12_fa9_11_f_u_arrmul12_and9_11_y0;
  wire f_u_arrmul12_fa9_11_f_u_arrmul12_fa10_10_y2;
  wire f_u_arrmul12_fa9_11_y0;
  wire f_u_arrmul12_fa9_11_y1;
  wire f_u_arrmul12_fa9_11_f_u_arrmul12_fa8_11_y4;
  wire f_u_arrmul12_fa9_11_y2;
  wire f_u_arrmul12_fa9_11_y3;
  wire f_u_arrmul12_fa9_11_y4;
  wire f_u_arrmul12_and10_11_a_10;
  wire f_u_arrmul12_and10_11_b_11;
  wire f_u_arrmul12_and10_11_y0;
  wire f_u_arrmul12_fa10_11_f_u_arrmul12_and10_11_y0;
  wire f_u_arrmul12_fa10_11_f_u_arrmul12_fa11_10_y2;
  wire f_u_arrmul12_fa10_11_y0;
  wire f_u_arrmul12_fa10_11_y1;
  wire f_u_arrmul12_fa10_11_f_u_arrmul12_fa9_11_y4;
  wire f_u_arrmul12_fa10_11_y2;
  wire f_u_arrmul12_fa10_11_y3;
  wire f_u_arrmul12_fa10_11_y4;
  wire f_u_arrmul12_and11_11_a_11;
  wire f_u_arrmul12_and11_11_b_11;
  wire f_u_arrmul12_and11_11_y0;
  wire f_u_arrmul12_fa11_11_f_u_arrmul12_and11_11_y0;
  wire f_u_arrmul12_fa11_11_f_u_arrmul12_fa11_10_y4;
  wire f_u_arrmul12_fa11_11_y0;
  wire f_u_arrmul12_fa11_11_y1;
  wire f_u_arrmul12_fa11_11_f_u_arrmul12_fa10_11_y4;
  wire f_u_arrmul12_fa11_11_y2;
  wire f_u_arrmul12_fa11_11_y3;
  wire f_u_arrmul12_fa11_11_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign f_u_arrmul12_and0_0_a_0 = a_0;
  assign f_u_arrmul12_and0_0_b_0 = b_0;
  assign f_u_arrmul12_and0_0_y0 = f_u_arrmul12_and0_0_a_0 & f_u_arrmul12_and0_0_b_0;
  assign f_u_arrmul12_and1_0_a_1 = a_1;
  assign f_u_arrmul12_and1_0_b_0 = b_0;
  assign f_u_arrmul12_and1_0_y0 = f_u_arrmul12_and1_0_a_1 & f_u_arrmul12_and1_0_b_0;
  assign f_u_arrmul12_and2_0_a_2 = a_2;
  assign f_u_arrmul12_and2_0_b_0 = b_0;
  assign f_u_arrmul12_and2_0_y0 = f_u_arrmul12_and2_0_a_2 & f_u_arrmul12_and2_0_b_0;
  assign f_u_arrmul12_and3_0_a_3 = a_3;
  assign f_u_arrmul12_and3_0_b_0 = b_0;
  assign f_u_arrmul12_and3_0_y0 = f_u_arrmul12_and3_0_a_3 & f_u_arrmul12_and3_0_b_0;
  assign f_u_arrmul12_and4_0_a_4 = a_4;
  assign f_u_arrmul12_and4_0_b_0 = b_0;
  assign f_u_arrmul12_and4_0_y0 = f_u_arrmul12_and4_0_a_4 & f_u_arrmul12_and4_0_b_0;
  assign f_u_arrmul12_and5_0_a_5 = a_5;
  assign f_u_arrmul12_and5_0_b_0 = b_0;
  assign f_u_arrmul12_and5_0_y0 = f_u_arrmul12_and5_0_a_5 & f_u_arrmul12_and5_0_b_0;
  assign f_u_arrmul12_and6_0_a_6 = a_6;
  assign f_u_arrmul12_and6_0_b_0 = b_0;
  assign f_u_arrmul12_and6_0_y0 = f_u_arrmul12_and6_0_a_6 & f_u_arrmul12_and6_0_b_0;
  assign f_u_arrmul12_and7_0_a_7 = a_7;
  assign f_u_arrmul12_and7_0_b_0 = b_0;
  assign f_u_arrmul12_and7_0_y0 = f_u_arrmul12_and7_0_a_7 & f_u_arrmul12_and7_0_b_0;
  assign f_u_arrmul12_and8_0_a_8 = a_8;
  assign f_u_arrmul12_and8_0_b_0 = b_0;
  assign f_u_arrmul12_and8_0_y0 = f_u_arrmul12_and8_0_a_8 & f_u_arrmul12_and8_0_b_0;
  assign f_u_arrmul12_and9_0_a_9 = a_9;
  assign f_u_arrmul12_and9_0_b_0 = b_0;
  assign f_u_arrmul12_and9_0_y0 = f_u_arrmul12_and9_0_a_9 & f_u_arrmul12_and9_0_b_0;
  assign f_u_arrmul12_and10_0_a_10 = a_10;
  assign f_u_arrmul12_and10_0_b_0 = b_0;
  assign f_u_arrmul12_and10_0_y0 = f_u_arrmul12_and10_0_a_10 & f_u_arrmul12_and10_0_b_0;
  assign f_u_arrmul12_and11_0_a_11 = a_11;
  assign f_u_arrmul12_and11_0_b_0 = b_0;
  assign f_u_arrmul12_and11_0_y0 = f_u_arrmul12_and11_0_a_11 & f_u_arrmul12_and11_0_b_0;
  assign f_u_arrmul12_and0_1_a_0 = a_0;
  assign f_u_arrmul12_and0_1_b_1 = b_1;
  assign f_u_arrmul12_and0_1_y0 = f_u_arrmul12_and0_1_a_0 & f_u_arrmul12_and0_1_b_1;
  assign f_u_arrmul12_ha0_1_f_u_arrmul12_and0_1_y0 = f_u_arrmul12_and0_1_y0;
  assign f_u_arrmul12_ha0_1_f_u_arrmul12_and1_0_y0 = f_u_arrmul12_and1_0_y0;
  assign f_u_arrmul12_ha0_1_y0 = f_u_arrmul12_ha0_1_f_u_arrmul12_and0_1_y0 ^ f_u_arrmul12_ha0_1_f_u_arrmul12_and1_0_y0;
  assign f_u_arrmul12_ha0_1_y1 = f_u_arrmul12_ha0_1_f_u_arrmul12_and0_1_y0 & f_u_arrmul12_ha0_1_f_u_arrmul12_and1_0_y0;
  assign f_u_arrmul12_and1_1_a_1 = a_1;
  assign f_u_arrmul12_and1_1_b_1 = b_1;
  assign f_u_arrmul12_and1_1_y0 = f_u_arrmul12_and1_1_a_1 & f_u_arrmul12_and1_1_b_1;
  assign f_u_arrmul12_fa1_1_f_u_arrmul12_and1_1_y0 = f_u_arrmul12_and1_1_y0;
  assign f_u_arrmul12_fa1_1_f_u_arrmul12_and2_0_y0 = f_u_arrmul12_and2_0_y0;
  assign f_u_arrmul12_fa1_1_f_u_arrmul12_ha0_1_y1 = f_u_arrmul12_ha0_1_y1;
  assign f_u_arrmul12_fa1_1_y0 = f_u_arrmul12_fa1_1_f_u_arrmul12_and1_1_y0 ^ f_u_arrmul12_fa1_1_f_u_arrmul12_and2_0_y0;
  assign f_u_arrmul12_fa1_1_y1 = f_u_arrmul12_fa1_1_f_u_arrmul12_and1_1_y0 & f_u_arrmul12_fa1_1_f_u_arrmul12_and2_0_y0;
  assign f_u_arrmul12_fa1_1_y2 = f_u_arrmul12_fa1_1_y0 ^ f_u_arrmul12_fa1_1_f_u_arrmul12_ha0_1_y1;
  assign f_u_arrmul12_fa1_1_y3 = f_u_arrmul12_fa1_1_y0 & f_u_arrmul12_fa1_1_f_u_arrmul12_ha0_1_y1;
  assign f_u_arrmul12_fa1_1_y4 = f_u_arrmul12_fa1_1_y1 | f_u_arrmul12_fa1_1_y3;
  assign f_u_arrmul12_and2_1_a_2 = a_2;
  assign f_u_arrmul12_and2_1_b_1 = b_1;
  assign f_u_arrmul12_and2_1_y0 = f_u_arrmul12_and2_1_a_2 & f_u_arrmul12_and2_1_b_1;
  assign f_u_arrmul12_fa2_1_f_u_arrmul12_and2_1_y0 = f_u_arrmul12_and2_1_y0;
  assign f_u_arrmul12_fa2_1_f_u_arrmul12_and3_0_y0 = f_u_arrmul12_and3_0_y0;
  assign f_u_arrmul12_fa2_1_f_u_arrmul12_fa1_1_y4 = f_u_arrmul12_fa1_1_y4;
  assign f_u_arrmul12_fa2_1_y0 = f_u_arrmul12_fa2_1_f_u_arrmul12_and2_1_y0 ^ f_u_arrmul12_fa2_1_f_u_arrmul12_and3_0_y0;
  assign f_u_arrmul12_fa2_1_y1 = f_u_arrmul12_fa2_1_f_u_arrmul12_and2_1_y0 & f_u_arrmul12_fa2_1_f_u_arrmul12_and3_0_y0;
  assign f_u_arrmul12_fa2_1_y2 = f_u_arrmul12_fa2_1_y0 ^ f_u_arrmul12_fa2_1_f_u_arrmul12_fa1_1_y4;
  assign f_u_arrmul12_fa2_1_y3 = f_u_arrmul12_fa2_1_y0 & f_u_arrmul12_fa2_1_f_u_arrmul12_fa1_1_y4;
  assign f_u_arrmul12_fa2_1_y4 = f_u_arrmul12_fa2_1_y1 | f_u_arrmul12_fa2_1_y3;
  assign f_u_arrmul12_and3_1_a_3 = a_3;
  assign f_u_arrmul12_and3_1_b_1 = b_1;
  assign f_u_arrmul12_and3_1_y0 = f_u_arrmul12_and3_1_a_3 & f_u_arrmul12_and3_1_b_1;
  assign f_u_arrmul12_fa3_1_f_u_arrmul12_and3_1_y0 = f_u_arrmul12_and3_1_y0;
  assign f_u_arrmul12_fa3_1_f_u_arrmul12_and4_0_y0 = f_u_arrmul12_and4_0_y0;
  assign f_u_arrmul12_fa3_1_f_u_arrmul12_fa2_1_y4 = f_u_arrmul12_fa2_1_y4;
  assign f_u_arrmul12_fa3_1_y0 = f_u_arrmul12_fa3_1_f_u_arrmul12_and3_1_y0 ^ f_u_arrmul12_fa3_1_f_u_arrmul12_and4_0_y0;
  assign f_u_arrmul12_fa3_1_y1 = f_u_arrmul12_fa3_1_f_u_arrmul12_and3_1_y0 & f_u_arrmul12_fa3_1_f_u_arrmul12_and4_0_y0;
  assign f_u_arrmul12_fa3_1_y2 = f_u_arrmul12_fa3_1_y0 ^ f_u_arrmul12_fa3_1_f_u_arrmul12_fa2_1_y4;
  assign f_u_arrmul12_fa3_1_y3 = f_u_arrmul12_fa3_1_y0 & f_u_arrmul12_fa3_1_f_u_arrmul12_fa2_1_y4;
  assign f_u_arrmul12_fa3_1_y4 = f_u_arrmul12_fa3_1_y1 | f_u_arrmul12_fa3_1_y3;
  assign f_u_arrmul12_and4_1_a_4 = a_4;
  assign f_u_arrmul12_and4_1_b_1 = b_1;
  assign f_u_arrmul12_and4_1_y0 = f_u_arrmul12_and4_1_a_4 & f_u_arrmul12_and4_1_b_1;
  assign f_u_arrmul12_fa4_1_f_u_arrmul12_and4_1_y0 = f_u_arrmul12_and4_1_y0;
  assign f_u_arrmul12_fa4_1_f_u_arrmul12_and5_0_y0 = f_u_arrmul12_and5_0_y0;
  assign f_u_arrmul12_fa4_1_f_u_arrmul12_fa3_1_y4 = f_u_arrmul12_fa3_1_y4;
  assign f_u_arrmul12_fa4_1_y0 = f_u_arrmul12_fa4_1_f_u_arrmul12_and4_1_y0 ^ f_u_arrmul12_fa4_1_f_u_arrmul12_and5_0_y0;
  assign f_u_arrmul12_fa4_1_y1 = f_u_arrmul12_fa4_1_f_u_arrmul12_and4_1_y0 & f_u_arrmul12_fa4_1_f_u_arrmul12_and5_0_y0;
  assign f_u_arrmul12_fa4_1_y2 = f_u_arrmul12_fa4_1_y0 ^ f_u_arrmul12_fa4_1_f_u_arrmul12_fa3_1_y4;
  assign f_u_arrmul12_fa4_1_y3 = f_u_arrmul12_fa4_1_y0 & f_u_arrmul12_fa4_1_f_u_arrmul12_fa3_1_y4;
  assign f_u_arrmul12_fa4_1_y4 = f_u_arrmul12_fa4_1_y1 | f_u_arrmul12_fa4_1_y3;
  assign f_u_arrmul12_and5_1_a_5 = a_5;
  assign f_u_arrmul12_and5_1_b_1 = b_1;
  assign f_u_arrmul12_and5_1_y0 = f_u_arrmul12_and5_1_a_5 & f_u_arrmul12_and5_1_b_1;
  assign f_u_arrmul12_fa5_1_f_u_arrmul12_and5_1_y0 = f_u_arrmul12_and5_1_y0;
  assign f_u_arrmul12_fa5_1_f_u_arrmul12_and6_0_y0 = f_u_arrmul12_and6_0_y0;
  assign f_u_arrmul12_fa5_1_f_u_arrmul12_fa4_1_y4 = f_u_arrmul12_fa4_1_y4;
  assign f_u_arrmul12_fa5_1_y0 = f_u_arrmul12_fa5_1_f_u_arrmul12_and5_1_y0 ^ f_u_arrmul12_fa5_1_f_u_arrmul12_and6_0_y0;
  assign f_u_arrmul12_fa5_1_y1 = f_u_arrmul12_fa5_1_f_u_arrmul12_and5_1_y0 & f_u_arrmul12_fa5_1_f_u_arrmul12_and6_0_y0;
  assign f_u_arrmul12_fa5_1_y2 = f_u_arrmul12_fa5_1_y0 ^ f_u_arrmul12_fa5_1_f_u_arrmul12_fa4_1_y4;
  assign f_u_arrmul12_fa5_1_y3 = f_u_arrmul12_fa5_1_y0 & f_u_arrmul12_fa5_1_f_u_arrmul12_fa4_1_y4;
  assign f_u_arrmul12_fa5_1_y4 = f_u_arrmul12_fa5_1_y1 | f_u_arrmul12_fa5_1_y3;
  assign f_u_arrmul12_and6_1_a_6 = a_6;
  assign f_u_arrmul12_and6_1_b_1 = b_1;
  assign f_u_arrmul12_and6_1_y0 = f_u_arrmul12_and6_1_a_6 & f_u_arrmul12_and6_1_b_1;
  assign f_u_arrmul12_fa6_1_f_u_arrmul12_and6_1_y0 = f_u_arrmul12_and6_1_y0;
  assign f_u_arrmul12_fa6_1_f_u_arrmul12_and7_0_y0 = f_u_arrmul12_and7_0_y0;
  assign f_u_arrmul12_fa6_1_f_u_arrmul12_fa5_1_y4 = f_u_arrmul12_fa5_1_y4;
  assign f_u_arrmul12_fa6_1_y0 = f_u_arrmul12_fa6_1_f_u_arrmul12_and6_1_y0 ^ f_u_arrmul12_fa6_1_f_u_arrmul12_and7_0_y0;
  assign f_u_arrmul12_fa6_1_y1 = f_u_arrmul12_fa6_1_f_u_arrmul12_and6_1_y0 & f_u_arrmul12_fa6_1_f_u_arrmul12_and7_0_y0;
  assign f_u_arrmul12_fa6_1_y2 = f_u_arrmul12_fa6_1_y0 ^ f_u_arrmul12_fa6_1_f_u_arrmul12_fa5_1_y4;
  assign f_u_arrmul12_fa6_1_y3 = f_u_arrmul12_fa6_1_y0 & f_u_arrmul12_fa6_1_f_u_arrmul12_fa5_1_y4;
  assign f_u_arrmul12_fa6_1_y4 = f_u_arrmul12_fa6_1_y1 | f_u_arrmul12_fa6_1_y3;
  assign f_u_arrmul12_and7_1_a_7 = a_7;
  assign f_u_arrmul12_and7_1_b_1 = b_1;
  assign f_u_arrmul12_and7_1_y0 = f_u_arrmul12_and7_1_a_7 & f_u_arrmul12_and7_1_b_1;
  assign f_u_arrmul12_fa7_1_f_u_arrmul12_and7_1_y0 = f_u_arrmul12_and7_1_y0;
  assign f_u_arrmul12_fa7_1_f_u_arrmul12_and8_0_y0 = f_u_arrmul12_and8_0_y0;
  assign f_u_arrmul12_fa7_1_f_u_arrmul12_fa6_1_y4 = f_u_arrmul12_fa6_1_y4;
  assign f_u_arrmul12_fa7_1_y0 = f_u_arrmul12_fa7_1_f_u_arrmul12_and7_1_y0 ^ f_u_arrmul12_fa7_1_f_u_arrmul12_and8_0_y0;
  assign f_u_arrmul12_fa7_1_y1 = f_u_arrmul12_fa7_1_f_u_arrmul12_and7_1_y0 & f_u_arrmul12_fa7_1_f_u_arrmul12_and8_0_y0;
  assign f_u_arrmul12_fa7_1_y2 = f_u_arrmul12_fa7_1_y0 ^ f_u_arrmul12_fa7_1_f_u_arrmul12_fa6_1_y4;
  assign f_u_arrmul12_fa7_1_y3 = f_u_arrmul12_fa7_1_y0 & f_u_arrmul12_fa7_1_f_u_arrmul12_fa6_1_y4;
  assign f_u_arrmul12_fa7_1_y4 = f_u_arrmul12_fa7_1_y1 | f_u_arrmul12_fa7_1_y3;
  assign f_u_arrmul12_and8_1_a_8 = a_8;
  assign f_u_arrmul12_and8_1_b_1 = b_1;
  assign f_u_arrmul12_and8_1_y0 = f_u_arrmul12_and8_1_a_8 & f_u_arrmul12_and8_1_b_1;
  assign f_u_arrmul12_fa8_1_f_u_arrmul12_and8_1_y0 = f_u_arrmul12_and8_1_y0;
  assign f_u_arrmul12_fa8_1_f_u_arrmul12_and9_0_y0 = f_u_arrmul12_and9_0_y0;
  assign f_u_arrmul12_fa8_1_f_u_arrmul12_fa7_1_y4 = f_u_arrmul12_fa7_1_y4;
  assign f_u_arrmul12_fa8_1_y0 = f_u_arrmul12_fa8_1_f_u_arrmul12_and8_1_y0 ^ f_u_arrmul12_fa8_1_f_u_arrmul12_and9_0_y0;
  assign f_u_arrmul12_fa8_1_y1 = f_u_arrmul12_fa8_1_f_u_arrmul12_and8_1_y0 & f_u_arrmul12_fa8_1_f_u_arrmul12_and9_0_y0;
  assign f_u_arrmul12_fa8_1_y2 = f_u_arrmul12_fa8_1_y0 ^ f_u_arrmul12_fa8_1_f_u_arrmul12_fa7_1_y4;
  assign f_u_arrmul12_fa8_1_y3 = f_u_arrmul12_fa8_1_y0 & f_u_arrmul12_fa8_1_f_u_arrmul12_fa7_1_y4;
  assign f_u_arrmul12_fa8_1_y4 = f_u_arrmul12_fa8_1_y1 | f_u_arrmul12_fa8_1_y3;
  assign f_u_arrmul12_and9_1_a_9 = a_9;
  assign f_u_arrmul12_and9_1_b_1 = b_1;
  assign f_u_arrmul12_and9_1_y0 = f_u_arrmul12_and9_1_a_9 & f_u_arrmul12_and9_1_b_1;
  assign f_u_arrmul12_fa9_1_f_u_arrmul12_and9_1_y0 = f_u_arrmul12_and9_1_y0;
  assign f_u_arrmul12_fa9_1_f_u_arrmul12_and10_0_y0 = f_u_arrmul12_and10_0_y0;
  assign f_u_arrmul12_fa9_1_f_u_arrmul12_fa8_1_y4 = f_u_arrmul12_fa8_1_y4;
  assign f_u_arrmul12_fa9_1_y0 = f_u_arrmul12_fa9_1_f_u_arrmul12_and9_1_y0 ^ f_u_arrmul12_fa9_1_f_u_arrmul12_and10_0_y0;
  assign f_u_arrmul12_fa9_1_y1 = f_u_arrmul12_fa9_1_f_u_arrmul12_and9_1_y0 & f_u_arrmul12_fa9_1_f_u_arrmul12_and10_0_y0;
  assign f_u_arrmul12_fa9_1_y2 = f_u_arrmul12_fa9_1_y0 ^ f_u_arrmul12_fa9_1_f_u_arrmul12_fa8_1_y4;
  assign f_u_arrmul12_fa9_1_y3 = f_u_arrmul12_fa9_1_y0 & f_u_arrmul12_fa9_1_f_u_arrmul12_fa8_1_y4;
  assign f_u_arrmul12_fa9_1_y4 = f_u_arrmul12_fa9_1_y1 | f_u_arrmul12_fa9_1_y3;
  assign f_u_arrmul12_and10_1_a_10 = a_10;
  assign f_u_arrmul12_and10_1_b_1 = b_1;
  assign f_u_arrmul12_and10_1_y0 = f_u_arrmul12_and10_1_a_10 & f_u_arrmul12_and10_1_b_1;
  assign f_u_arrmul12_fa10_1_f_u_arrmul12_and10_1_y0 = f_u_arrmul12_and10_1_y0;
  assign f_u_arrmul12_fa10_1_f_u_arrmul12_and11_0_y0 = f_u_arrmul12_and11_0_y0;
  assign f_u_arrmul12_fa10_1_f_u_arrmul12_fa9_1_y4 = f_u_arrmul12_fa9_1_y4;
  assign f_u_arrmul12_fa10_1_y0 = f_u_arrmul12_fa10_1_f_u_arrmul12_and10_1_y0 ^ f_u_arrmul12_fa10_1_f_u_arrmul12_and11_0_y0;
  assign f_u_arrmul12_fa10_1_y1 = f_u_arrmul12_fa10_1_f_u_arrmul12_and10_1_y0 & f_u_arrmul12_fa10_1_f_u_arrmul12_and11_0_y0;
  assign f_u_arrmul12_fa10_1_y2 = f_u_arrmul12_fa10_1_y0 ^ f_u_arrmul12_fa10_1_f_u_arrmul12_fa9_1_y4;
  assign f_u_arrmul12_fa10_1_y3 = f_u_arrmul12_fa10_1_y0 & f_u_arrmul12_fa10_1_f_u_arrmul12_fa9_1_y4;
  assign f_u_arrmul12_fa10_1_y4 = f_u_arrmul12_fa10_1_y1 | f_u_arrmul12_fa10_1_y3;
  assign f_u_arrmul12_and11_1_a_11 = a_11;
  assign f_u_arrmul12_and11_1_b_1 = b_1;
  assign f_u_arrmul12_and11_1_y0 = f_u_arrmul12_and11_1_a_11 & f_u_arrmul12_and11_1_b_1;
  assign f_u_arrmul12_ha11_1_f_u_arrmul12_and11_1_y0 = f_u_arrmul12_and11_1_y0;
  assign f_u_arrmul12_ha11_1_f_u_arrmul12_fa10_1_y4 = f_u_arrmul12_fa10_1_y4;
  assign f_u_arrmul12_ha11_1_y0 = f_u_arrmul12_ha11_1_f_u_arrmul12_and11_1_y0 ^ f_u_arrmul12_ha11_1_f_u_arrmul12_fa10_1_y4;
  assign f_u_arrmul12_ha11_1_y1 = f_u_arrmul12_ha11_1_f_u_arrmul12_and11_1_y0 & f_u_arrmul12_ha11_1_f_u_arrmul12_fa10_1_y4;
  assign f_u_arrmul12_and0_2_a_0 = a_0;
  assign f_u_arrmul12_and0_2_b_2 = b_2;
  assign f_u_arrmul12_and0_2_y0 = f_u_arrmul12_and0_2_a_0 & f_u_arrmul12_and0_2_b_2;
  assign f_u_arrmul12_ha0_2_f_u_arrmul12_and0_2_y0 = f_u_arrmul12_and0_2_y0;
  assign f_u_arrmul12_ha0_2_f_u_arrmul12_fa1_1_y2 = f_u_arrmul12_fa1_1_y2;
  assign f_u_arrmul12_ha0_2_y0 = f_u_arrmul12_ha0_2_f_u_arrmul12_and0_2_y0 ^ f_u_arrmul12_ha0_2_f_u_arrmul12_fa1_1_y2;
  assign f_u_arrmul12_ha0_2_y1 = f_u_arrmul12_ha0_2_f_u_arrmul12_and0_2_y0 & f_u_arrmul12_ha0_2_f_u_arrmul12_fa1_1_y2;
  assign f_u_arrmul12_and1_2_a_1 = a_1;
  assign f_u_arrmul12_and1_2_b_2 = b_2;
  assign f_u_arrmul12_and1_2_y0 = f_u_arrmul12_and1_2_a_1 & f_u_arrmul12_and1_2_b_2;
  assign f_u_arrmul12_fa1_2_f_u_arrmul12_and1_2_y0 = f_u_arrmul12_and1_2_y0;
  assign f_u_arrmul12_fa1_2_f_u_arrmul12_fa2_1_y2 = f_u_arrmul12_fa2_1_y2;
  assign f_u_arrmul12_fa1_2_f_u_arrmul12_ha0_2_y1 = f_u_arrmul12_ha0_2_y1;
  assign f_u_arrmul12_fa1_2_y0 = f_u_arrmul12_fa1_2_f_u_arrmul12_and1_2_y0 ^ f_u_arrmul12_fa1_2_f_u_arrmul12_fa2_1_y2;
  assign f_u_arrmul12_fa1_2_y1 = f_u_arrmul12_fa1_2_f_u_arrmul12_and1_2_y0 & f_u_arrmul12_fa1_2_f_u_arrmul12_fa2_1_y2;
  assign f_u_arrmul12_fa1_2_y2 = f_u_arrmul12_fa1_2_y0 ^ f_u_arrmul12_fa1_2_f_u_arrmul12_ha0_2_y1;
  assign f_u_arrmul12_fa1_2_y3 = f_u_arrmul12_fa1_2_y0 & f_u_arrmul12_fa1_2_f_u_arrmul12_ha0_2_y1;
  assign f_u_arrmul12_fa1_2_y4 = f_u_arrmul12_fa1_2_y1 | f_u_arrmul12_fa1_2_y3;
  assign f_u_arrmul12_and2_2_a_2 = a_2;
  assign f_u_arrmul12_and2_2_b_2 = b_2;
  assign f_u_arrmul12_and2_2_y0 = f_u_arrmul12_and2_2_a_2 & f_u_arrmul12_and2_2_b_2;
  assign f_u_arrmul12_fa2_2_f_u_arrmul12_and2_2_y0 = f_u_arrmul12_and2_2_y0;
  assign f_u_arrmul12_fa2_2_f_u_arrmul12_fa3_1_y2 = f_u_arrmul12_fa3_1_y2;
  assign f_u_arrmul12_fa2_2_f_u_arrmul12_fa1_2_y4 = f_u_arrmul12_fa1_2_y4;
  assign f_u_arrmul12_fa2_2_y0 = f_u_arrmul12_fa2_2_f_u_arrmul12_and2_2_y0 ^ f_u_arrmul12_fa2_2_f_u_arrmul12_fa3_1_y2;
  assign f_u_arrmul12_fa2_2_y1 = f_u_arrmul12_fa2_2_f_u_arrmul12_and2_2_y0 & f_u_arrmul12_fa2_2_f_u_arrmul12_fa3_1_y2;
  assign f_u_arrmul12_fa2_2_y2 = f_u_arrmul12_fa2_2_y0 ^ f_u_arrmul12_fa2_2_f_u_arrmul12_fa1_2_y4;
  assign f_u_arrmul12_fa2_2_y3 = f_u_arrmul12_fa2_2_y0 & f_u_arrmul12_fa2_2_f_u_arrmul12_fa1_2_y4;
  assign f_u_arrmul12_fa2_2_y4 = f_u_arrmul12_fa2_2_y1 | f_u_arrmul12_fa2_2_y3;
  assign f_u_arrmul12_and3_2_a_3 = a_3;
  assign f_u_arrmul12_and3_2_b_2 = b_2;
  assign f_u_arrmul12_and3_2_y0 = f_u_arrmul12_and3_2_a_3 & f_u_arrmul12_and3_2_b_2;
  assign f_u_arrmul12_fa3_2_f_u_arrmul12_and3_2_y0 = f_u_arrmul12_and3_2_y0;
  assign f_u_arrmul12_fa3_2_f_u_arrmul12_fa4_1_y2 = f_u_arrmul12_fa4_1_y2;
  assign f_u_arrmul12_fa3_2_f_u_arrmul12_fa2_2_y4 = f_u_arrmul12_fa2_2_y4;
  assign f_u_arrmul12_fa3_2_y0 = f_u_arrmul12_fa3_2_f_u_arrmul12_and3_2_y0 ^ f_u_arrmul12_fa3_2_f_u_arrmul12_fa4_1_y2;
  assign f_u_arrmul12_fa3_2_y1 = f_u_arrmul12_fa3_2_f_u_arrmul12_and3_2_y0 & f_u_arrmul12_fa3_2_f_u_arrmul12_fa4_1_y2;
  assign f_u_arrmul12_fa3_2_y2 = f_u_arrmul12_fa3_2_y0 ^ f_u_arrmul12_fa3_2_f_u_arrmul12_fa2_2_y4;
  assign f_u_arrmul12_fa3_2_y3 = f_u_arrmul12_fa3_2_y0 & f_u_arrmul12_fa3_2_f_u_arrmul12_fa2_2_y4;
  assign f_u_arrmul12_fa3_2_y4 = f_u_arrmul12_fa3_2_y1 | f_u_arrmul12_fa3_2_y3;
  assign f_u_arrmul12_and4_2_a_4 = a_4;
  assign f_u_arrmul12_and4_2_b_2 = b_2;
  assign f_u_arrmul12_and4_2_y0 = f_u_arrmul12_and4_2_a_4 & f_u_arrmul12_and4_2_b_2;
  assign f_u_arrmul12_fa4_2_f_u_arrmul12_and4_2_y0 = f_u_arrmul12_and4_2_y0;
  assign f_u_arrmul12_fa4_2_f_u_arrmul12_fa5_1_y2 = f_u_arrmul12_fa5_1_y2;
  assign f_u_arrmul12_fa4_2_f_u_arrmul12_fa3_2_y4 = f_u_arrmul12_fa3_2_y4;
  assign f_u_arrmul12_fa4_2_y0 = f_u_arrmul12_fa4_2_f_u_arrmul12_and4_2_y0 ^ f_u_arrmul12_fa4_2_f_u_arrmul12_fa5_1_y2;
  assign f_u_arrmul12_fa4_2_y1 = f_u_arrmul12_fa4_2_f_u_arrmul12_and4_2_y0 & f_u_arrmul12_fa4_2_f_u_arrmul12_fa5_1_y2;
  assign f_u_arrmul12_fa4_2_y2 = f_u_arrmul12_fa4_2_y0 ^ f_u_arrmul12_fa4_2_f_u_arrmul12_fa3_2_y4;
  assign f_u_arrmul12_fa4_2_y3 = f_u_arrmul12_fa4_2_y0 & f_u_arrmul12_fa4_2_f_u_arrmul12_fa3_2_y4;
  assign f_u_arrmul12_fa4_2_y4 = f_u_arrmul12_fa4_2_y1 | f_u_arrmul12_fa4_2_y3;
  assign f_u_arrmul12_and5_2_a_5 = a_5;
  assign f_u_arrmul12_and5_2_b_2 = b_2;
  assign f_u_arrmul12_and5_2_y0 = f_u_arrmul12_and5_2_a_5 & f_u_arrmul12_and5_2_b_2;
  assign f_u_arrmul12_fa5_2_f_u_arrmul12_and5_2_y0 = f_u_arrmul12_and5_2_y0;
  assign f_u_arrmul12_fa5_2_f_u_arrmul12_fa6_1_y2 = f_u_arrmul12_fa6_1_y2;
  assign f_u_arrmul12_fa5_2_f_u_arrmul12_fa4_2_y4 = f_u_arrmul12_fa4_2_y4;
  assign f_u_arrmul12_fa5_2_y0 = f_u_arrmul12_fa5_2_f_u_arrmul12_and5_2_y0 ^ f_u_arrmul12_fa5_2_f_u_arrmul12_fa6_1_y2;
  assign f_u_arrmul12_fa5_2_y1 = f_u_arrmul12_fa5_2_f_u_arrmul12_and5_2_y0 & f_u_arrmul12_fa5_2_f_u_arrmul12_fa6_1_y2;
  assign f_u_arrmul12_fa5_2_y2 = f_u_arrmul12_fa5_2_y0 ^ f_u_arrmul12_fa5_2_f_u_arrmul12_fa4_2_y4;
  assign f_u_arrmul12_fa5_2_y3 = f_u_arrmul12_fa5_2_y0 & f_u_arrmul12_fa5_2_f_u_arrmul12_fa4_2_y4;
  assign f_u_arrmul12_fa5_2_y4 = f_u_arrmul12_fa5_2_y1 | f_u_arrmul12_fa5_2_y3;
  assign f_u_arrmul12_and6_2_a_6 = a_6;
  assign f_u_arrmul12_and6_2_b_2 = b_2;
  assign f_u_arrmul12_and6_2_y0 = f_u_arrmul12_and6_2_a_6 & f_u_arrmul12_and6_2_b_2;
  assign f_u_arrmul12_fa6_2_f_u_arrmul12_and6_2_y0 = f_u_arrmul12_and6_2_y0;
  assign f_u_arrmul12_fa6_2_f_u_arrmul12_fa7_1_y2 = f_u_arrmul12_fa7_1_y2;
  assign f_u_arrmul12_fa6_2_f_u_arrmul12_fa5_2_y4 = f_u_arrmul12_fa5_2_y4;
  assign f_u_arrmul12_fa6_2_y0 = f_u_arrmul12_fa6_2_f_u_arrmul12_and6_2_y0 ^ f_u_arrmul12_fa6_2_f_u_arrmul12_fa7_1_y2;
  assign f_u_arrmul12_fa6_2_y1 = f_u_arrmul12_fa6_2_f_u_arrmul12_and6_2_y0 & f_u_arrmul12_fa6_2_f_u_arrmul12_fa7_1_y2;
  assign f_u_arrmul12_fa6_2_y2 = f_u_arrmul12_fa6_2_y0 ^ f_u_arrmul12_fa6_2_f_u_arrmul12_fa5_2_y4;
  assign f_u_arrmul12_fa6_2_y3 = f_u_arrmul12_fa6_2_y0 & f_u_arrmul12_fa6_2_f_u_arrmul12_fa5_2_y4;
  assign f_u_arrmul12_fa6_2_y4 = f_u_arrmul12_fa6_2_y1 | f_u_arrmul12_fa6_2_y3;
  assign f_u_arrmul12_and7_2_a_7 = a_7;
  assign f_u_arrmul12_and7_2_b_2 = b_2;
  assign f_u_arrmul12_and7_2_y0 = f_u_arrmul12_and7_2_a_7 & f_u_arrmul12_and7_2_b_2;
  assign f_u_arrmul12_fa7_2_f_u_arrmul12_and7_2_y0 = f_u_arrmul12_and7_2_y0;
  assign f_u_arrmul12_fa7_2_f_u_arrmul12_fa8_1_y2 = f_u_arrmul12_fa8_1_y2;
  assign f_u_arrmul12_fa7_2_f_u_arrmul12_fa6_2_y4 = f_u_arrmul12_fa6_2_y4;
  assign f_u_arrmul12_fa7_2_y0 = f_u_arrmul12_fa7_2_f_u_arrmul12_and7_2_y0 ^ f_u_arrmul12_fa7_2_f_u_arrmul12_fa8_1_y2;
  assign f_u_arrmul12_fa7_2_y1 = f_u_arrmul12_fa7_2_f_u_arrmul12_and7_2_y0 & f_u_arrmul12_fa7_2_f_u_arrmul12_fa8_1_y2;
  assign f_u_arrmul12_fa7_2_y2 = f_u_arrmul12_fa7_2_y0 ^ f_u_arrmul12_fa7_2_f_u_arrmul12_fa6_2_y4;
  assign f_u_arrmul12_fa7_2_y3 = f_u_arrmul12_fa7_2_y0 & f_u_arrmul12_fa7_2_f_u_arrmul12_fa6_2_y4;
  assign f_u_arrmul12_fa7_2_y4 = f_u_arrmul12_fa7_2_y1 | f_u_arrmul12_fa7_2_y3;
  assign f_u_arrmul12_and8_2_a_8 = a_8;
  assign f_u_arrmul12_and8_2_b_2 = b_2;
  assign f_u_arrmul12_and8_2_y0 = f_u_arrmul12_and8_2_a_8 & f_u_arrmul12_and8_2_b_2;
  assign f_u_arrmul12_fa8_2_f_u_arrmul12_and8_2_y0 = f_u_arrmul12_and8_2_y0;
  assign f_u_arrmul12_fa8_2_f_u_arrmul12_fa9_1_y2 = f_u_arrmul12_fa9_1_y2;
  assign f_u_arrmul12_fa8_2_f_u_arrmul12_fa7_2_y4 = f_u_arrmul12_fa7_2_y4;
  assign f_u_arrmul12_fa8_2_y0 = f_u_arrmul12_fa8_2_f_u_arrmul12_and8_2_y0 ^ f_u_arrmul12_fa8_2_f_u_arrmul12_fa9_1_y2;
  assign f_u_arrmul12_fa8_2_y1 = f_u_arrmul12_fa8_2_f_u_arrmul12_and8_2_y0 & f_u_arrmul12_fa8_2_f_u_arrmul12_fa9_1_y2;
  assign f_u_arrmul12_fa8_2_y2 = f_u_arrmul12_fa8_2_y0 ^ f_u_arrmul12_fa8_2_f_u_arrmul12_fa7_2_y4;
  assign f_u_arrmul12_fa8_2_y3 = f_u_arrmul12_fa8_2_y0 & f_u_arrmul12_fa8_2_f_u_arrmul12_fa7_2_y4;
  assign f_u_arrmul12_fa8_2_y4 = f_u_arrmul12_fa8_2_y1 | f_u_arrmul12_fa8_2_y3;
  assign f_u_arrmul12_and9_2_a_9 = a_9;
  assign f_u_arrmul12_and9_2_b_2 = b_2;
  assign f_u_arrmul12_and9_2_y0 = f_u_arrmul12_and9_2_a_9 & f_u_arrmul12_and9_2_b_2;
  assign f_u_arrmul12_fa9_2_f_u_arrmul12_and9_2_y0 = f_u_arrmul12_and9_2_y0;
  assign f_u_arrmul12_fa9_2_f_u_arrmul12_fa10_1_y2 = f_u_arrmul12_fa10_1_y2;
  assign f_u_arrmul12_fa9_2_f_u_arrmul12_fa8_2_y4 = f_u_arrmul12_fa8_2_y4;
  assign f_u_arrmul12_fa9_2_y0 = f_u_arrmul12_fa9_2_f_u_arrmul12_and9_2_y0 ^ f_u_arrmul12_fa9_2_f_u_arrmul12_fa10_1_y2;
  assign f_u_arrmul12_fa9_2_y1 = f_u_arrmul12_fa9_2_f_u_arrmul12_and9_2_y0 & f_u_arrmul12_fa9_2_f_u_arrmul12_fa10_1_y2;
  assign f_u_arrmul12_fa9_2_y2 = f_u_arrmul12_fa9_2_y0 ^ f_u_arrmul12_fa9_2_f_u_arrmul12_fa8_2_y4;
  assign f_u_arrmul12_fa9_2_y3 = f_u_arrmul12_fa9_2_y0 & f_u_arrmul12_fa9_2_f_u_arrmul12_fa8_2_y4;
  assign f_u_arrmul12_fa9_2_y4 = f_u_arrmul12_fa9_2_y1 | f_u_arrmul12_fa9_2_y3;
  assign f_u_arrmul12_and10_2_a_10 = a_10;
  assign f_u_arrmul12_and10_2_b_2 = b_2;
  assign f_u_arrmul12_and10_2_y0 = f_u_arrmul12_and10_2_a_10 & f_u_arrmul12_and10_2_b_2;
  assign f_u_arrmul12_fa10_2_f_u_arrmul12_and10_2_y0 = f_u_arrmul12_and10_2_y0;
  assign f_u_arrmul12_fa10_2_f_u_arrmul12_ha11_1_y0 = f_u_arrmul12_ha11_1_y0;
  assign f_u_arrmul12_fa10_2_f_u_arrmul12_fa9_2_y4 = f_u_arrmul12_fa9_2_y4;
  assign f_u_arrmul12_fa10_2_y0 = f_u_arrmul12_fa10_2_f_u_arrmul12_and10_2_y0 ^ f_u_arrmul12_fa10_2_f_u_arrmul12_ha11_1_y0;
  assign f_u_arrmul12_fa10_2_y1 = f_u_arrmul12_fa10_2_f_u_arrmul12_and10_2_y0 & f_u_arrmul12_fa10_2_f_u_arrmul12_ha11_1_y0;
  assign f_u_arrmul12_fa10_2_y2 = f_u_arrmul12_fa10_2_y0 ^ f_u_arrmul12_fa10_2_f_u_arrmul12_fa9_2_y4;
  assign f_u_arrmul12_fa10_2_y3 = f_u_arrmul12_fa10_2_y0 & f_u_arrmul12_fa10_2_f_u_arrmul12_fa9_2_y4;
  assign f_u_arrmul12_fa10_2_y4 = f_u_arrmul12_fa10_2_y1 | f_u_arrmul12_fa10_2_y3;
  assign f_u_arrmul12_and11_2_a_11 = a_11;
  assign f_u_arrmul12_and11_2_b_2 = b_2;
  assign f_u_arrmul12_and11_2_y0 = f_u_arrmul12_and11_2_a_11 & f_u_arrmul12_and11_2_b_2;
  assign f_u_arrmul12_fa11_2_f_u_arrmul12_and11_2_y0 = f_u_arrmul12_and11_2_y0;
  assign f_u_arrmul12_fa11_2_f_u_arrmul12_ha11_1_y1 = f_u_arrmul12_ha11_1_y1;
  assign f_u_arrmul12_fa11_2_f_u_arrmul12_fa10_2_y4 = f_u_arrmul12_fa10_2_y4;
  assign f_u_arrmul12_fa11_2_y0 = f_u_arrmul12_fa11_2_f_u_arrmul12_and11_2_y0 ^ f_u_arrmul12_fa11_2_f_u_arrmul12_ha11_1_y1;
  assign f_u_arrmul12_fa11_2_y1 = f_u_arrmul12_fa11_2_f_u_arrmul12_and11_2_y0 & f_u_arrmul12_fa11_2_f_u_arrmul12_ha11_1_y1;
  assign f_u_arrmul12_fa11_2_y2 = f_u_arrmul12_fa11_2_y0 ^ f_u_arrmul12_fa11_2_f_u_arrmul12_fa10_2_y4;
  assign f_u_arrmul12_fa11_2_y3 = f_u_arrmul12_fa11_2_y0 & f_u_arrmul12_fa11_2_f_u_arrmul12_fa10_2_y4;
  assign f_u_arrmul12_fa11_2_y4 = f_u_arrmul12_fa11_2_y1 | f_u_arrmul12_fa11_2_y3;
  assign f_u_arrmul12_and0_3_a_0 = a_0;
  assign f_u_arrmul12_and0_3_b_3 = b_3;
  assign f_u_arrmul12_and0_3_y0 = f_u_arrmul12_and0_3_a_0 & f_u_arrmul12_and0_3_b_3;
  assign f_u_arrmul12_ha0_3_f_u_arrmul12_and0_3_y0 = f_u_arrmul12_and0_3_y0;
  assign f_u_arrmul12_ha0_3_f_u_arrmul12_fa1_2_y2 = f_u_arrmul12_fa1_2_y2;
  assign f_u_arrmul12_ha0_3_y0 = f_u_arrmul12_ha0_3_f_u_arrmul12_and0_3_y0 ^ f_u_arrmul12_ha0_3_f_u_arrmul12_fa1_2_y2;
  assign f_u_arrmul12_ha0_3_y1 = f_u_arrmul12_ha0_3_f_u_arrmul12_and0_3_y0 & f_u_arrmul12_ha0_3_f_u_arrmul12_fa1_2_y2;
  assign f_u_arrmul12_and1_3_a_1 = a_1;
  assign f_u_arrmul12_and1_3_b_3 = b_3;
  assign f_u_arrmul12_and1_3_y0 = f_u_arrmul12_and1_3_a_1 & f_u_arrmul12_and1_3_b_3;
  assign f_u_arrmul12_fa1_3_f_u_arrmul12_and1_3_y0 = f_u_arrmul12_and1_3_y0;
  assign f_u_arrmul12_fa1_3_f_u_arrmul12_fa2_2_y2 = f_u_arrmul12_fa2_2_y2;
  assign f_u_arrmul12_fa1_3_f_u_arrmul12_ha0_3_y1 = f_u_arrmul12_ha0_3_y1;
  assign f_u_arrmul12_fa1_3_y0 = f_u_arrmul12_fa1_3_f_u_arrmul12_and1_3_y0 ^ f_u_arrmul12_fa1_3_f_u_arrmul12_fa2_2_y2;
  assign f_u_arrmul12_fa1_3_y1 = f_u_arrmul12_fa1_3_f_u_arrmul12_and1_3_y0 & f_u_arrmul12_fa1_3_f_u_arrmul12_fa2_2_y2;
  assign f_u_arrmul12_fa1_3_y2 = f_u_arrmul12_fa1_3_y0 ^ f_u_arrmul12_fa1_3_f_u_arrmul12_ha0_3_y1;
  assign f_u_arrmul12_fa1_3_y3 = f_u_arrmul12_fa1_3_y0 & f_u_arrmul12_fa1_3_f_u_arrmul12_ha0_3_y1;
  assign f_u_arrmul12_fa1_3_y4 = f_u_arrmul12_fa1_3_y1 | f_u_arrmul12_fa1_3_y3;
  assign f_u_arrmul12_and2_3_a_2 = a_2;
  assign f_u_arrmul12_and2_3_b_3 = b_3;
  assign f_u_arrmul12_and2_3_y0 = f_u_arrmul12_and2_3_a_2 & f_u_arrmul12_and2_3_b_3;
  assign f_u_arrmul12_fa2_3_f_u_arrmul12_and2_3_y0 = f_u_arrmul12_and2_3_y0;
  assign f_u_arrmul12_fa2_3_f_u_arrmul12_fa3_2_y2 = f_u_arrmul12_fa3_2_y2;
  assign f_u_arrmul12_fa2_3_f_u_arrmul12_fa1_3_y4 = f_u_arrmul12_fa1_3_y4;
  assign f_u_arrmul12_fa2_3_y0 = f_u_arrmul12_fa2_3_f_u_arrmul12_and2_3_y0 ^ f_u_arrmul12_fa2_3_f_u_arrmul12_fa3_2_y2;
  assign f_u_arrmul12_fa2_3_y1 = f_u_arrmul12_fa2_3_f_u_arrmul12_and2_3_y0 & f_u_arrmul12_fa2_3_f_u_arrmul12_fa3_2_y2;
  assign f_u_arrmul12_fa2_3_y2 = f_u_arrmul12_fa2_3_y0 ^ f_u_arrmul12_fa2_3_f_u_arrmul12_fa1_3_y4;
  assign f_u_arrmul12_fa2_3_y3 = f_u_arrmul12_fa2_3_y0 & f_u_arrmul12_fa2_3_f_u_arrmul12_fa1_3_y4;
  assign f_u_arrmul12_fa2_3_y4 = f_u_arrmul12_fa2_3_y1 | f_u_arrmul12_fa2_3_y3;
  assign f_u_arrmul12_and3_3_a_3 = a_3;
  assign f_u_arrmul12_and3_3_b_3 = b_3;
  assign f_u_arrmul12_and3_3_y0 = f_u_arrmul12_and3_3_a_3 & f_u_arrmul12_and3_3_b_3;
  assign f_u_arrmul12_fa3_3_f_u_arrmul12_and3_3_y0 = f_u_arrmul12_and3_3_y0;
  assign f_u_arrmul12_fa3_3_f_u_arrmul12_fa4_2_y2 = f_u_arrmul12_fa4_2_y2;
  assign f_u_arrmul12_fa3_3_f_u_arrmul12_fa2_3_y4 = f_u_arrmul12_fa2_3_y4;
  assign f_u_arrmul12_fa3_3_y0 = f_u_arrmul12_fa3_3_f_u_arrmul12_and3_3_y0 ^ f_u_arrmul12_fa3_3_f_u_arrmul12_fa4_2_y2;
  assign f_u_arrmul12_fa3_3_y1 = f_u_arrmul12_fa3_3_f_u_arrmul12_and3_3_y0 & f_u_arrmul12_fa3_3_f_u_arrmul12_fa4_2_y2;
  assign f_u_arrmul12_fa3_3_y2 = f_u_arrmul12_fa3_3_y0 ^ f_u_arrmul12_fa3_3_f_u_arrmul12_fa2_3_y4;
  assign f_u_arrmul12_fa3_3_y3 = f_u_arrmul12_fa3_3_y0 & f_u_arrmul12_fa3_3_f_u_arrmul12_fa2_3_y4;
  assign f_u_arrmul12_fa3_3_y4 = f_u_arrmul12_fa3_3_y1 | f_u_arrmul12_fa3_3_y3;
  assign f_u_arrmul12_and4_3_a_4 = a_4;
  assign f_u_arrmul12_and4_3_b_3 = b_3;
  assign f_u_arrmul12_and4_3_y0 = f_u_arrmul12_and4_3_a_4 & f_u_arrmul12_and4_3_b_3;
  assign f_u_arrmul12_fa4_3_f_u_arrmul12_and4_3_y0 = f_u_arrmul12_and4_3_y0;
  assign f_u_arrmul12_fa4_3_f_u_arrmul12_fa5_2_y2 = f_u_arrmul12_fa5_2_y2;
  assign f_u_arrmul12_fa4_3_f_u_arrmul12_fa3_3_y4 = f_u_arrmul12_fa3_3_y4;
  assign f_u_arrmul12_fa4_3_y0 = f_u_arrmul12_fa4_3_f_u_arrmul12_and4_3_y0 ^ f_u_arrmul12_fa4_3_f_u_arrmul12_fa5_2_y2;
  assign f_u_arrmul12_fa4_3_y1 = f_u_arrmul12_fa4_3_f_u_arrmul12_and4_3_y0 & f_u_arrmul12_fa4_3_f_u_arrmul12_fa5_2_y2;
  assign f_u_arrmul12_fa4_3_y2 = f_u_arrmul12_fa4_3_y0 ^ f_u_arrmul12_fa4_3_f_u_arrmul12_fa3_3_y4;
  assign f_u_arrmul12_fa4_3_y3 = f_u_arrmul12_fa4_3_y0 & f_u_arrmul12_fa4_3_f_u_arrmul12_fa3_3_y4;
  assign f_u_arrmul12_fa4_3_y4 = f_u_arrmul12_fa4_3_y1 | f_u_arrmul12_fa4_3_y3;
  assign f_u_arrmul12_and5_3_a_5 = a_5;
  assign f_u_arrmul12_and5_3_b_3 = b_3;
  assign f_u_arrmul12_and5_3_y0 = f_u_arrmul12_and5_3_a_5 & f_u_arrmul12_and5_3_b_3;
  assign f_u_arrmul12_fa5_3_f_u_arrmul12_and5_3_y0 = f_u_arrmul12_and5_3_y0;
  assign f_u_arrmul12_fa5_3_f_u_arrmul12_fa6_2_y2 = f_u_arrmul12_fa6_2_y2;
  assign f_u_arrmul12_fa5_3_f_u_arrmul12_fa4_3_y4 = f_u_arrmul12_fa4_3_y4;
  assign f_u_arrmul12_fa5_3_y0 = f_u_arrmul12_fa5_3_f_u_arrmul12_and5_3_y0 ^ f_u_arrmul12_fa5_3_f_u_arrmul12_fa6_2_y2;
  assign f_u_arrmul12_fa5_3_y1 = f_u_arrmul12_fa5_3_f_u_arrmul12_and5_3_y0 & f_u_arrmul12_fa5_3_f_u_arrmul12_fa6_2_y2;
  assign f_u_arrmul12_fa5_3_y2 = f_u_arrmul12_fa5_3_y0 ^ f_u_arrmul12_fa5_3_f_u_arrmul12_fa4_3_y4;
  assign f_u_arrmul12_fa5_3_y3 = f_u_arrmul12_fa5_3_y0 & f_u_arrmul12_fa5_3_f_u_arrmul12_fa4_3_y4;
  assign f_u_arrmul12_fa5_3_y4 = f_u_arrmul12_fa5_3_y1 | f_u_arrmul12_fa5_3_y3;
  assign f_u_arrmul12_and6_3_a_6 = a_6;
  assign f_u_arrmul12_and6_3_b_3 = b_3;
  assign f_u_arrmul12_and6_3_y0 = f_u_arrmul12_and6_3_a_6 & f_u_arrmul12_and6_3_b_3;
  assign f_u_arrmul12_fa6_3_f_u_arrmul12_and6_3_y0 = f_u_arrmul12_and6_3_y0;
  assign f_u_arrmul12_fa6_3_f_u_arrmul12_fa7_2_y2 = f_u_arrmul12_fa7_2_y2;
  assign f_u_arrmul12_fa6_3_f_u_arrmul12_fa5_3_y4 = f_u_arrmul12_fa5_3_y4;
  assign f_u_arrmul12_fa6_3_y0 = f_u_arrmul12_fa6_3_f_u_arrmul12_and6_3_y0 ^ f_u_arrmul12_fa6_3_f_u_arrmul12_fa7_2_y2;
  assign f_u_arrmul12_fa6_3_y1 = f_u_arrmul12_fa6_3_f_u_arrmul12_and6_3_y0 & f_u_arrmul12_fa6_3_f_u_arrmul12_fa7_2_y2;
  assign f_u_arrmul12_fa6_3_y2 = f_u_arrmul12_fa6_3_y0 ^ f_u_arrmul12_fa6_3_f_u_arrmul12_fa5_3_y4;
  assign f_u_arrmul12_fa6_3_y3 = f_u_arrmul12_fa6_3_y0 & f_u_arrmul12_fa6_3_f_u_arrmul12_fa5_3_y4;
  assign f_u_arrmul12_fa6_3_y4 = f_u_arrmul12_fa6_3_y1 | f_u_arrmul12_fa6_3_y3;
  assign f_u_arrmul12_and7_3_a_7 = a_7;
  assign f_u_arrmul12_and7_3_b_3 = b_3;
  assign f_u_arrmul12_and7_3_y0 = f_u_arrmul12_and7_3_a_7 & f_u_arrmul12_and7_3_b_3;
  assign f_u_arrmul12_fa7_3_f_u_arrmul12_and7_3_y0 = f_u_arrmul12_and7_3_y0;
  assign f_u_arrmul12_fa7_3_f_u_arrmul12_fa8_2_y2 = f_u_arrmul12_fa8_2_y2;
  assign f_u_arrmul12_fa7_3_f_u_arrmul12_fa6_3_y4 = f_u_arrmul12_fa6_3_y4;
  assign f_u_arrmul12_fa7_3_y0 = f_u_arrmul12_fa7_3_f_u_arrmul12_and7_3_y0 ^ f_u_arrmul12_fa7_3_f_u_arrmul12_fa8_2_y2;
  assign f_u_arrmul12_fa7_3_y1 = f_u_arrmul12_fa7_3_f_u_arrmul12_and7_3_y0 & f_u_arrmul12_fa7_3_f_u_arrmul12_fa8_2_y2;
  assign f_u_arrmul12_fa7_3_y2 = f_u_arrmul12_fa7_3_y0 ^ f_u_arrmul12_fa7_3_f_u_arrmul12_fa6_3_y4;
  assign f_u_arrmul12_fa7_3_y3 = f_u_arrmul12_fa7_3_y0 & f_u_arrmul12_fa7_3_f_u_arrmul12_fa6_3_y4;
  assign f_u_arrmul12_fa7_3_y4 = f_u_arrmul12_fa7_3_y1 | f_u_arrmul12_fa7_3_y3;
  assign f_u_arrmul12_and8_3_a_8 = a_8;
  assign f_u_arrmul12_and8_3_b_3 = b_3;
  assign f_u_arrmul12_and8_3_y0 = f_u_arrmul12_and8_3_a_8 & f_u_arrmul12_and8_3_b_3;
  assign f_u_arrmul12_fa8_3_f_u_arrmul12_and8_3_y0 = f_u_arrmul12_and8_3_y0;
  assign f_u_arrmul12_fa8_3_f_u_arrmul12_fa9_2_y2 = f_u_arrmul12_fa9_2_y2;
  assign f_u_arrmul12_fa8_3_f_u_arrmul12_fa7_3_y4 = f_u_arrmul12_fa7_3_y4;
  assign f_u_arrmul12_fa8_3_y0 = f_u_arrmul12_fa8_3_f_u_arrmul12_and8_3_y0 ^ f_u_arrmul12_fa8_3_f_u_arrmul12_fa9_2_y2;
  assign f_u_arrmul12_fa8_3_y1 = f_u_arrmul12_fa8_3_f_u_arrmul12_and8_3_y0 & f_u_arrmul12_fa8_3_f_u_arrmul12_fa9_2_y2;
  assign f_u_arrmul12_fa8_3_y2 = f_u_arrmul12_fa8_3_y0 ^ f_u_arrmul12_fa8_3_f_u_arrmul12_fa7_3_y4;
  assign f_u_arrmul12_fa8_3_y3 = f_u_arrmul12_fa8_3_y0 & f_u_arrmul12_fa8_3_f_u_arrmul12_fa7_3_y4;
  assign f_u_arrmul12_fa8_3_y4 = f_u_arrmul12_fa8_3_y1 | f_u_arrmul12_fa8_3_y3;
  assign f_u_arrmul12_and9_3_a_9 = a_9;
  assign f_u_arrmul12_and9_3_b_3 = b_3;
  assign f_u_arrmul12_and9_3_y0 = f_u_arrmul12_and9_3_a_9 & f_u_arrmul12_and9_3_b_3;
  assign f_u_arrmul12_fa9_3_f_u_arrmul12_and9_3_y0 = f_u_arrmul12_and9_3_y0;
  assign f_u_arrmul12_fa9_3_f_u_arrmul12_fa10_2_y2 = f_u_arrmul12_fa10_2_y2;
  assign f_u_arrmul12_fa9_3_f_u_arrmul12_fa8_3_y4 = f_u_arrmul12_fa8_3_y4;
  assign f_u_arrmul12_fa9_3_y0 = f_u_arrmul12_fa9_3_f_u_arrmul12_and9_3_y0 ^ f_u_arrmul12_fa9_3_f_u_arrmul12_fa10_2_y2;
  assign f_u_arrmul12_fa9_3_y1 = f_u_arrmul12_fa9_3_f_u_arrmul12_and9_3_y0 & f_u_arrmul12_fa9_3_f_u_arrmul12_fa10_2_y2;
  assign f_u_arrmul12_fa9_3_y2 = f_u_arrmul12_fa9_3_y0 ^ f_u_arrmul12_fa9_3_f_u_arrmul12_fa8_3_y4;
  assign f_u_arrmul12_fa9_3_y3 = f_u_arrmul12_fa9_3_y0 & f_u_arrmul12_fa9_3_f_u_arrmul12_fa8_3_y4;
  assign f_u_arrmul12_fa9_3_y4 = f_u_arrmul12_fa9_3_y1 | f_u_arrmul12_fa9_3_y3;
  assign f_u_arrmul12_and10_3_a_10 = a_10;
  assign f_u_arrmul12_and10_3_b_3 = b_3;
  assign f_u_arrmul12_and10_3_y0 = f_u_arrmul12_and10_3_a_10 & f_u_arrmul12_and10_3_b_3;
  assign f_u_arrmul12_fa10_3_f_u_arrmul12_and10_3_y0 = f_u_arrmul12_and10_3_y0;
  assign f_u_arrmul12_fa10_3_f_u_arrmul12_fa11_2_y2 = f_u_arrmul12_fa11_2_y2;
  assign f_u_arrmul12_fa10_3_f_u_arrmul12_fa9_3_y4 = f_u_arrmul12_fa9_3_y4;
  assign f_u_arrmul12_fa10_3_y0 = f_u_arrmul12_fa10_3_f_u_arrmul12_and10_3_y0 ^ f_u_arrmul12_fa10_3_f_u_arrmul12_fa11_2_y2;
  assign f_u_arrmul12_fa10_3_y1 = f_u_arrmul12_fa10_3_f_u_arrmul12_and10_3_y0 & f_u_arrmul12_fa10_3_f_u_arrmul12_fa11_2_y2;
  assign f_u_arrmul12_fa10_3_y2 = f_u_arrmul12_fa10_3_y0 ^ f_u_arrmul12_fa10_3_f_u_arrmul12_fa9_3_y4;
  assign f_u_arrmul12_fa10_3_y3 = f_u_arrmul12_fa10_3_y0 & f_u_arrmul12_fa10_3_f_u_arrmul12_fa9_3_y4;
  assign f_u_arrmul12_fa10_3_y4 = f_u_arrmul12_fa10_3_y1 | f_u_arrmul12_fa10_3_y3;
  assign f_u_arrmul12_and11_3_a_11 = a_11;
  assign f_u_arrmul12_and11_3_b_3 = b_3;
  assign f_u_arrmul12_and11_3_y0 = f_u_arrmul12_and11_3_a_11 & f_u_arrmul12_and11_3_b_3;
  assign f_u_arrmul12_fa11_3_f_u_arrmul12_and11_3_y0 = f_u_arrmul12_and11_3_y0;
  assign f_u_arrmul12_fa11_3_f_u_arrmul12_fa11_2_y4 = f_u_arrmul12_fa11_2_y4;
  assign f_u_arrmul12_fa11_3_f_u_arrmul12_fa10_3_y4 = f_u_arrmul12_fa10_3_y4;
  assign f_u_arrmul12_fa11_3_y0 = f_u_arrmul12_fa11_3_f_u_arrmul12_and11_3_y0 ^ f_u_arrmul12_fa11_3_f_u_arrmul12_fa11_2_y4;
  assign f_u_arrmul12_fa11_3_y1 = f_u_arrmul12_fa11_3_f_u_arrmul12_and11_3_y0 & f_u_arrmul12_fa11_3_f_u_arrmul12_fa11_2_y4;
  assign f_u_arrmul12_fa11_3_y2 = f_u_arrmul12_fa11_3_y0 ^ f_u_arrmul12_fa11_3_f_u_arrmul12_fa10_3_y4;
  assign f_u_arrmul12_fa11_3_y3 = f_u_arrmul12_fa11_3_y0 & f_u_arrmul12_fa11_3_f_u_arrmul12_fa10_3_y4;
  assign f_u_arrmul12_fa11_3_y4 = f_u_arrmul12_fa11_3_y1 | f_u_arrmul12_fa11_3_y3;
  assign f_u_arrmul12_and0_4_a_0 = a_0;
  assign f_u_arrmul12_and0_4_b_4 = b_4;
  assign f_u_arrmul12_and0_4_y0 = f_u_arrmul12_and0_4_a_0 & f_u_arrmul12_and0_4_b_4;
  assign f_u_arrmul12_ha0_4_f_u_arrmul12_and0_4_y0 = f_u_arrmul12_and0_4_y0;
  assign f_u_arrmul12_ha0_4_f_u_arrmul12_fa1_3_y2 = f_u_arrmul12_fa1_3_y2;
  assign f_u_arrmul12_ha0_4_y0 = f_u_arrmul12_ha0_4_f_u_arrmul12_and0_4_y0 ^ f_u_arrmul12_ha0_4_f_u_arrmul12_fa1_3_y2;
  assign f_u_arrmul12_ha0_4_y1 = f_u_arrmul12_ha0_4_f_u_arrmul12_and0_4_y0 & f_u_arrmul12_ha0_4_f_u_arrmul12_fa1_3_y2;
  assign f_u_arrmul12_and1_4_a_1 = a_1;
  assign f_u_arrmul12_and1_4_b_4 = b_4;
  assign f_u_arrmul12_and1_4_y0 = f_u_arrmul12_and1_4_a_1 & f_u_arrmul12_and1_4_b_4;
  assign f_u_arrmul12_fa1_4_f_u_arrmul12_and1_4_y0 = f_u_arrmul12_and1_4_y0;
  assign f_u_arrmul12_fa1_4_f_u_arrmul12_fa2_3_y2 = f_u_arrmul12_fa2_3_y2;
  assign f_u_arrmul12_fa1_4_f_u_arrmul12_ha0_4_y1 = f_u_arrmul12_ha0_4_y1;
  assign f_u_arrmul12_fa1_4_y0 = f_u_arrmul12_fa1_4_f_u_arrmul12_and1_4_y0 ^ f_u_arrmul12_fa1_4_f_u_arrmul12_fa2_3_y2;
  assign f_u_arrmul12_fa1_4_y1 = f_u_arrmul12_fa1_4_f_u_arrmul12_and1_4_y0 & f_u_arrmul12_fa1_4_f_u_arrmul12_fa2_3_y2;
  assign f_u_arrmul12_fa1_4_y2 = f_u_arrmul12_fa1_4_y0 ^ f_u_arrmul12_fa1_4_f_u_arrmul12_ha0_4_y1;
  assign f_u_arrmul12_fa1_4_y3 = f_u_arrmul12_fa1_4_y0 & f_u_arrmul12_fa1_4_f_u_arrmul12_ha0_4_y1;
  assign f_u_arrmul12_fa1_4_y4 = f_u_arrmul12_fa1_4_y1 | f_u_arrmul12_fa1_4_y3;
  assign f_u_arrmul12_and2_4_a_2 = a_2;
  assign f_u_arrmul12_and2_4_b_4 = b_4;
  assign f_u_arrmul12_and2_4_y0 = f_u_arrmul12_and2_4_a_2 & f_u_arrmul12_and2_4_b_4;
  assign f_u_arrmul12_fa2_4_f_u_arrmul12_and2_4_y0 = f_u_arrmul12_and2_4_y0;
  assign f_u_arrmul12_fa2_4_f_u_arrmul12_fa3_3_y2 = f_u_arrmul12_fa3_3_y2;
  assign f_u_arrmul12_fa2_4_f_u_arrmul12_fa1_4_y4 = f_u_arrmul12_fa1_4_y4;
  assign f_u_arrmul12_fa2_4_y0 = f_u_arrmul12_fa2_4_f_u_arrmul12_and2_4_y0 ^ f_u_arrmul12_fa2_4_f_u_arrmul12_fa3_3_y2;
  assign f_u_arrmul12_fa2_4_y1 = f_u_arrmul12_fa2_4_f_u_arrmul12_and2_4_y0 & f_u_arrmul12_fa2_4_f_u_arrmul12_fa3_3_y2;
  assign f_u_arrmul12_fa2_4_y2 = f_u_arrmul12_fa2_4_y0 ^ f_u_arrmul12_fa2_4_f_u_arrmul12_fa1_4_y4;
  assign f_u_arrmul12_fa2_4_y3 = f_u_arrmul12_fa2_4_y0 & f_u_arrmul12_fa2_4_f_u_arrmul12_fa1_4_y4;
  assign f_u_arrmul12_fa2_4_y4 = f_u_arrmul12_fa2_4_y1 | f_u_arrmul12_fa2_4_y3;
  assign f_u_arrmul12_and3_4_a_3 = a_3;
  assign f_u_arrmul12_and3_4_b_4 = b_4;
  assign f_u_arrmul12_and3_4_y0 = f_u_arrmul12_and3_4_a_3 & f_u_arrmul12_and3_4_b_4;
  assign f_u_arrmul12_fa3_4_f_u_arrmul12_and3_4_y0 = f_u_arrmul12_and3_4_y0;
  assign f_u_arrmul12_fa3_4_f_u_arrmul12_fa4_3_y2 = f_u_arrmul12_fa4_3_y2;
  assign f_u_arrmul12_fa3_4_f_u_arrmul12_fa2_4_y4 = f_u_arrmul12_fa2_4_y4;
  assign f_u_arrmul12_fa3_4_y0 = f_u_arrmul12_fa3_4_f_u_arrmul12_and3_4_y0 ^ f_u_arrmul12_fa3_4_f_u_arrmul12_fa4_3_y2;
  assign f_u_arrmul12_fa3_4_y1 = f_u_arrmul12_fa3_4_f_u_arrmul12_and3_4_y0 & f_u_arrmul12_fa3_4_f_u_arrmul12_fa4_3_y2;
  assign f_u_arrmul12_fa3_4_y2 = f_u_arrmul12_fa3_4_y0 ^ f_u_arrmul12_fa3_4_f_u_arrmul12_fa2_4_y4;
  assign f_u_arrmul12_fa3_4_y3 = f_u_arrmul12_fa3_4_y0 & f_u_arrmul12_fa3_4_f_u_arrmul12_fa2_4_y4;
  assign f_u_arrmul12_fa3_4_y4 = f_u_arrmul12_fa3_4_y1 | f_u_arrmul12_fa3_4_y3;
  assign f_u_arrmul12_and4_4_a_4 = a_4;
  assign f_u_arrmul12_and4_4_b_4 = b_4;
  assign f_u_arrmul12_and4_4_y0 = f_u_arrmul12_and4_4_a_4 & f_u_arrmul12_and4_4_b_4;
  assign f_u_arrmul12_fa4_4_f_u_arrmul12_and4_4_y0 = f_u_arrmul12_and4_4_y0;
  assign f_u_arrmul12_fa4_4_f_u_arrmul12_fa5_3_y2 = f_u_arrmul12_fa5_3_y2;
  assign f_u_arrmul12_fa4_4_f_u_arrmul12_fa3_4_y4 = f_u_arrmul12_fa3_4_y4;
  assign f_u_arrmul12_fa4_4_y0 = f_u_arrmul12_fa4_4_f_u_arrmul12_and4_4_y0 ^ f_u_arrmul12_fa4_4_f_u_arrmul12_fa5_3_y2;
  assign f_u_arrmul12_fa4_4_y1 = f_u_arrmul12_fa4_4_f_u_arrmul12_and4_4_y0 & f_u_arrmul12_fa4_4_f_u_arrmul12_fa5_3_y2;
  assign f_u_arrmul12_fa4_4_y2 = f_u_arrmul12_fa4_4_y0 ^ f_u_arrmul12_fa4_4_f_u_arrmul12_fa3_4_y4;
  assign f_u_arrmul12_fa4_4_y3 = f_u_arrmul12_fa4_4_y0 & f_u_arrmul12_fa4_4_f_u_arrmul12_fa3_4_y4;
  assign f_u_arrmul12_fa4_4_y4 = f_u_arrmul12_fa4_4_y1 | f_u_arrmul12_fa4_4_y3;
  assign f_u_arrmul12_and5_4_a_5 = a_5;
  assign f_u_arrmul12_and5_4_b_4 = b_4;
  assign f_u_arrmul12_and5_4_y0 = f_u_arrmul12_and5_4_a_5 & f_u_arrmul12_and5_4_b_4;
  assign f_u_arrmul12_fa5_4_f_u_arrmul12_and5_4_y0 = f_u_arrmul12_and5_4_y0;
  assign f_u_arrmul12_fa5_4_f_u_arrmul12_fa6_3_y2 = f_u_arrmul12_fa6_3_y2;
  assign f_u_arrmul12_fa5_4_f_u_arrmul12_fa4_4_y4 = f_u_arrmul12_fa4_4_y4;
  assign f_u_arrmul12_fa5_4_y0 = f_u_arrmul12_fa5_4_f_u_arrmul12_and5_4_y0 ^ f_u_arrmul12_fa5_4_f_u_arrmul12_fa6_3_y2;
  assign f_u_arrmul12_fa5_4_y1 = f_u_arrmul12_fa5_4_f_u_arrmul12_and5_4_y0 & f_u_arrmul12_fa5_4_f_u_arrmul12_fa6_3_y2;
  assign f_u_arrmul12_fa5_4_y2 = f_u_arrmul12_fa5_4_y0 ^ f_u_arrmul12_fa5_4_f_u_arrmul12_fa4_4_y4;
  assign f_u_arrmul12_fa5_4_y3 = f_u_arrmul12_fa5_4_y0 & f_u_arrmul12_fa5_4_f_u_arrmul12_fa4_4_y4;
  assign f_u_arrmul12_fa5_4_y4 = f_u_arrmul12_fa5_4_y1 | f_u_arrmul12_fa5_4_y3;
  assign f_u_arrmul12_and6_4_a_6 = a_6;
  assign f_u_arrmul12_and6_4_b_4 = b_4;
  assign f_u_arrmul12_and6_4_y0 = f_u_arrmul12_and6_4_a_6 & f_u_arrmul12_and6_4_b_4;
  assign f_u_arrmul12_fa6_4_f_u_arrmul12_and6_4_y0 = f_u_arrmul12_and6_4_y0;
  assign f_u_arrmul12_fa6_4_f_u_arrmul12_fa7_3_y2 = f_u_arrmul12_fa7_3_y2;
  assign f_u_arrmul12_fa6_4_f_u_arrmul12_fa5_4_y4 = f_u_arrmul12_fa5_4_y4;
  assign f_u_arrmul12_fa6_4_y0 = f_u_arrmul12_fa6_4_f_u_arrmul12_and6_4_y0 ^ f_u_arrmul12_fa6_4_f_u_arrmul12_fa7_3_y2;
  assign f_u_arrmul12_fa6_4_y1 = f_u_arrmul12_fa6_4_f_u_arrmul12_and6_4_y0 & f_u_arrmul12_fa6_4_f_u_arrmul12_fa7_3_y2;
  assign f_u_arrmul12_fa6_4_y2 = f_u_arrmul12_fa6_4_y0 ^ f_u_arrmul12_fa6_4_f_u_arrmul12_fa5_4_y4;
  assign f_u_arrmul12_fa6_4_y3 = f_u_arrmul12_fa6_4_y0 & f_u_arrmul12_fa6_4_f_u_arrmul12_fa5_4_y4;
  assign f_u_arrmul12_fa6_4_y4 = f_u_arrmul12_fa6_4_y1 | f_u_arrmul12_fa6_4_y3;
  assign f_u_arrmul12_and7_4_a_7 = a_7;
  assign f_u_arrmul12_and7_4_b_4 = b_4;
  assign f_u_arrmul12_and7_4_y0 = f_u_arrmul12_and7_4_a_7 & f_u_arrmul12_and7_4_b_4;
  assign f_u_arrmul12_fa7_4_f_u_arrmul12_and7_4_y0 = f_u_arrmul12_and7_4_y0;
  assign f_u_arrmul12_fa7_4_f_u_arrmul12_fa8_3_y2 = f_u_arrmul12_fa8_3_y2;
  assign f_u_arrmul12_fa7_4_f_u_arrmul12_fa6_4_y4 = f_u_arrmul12_fa6_4_y4;
  assign f_u_arrmul12_fa7_4_y0 = f_u_arrmul12_fa7_4_f_u_arrmul12_and7_4_y0 ^ f_u_arrmul12_fa7_4_f_u_arrmul12_fa8_3_y2;
  assign f_u_arrmul12_fa7_4_y1 = f_u_arrmul12_fa7_4_f_u_arrmul12_and7_4_y0 & f_u_arrmul12_fa7_4_f_u_arrmul12_fa8_3_y2;
  assign f_u_arrmul12_fa7_4_y2 = f_u_arrmul12_fa7_4_y0 ^ f_u_arrmul12_fa7_4_f_u_arrmul12_fa6_4_y4;
  assign f_u_arrmul12_fa7_4_y3 = f_u_arrmul12_fa7_4_y0 & f_u_arrmul12_fa7_4_f_u_arrmul12_fa6_4_y4;
  assign f_u_arrmul12_fa7_4_y4 = f_u_arrmul12_fa7_4_y1 | f_u_arrmul12_fa7_4_y3;
  assign f_u_arrmul12_and8_4_a_8 = a_8;
  assign f_u_arrmul12_and8_4_b_4 = b_4;
  assign f_u_arrmul12_and8_4_y0 = f_u_arrmul12_and8_4_a_8 & f_u_arrmul12_and8_4_b_4;
  assign f_u_arrmul12_fa8_4_f_u_arrmul12_and8_4_y0 = f_u_arrmul12_and8_4_y0;
  assign f_u_arrmul12_fa8_4_f_u_arrmul12_fa9_3_y2 = f_u_arrmul12_fa9_3_y2;
  assign f_u_arrmul12_fa8_4_f_u_arrmul12_fa7_4_y4 = f_u_arrmul12_fa7_4_y4;
  assign f_u_arrmul12_fa8_4_y0 = f_u_arrmul12_fa8_4_f_u_arrmul12_and8_4_y0 ^ f_u_arrmul12_fa8_4_f_u_arrmul12_fa9_3_y2;
  assign f_u_arrmul12_fa8_4_y1 = f_u_arrmul12_fa8_4_f_u_arrmul12_and8_4_y0 & f_u_arrmul12_fa8_4_f_u_arrmul12_fa9_3_y2;
  assign f_u_arrmul12_fa8_4_y2 = f_u_arrmul12_fa8_4_y0 ^ f_u_arrmul12_fa8_4_f_u_arrmul12_fa7_4_y4;
  assign f_u_arrmul12_fa8_4_y3 = f_u_arrmul12_fa8_4_y0 & f_u_arrmul12_fa8_4_f_u_arrmul12_fa7_4_y4;
  assign f_u_arrmul12_fa8_4_y4 = f_u_arrmul12_fa8_4_y1 | f_u_arrmul12_fa8_4_y3;
  assign f_u_arrmul12_and9_4_a_9 = a_9;
  assign f_u_arrmul12_and9_4_b_4 = b_4;
  assign f_u_arrmul12_and9_4_y0 = f_u_arrmul12_and9_4_a_9 & f_u_arrmul12_and9_4_b_4;
  assign f_u_arrmul12_fa9_4_f_u_arrmul12_and9_4_y0 = f_u_arrmul12_and9_4_y0;
  assign f_u_arrmul12_fa9_4_f_u_arrmul12_fa10_3_y2 = f_u_arrmul12_fa10_3_y2;
  assign f_u_arrmul12_fa9_4_f_u_arrmul12_fa8_4_y4 = f_u_arrmul12_fa8_4_y4;
  assign f_u_arrmul12_fa9_4_y0 = f_u_arrmul12_fa9_4_f_u_arrmul12_and9_4_y0 ^ f_u_arrmul12_fa9_4_f_u_arrmul12_fa10_3_y2;
  assign f_u_arrmul12_fa9_4_y1 = f_u_arrmul12_fa9_4_f_u_arrmul12_and9_4_y0 & f_u_arrmul12_fa9_4_f_u_arrmul12_fa10_3_y2;
  assign f_u_arrmul12_fa9_4_y2 = f_u_arrmul12_fa9_4_y0 ^ f_u_arrmul12_fa9_4_f_u_arrmul12_fa8_4_y4;
  assign f_u_arrmul12_fa9_4_y3 = f_u_arrmul12_fa9_4_y0 & f_u_arrmul12_fa9_4_f_u_arrmul12_fa8_4_y4;
  assign f_u_arrmul12_fa9_4_y4 = f_u_arrmul12_fa9_4_y1 | f_u_arrmul12_fa9_4_y3;
  assign f_u_arrmul12_and10_4_a_10 = a_10;
  assign f_u_arrmul12_and10_4_b_4 = b_4;
  assign f_u_arrmul12_and10_4_y0 = f_u_arrmul12_and10_4_a_10 & f_u_arrmul12_and10_4_b_4;
  assign f_u_arrmul12_fa10_4_f_u_arrmul12_and10_4_y0 = f_u_arrmul12_and10_4_y0;
  assign f_u_arrmul12_fa10_4_f_u_arrmul12_fa11_3_y2 = f_u_arrmul12_fa11_3_y2;
  assign f_u_arrmul12_fa10_4_f_u_arrmul12_fa9_4_y4 = f_u_arrmul12_fa9_4_y4;
  assign f_u_arrmul12_fa10_4_y0 = f_u_arrmul12_fa10_4_f_u_arrmul12_and10_4_y0 ^ f_u_arrmul12_fa10_4_f_u_arrmul12_fa11_3_y2;
  assign f_u_arrmul12_fa10_4_y1 = f_u_arrmul12_fa10_4_f_u_arrmul12_and10_4_y0 & f_u_arrmul12_fa10_4_f_u_arrmul12_fa11_3_y2;
  assign f_u_arrmul12_fa10_4_y2 = f_u_arrmul12_fa10_4_y0 ^ f_u_arrmul12_fa10_4_f_u_arrmul12_fa9_4_y4;
  assign f_u_arrmul12_fa10_4_y3 = f_u_arrmul12_fa10_4_y0 & f_u_arrmul12_fa10_4_f_u_arrmul12_fa9_4_y4;
  assign f_u_arrmul12_fa10_4_y4 = f_u_arrmul12_fa10_4_y1 | f_u_arrmul12_fa10_4_y3;
  assign f_u_arrmul12_and11_4_a_11 = a_11;
  assign f_u_arrmul12_and11_4_b_4 = b_4;
  assign f_u_arrmul12_and11_4_y0 = f_u_arrmul12_and11_4_a_11 & f_u_arrmul12_and11_4_b_4;
  assign f_u_arrmul12_fa11_4_f_u_arrmul12_and11_4_y0 = f_u_arrmul12_and11_4_y0;
  assign f_u_arrmul12_fa11_4_f_u_arrmul12_fa11_3_y4 = f_u_arrmul12_fa11_3_y4;
  assign f_u_arrmul12_fa11_4_f_u_arrmul12_fa10_4_y4 = f_u_arrmul12_fa10_4_y4;
  assign f_u_arrmul12_fa11_4_y0 = f_u_arrmul12_fa11_4_f_u_arrmul12_and11_4_y0 ^ f_u_arrmul12_fa11_4_f_u_arrmul12_fa11_3_y4;
  assign f_u_arrmul12_fa11_4_y1 = f_u_arrmul12_fa11_4_f_u_arrmul12_and11_4_y0 & f_u_arrmul12_fa11_4_f_u_arrmul12_fa11_3_y4;
  assign f_u_arrmul12_fa11_4_y2 = f_u_arrmul12_fa11_4_y0 ^ f_u_arrmul12_fa11_4_f_u_arrmul12_fa10_4_y4;
  assign f_u_arrmul12_fa11_4_y3 = f_u_arrmul12_fa11_4_y0 & f_u_arrmul12_fa11_4_f_u_arrmul12_fa10_4_y4;
  assign f_u_arrmul12_fa11_4_y4 = f_u_arrmul12_fa11_4_y1 | f_u_arrmul12_fa11_4_y3;
  assign f_u_arrmul12_and0_5_a_0 = a_0;
  assign f_u_arrmul12_and0_5_b_5 = b_5;
  assign f_u_arrmul12_and0_5_y0 = f_u_arrmul12_and0_5_a_0 & f_u_arrmul12_and0_5_b_5;
  assign f_u_arrmul12_ha0_5_f_u_arrmul12_and0_5_y0 = f_u_arrmul12_and0_5_y0;
  assign f_u_arrmul12_ha0_5_f_u_arrmul12_fa1_4_y2 = f_u_arrmul12_fa1_4_y2;
  assign f_u_arrmul12_ha0_5_y0 = f_u_arrmul12_ha0_5_f_u_arrmul12_and0_5_y0 ^ f_u_arrmul12_ha0_5_f_u_arrmul12_fa1_4_y2;
  assign f_u_arrmul12_ha0_5_y1 = f_u_arrmul12_ha0_5_f_u_arrmul12_and0_5_y0 & f_u_arrmul12_ha0_5_f_u_arrmul12_fa1_4_y2;
  assign f_u_arrmul12_and1_5_a_1 = a_1;
  assign f_u_arrmul12_and1_5_b_5 = b_5;
  assign f_u_arrmul12_and1_5_y0 = f_u_arrmul12_and1_5_a_1 & f_u_arrmul12_and1_5_b_5;
  assign f_u_arrmul12_fa1_5_f_u_arrmul12_and1_5_y0 = f_u_arrmul12_and1_5_y0;
  assign f_u_arrmul12_fa1_5_f_u_arrmul12_fa2_4_y2 = f_u_arrmul12_fa2_4_y2;
  assign f_u_arrmul12_fa1_5_f_u_arrmul12_ha0_5_y1 = f_u_arrmul12_ha0_5_y1;
  assign f_u_arrmul12_fa1_5_y0 = f_u_arrmul12_fa1_5_f_u_arrmul12_and1_5_y0 ^ f_u_arrmul12_fa1_5_f_u_arrmul12_fa2_4_y2;
  assign f_u_arrmul12_fa1_5_y1 = f_u_arrmul12_fa1_5_f_u_arrmul12_and1_5_y0 & f_u_arrmul12_fa1_5_f_u_arrmul12_fa2_4_y2;
  assign f_u_arrmul12_fa1_5_y2 = f_u_arrmul12_fa1_5_y0 ^ f_u_arrmul12_fa1_5_f_u_arrmul12_ha0_5_y1;
  assign f_u_arrmul12_fa1_5_y3 = f_u_arrmul12_fa1_5_y0 & f_u_arrmul12_fa1_5_f_u_arrmul12_ha0_5_y1;
  assign f_u_arrmul12_fa1_5_y4 = f_u_arrmul12_fa1_5_y1 | f_u_arrmul12_fa1_5_y3;
  assign f_u_arrmul12_and2_5_a_2 = a_2;
  assign f_u_arrmul12_and2_5_b_5 = b_5;
  assign f_u_arrmul12_and2_5_y0 = f_u_arrmul12_and2_5_a_2 & f_u_arrmul12_and2_5_b_5;
  assign f_u_arrmul12_fa2_5_f_u_arrmul12_and2_5_y0 = f_u_arrmul12_and2_5_y0;
  assign f_u_arrmul12_fa2_5_f_u_arrmul12_fa3_4_y2 = f_u_arrmul12_fa3_4_y2;
  assign f_u_arrmul12_fa2_5_f_u_arrmul12_fa1_5_y4 = f_u_arrmul12_fa1_5_y4;
  assign f_u_arrmul12_fa2_5_y0 = f_u_arrmul12_fa2_5_f_u_arrmul12_and2_5_y0 ^ f_u_arrmul12_fa2_5_f_u_arrmul12_fa3_4_y2;
  assign f_u_arrmul12_fa2_5_y1 = f_u_arrmul12_fa2_5_f_u_arrmul12_and2_5_y0 & f_u_arrmul12_fa2_5_f_u_arrmul12_fa3_4_y2;
  assign f_u_arrmul12_fa2_5_y2 = f_u_arrmul12_fa2_5_y0 ^ f_u_arrmul12_fa2_5_f_u_arrmul12_fa1_5_y4;
  assign f_u_arrmul12_fa2_5_y3 = f_u_arrmul12_fa2_5_y0 & f_u_arrmul12_fa2_5_f_u_arrmul12_fa1_5_y4;
  assign f_u_arrmul12_fa2_5_y4 = f_u_arrmul12_fa2_5_y1 | f_u_arrmul12_fa2_5_y3;
  assign f_u_arrmul12_and3_5_a_3 = a_3;
  assign f_u_arrmul12_and3_5_b_5 = b_5;
  assign f_u_arrmul12_and3_5_y0 = f_u_arrmul12_and3_5_a_3 & f_u_arrmul12_and3_5_b_5;
  assign f_u_arrmul12_fa3_5_f_u_arrmul12_and3_5_y0 = f_u_arrmul12_and3_5_y0;
  assign f_u_arrmul12_fa3_5_f_u_arrmul12_fa4_4_y2 = f_u_arrmul12_fa4_4_y2;
  assign f_u_arrmul12_fa3_5_f_u_arrmul12_fa2_5_y4 = f_u_arrmul12_fa2_5_y4;
  assign f_u_arrmul12_fa3_5_y0 = f_u_arrmul12_fa3_5_f_u_arrmul12_and3_5_y0 ^ f_u_arrmul12_fa3_5_f_u_arrmul12_fa4_4_y2;
  assign f_u_arrmul12_fa3_5_y1 = f_u_arrmul12_fa3_5_f_u_arrmul12_and3_5_y0 & f_u_arrmul12_fa3_5_f_u_arrmul12_fa4_4_y2;
  assign f_u_arrmul12_fa3_5_y2 = f_u_arrmul12_fa3_5_y0 ^ f_u_arrmul12_fa3_5_f_u_arrmul12_fa2_5_y4;
  assign f_u_arrmul12_fa3_5_y3 = f_u_arrmul12_fa3_5_y0 & f_u_arrmul12_fa3_5_f_u_arrmul12_fa2_5_y4;
  assign f_u_arrmul12_fa3_5_y4 = f_u_arrmul12_fa3_5_y1 | f_u_arrmul12_fa3_5_y3;
  assign f_u_arrmul12_and4_5_a_4 = a_4;
  assign f_u_arrmul12_and4_5_b_5 = b_5;
  assign f_u_arrmul12_and4_5_y0 = f_u_arrmul12_and4_5_a_4 & f_u_arrmul12_and4_5_b_5;
  assign f_u_arrmul12_fa4_5_f_u_arrmul12_and4_5_y0 = f_u_arrmul12_and4_5_y0;
  assign f_u_arrmul12_fa4_5_f_u_arrmul12_fa5_4_y2 = f_u_arrmul12_fa5_4_y2;
  assign f_u_arrmul12_fa4_5_f_u_arrmul12_fa3_5_y4 = f_u_arrmul12_fa3_5_y4;
  assign f_u_arrmul12_fa4_5_y0 = f_u_arrmul12_fa4_5_f_u_arrmul12_and4_5_y0 ^ f_u_arrmul12_fa4_5_f_u_arrmul12_fa5_4_y2;
  assign f_u_arrmul12_fa4_5_y1 = f_u_arrmul12_fa4_5_f_u_arrmul12_and4_5_y0 & f_u_arrmul12_fa4_5_f_u_arrmul12_fa5_4_y2;
  assign f_u_arrmul12_fa4_5_y2 = f_u_arrmul12_fa4_5_y0 ^ f_u_arrmul12_fa4_5_f_u_arrmul12_fa3_5_y4;
  assign f_u_arrmul12_fa4_5_y3 = f_u_arrmul12_fa4_5_y0 & f_u_arrmul12_fa4_5_f_u_arrmul12_fa3_5_y4;
  assign f_u_arrmul12_fa4_5_y4 = f_u_arrmul12_fa4_5_y1 | f_u_arrmul12_fa4_5_y3;
  assign f_u_arrmul12_and5_5_a_5 = a_5;
  assign f_u_arrmul12_and5_5_b_5 = b_5;
  assign f_u_arrmul12_and5_5_y0 = f_u_arrmul12_and5_5_a_5 & f_u_arrmul12_and5_5_b_5;
  assign f_u_arrmul12_fa5_5_f_u_arrmul12_and5_5_y0 = f_u_arrmul12_and5_5_y0;
  assign f_u_arrmul12_fa5_5_f_u_arrmul12_fa6_4_y2 = f_u_arrmul12_fa6_4_y2;
  assign f_u_arrmul12_fa5_5_f_u_arrmul12_fa4_5_y4 = f_u_arrmul12_fa4_5_y4;
  assign f_u_arrmul12_fa5_5_y0 = f_u_arrmul12_fa5_5_f_u_arrmul12_and5_5_y0 ^ f_u_arrmul12_fa5_5_f_u_arrmul12_fa6_4_y2;
  assign f_u_arrmul12_fa5_5_y1 = f_u_arrmul12_fa5_5_f_u_arrmul12_and5_5_y0 & f_u_arrmul12_fa5_5_f_u_arrmul12_fa6_4_y2;
  assign f_u_arrmul12_fa5_5_y2 = f_u_arrmul12_fa5_5_y0 ^ f_u_arrmul12_fa5_5_f_u_arrmul12_fa4_5_y4;
  assign f_u_arrmul12_fa5_5_y3 = f_u_arrmul12_fa5_5_y0 & f_u_arrmul12_fa5_5_f_u_arrmul12_fa4_5_y4;
  assign f_u_arrmul12_fa5_5_y4 = f_u_arrmul12_fa5_5_y1 | f_u_arrmul12_fa5_5_y3;
  assign f_u_arrmul12_and6_5_a_6 = a_6;
  assign f_u_arrmul12_and6_5_b_5 = b_5;
  assign f_u_arrmul12_and6_5_y0 = f_u_arrmul12_and6_5_a_6 & f_u_arrmul12_and6_5_b_5;
  assign f_u_arrmul12_fa6_5_f_u_arrmul12_and6_5_y0 = f_u_arrmul12_and6_5_y0;
  assign f_u_arrmul12_fa6_5_f_u_arrmul12_fa7_4_y2 = f_u_arrmul12_fa7_4_y2;
  assign f_u_arrmul12_fa6_5_f_u_arrmul12_fa5_5_y4 = f_u_arrmul12_fa5_5_y4;
  assign f_u_arrmul12_fa6_5_y0 = f_u_arrmul12_fa6_5_f_u_arrmul12_and6_5_y0 ^ f_u_arrmul12_fa6_5_f_u_arrmul12_fa7_4_y2;
  assign f_u_arrmul12_fa6_5_y1 = f_u_arrmul12_fa6_5_f_u_arrmul12_and6_5_y0 & f_u_arrmul12_fa6_5_f_u_arrmul12_fa7_4_y2;
  assign f_u_arrmul12_fa6_5_y2 = f_u_arrmul12_fa6_5_y0 ^ f_u_arrmul12_fa6_5_f_u_arrmul12_fa5_5_y4;
  assign f_u_arrmul12_fa6_5_y3 = f_u_arrmul12_fa6_5_y0 & f_u_arrmul12_fa6_5_f_u_arrmul12_fa5_5_y4;
  assign f_u_arrmul12_fa6_5_y4 = f_u_arrmul12_fa6_5_y1 | f_u_arrmul12_fa6_5_y3;
  assign f_u_arrmul12_and7_5_a_7 = a_7;
  assign f_u_arrmul12_and7_5_b_5 = b_5;
  assign f_u_arrmul12_and7_5_y0 = f_u_arrmul12_and7_5_a_7 & f_u_arrmul12_and7_5_b_5;
  assign f_u_arrmul12_fa7_5_f_u_arrmul12_and7_5_y0 = f_u_arrmul12_and7_5_y0;
  assign f_u_arrmul12_fa7_5_f_u_arrmul12_fa8_4_y2 = f_u_arrmul12_fa8_4_y2;
  assign f_u_arrmul12_fa7_5_f_u_arrmul12_fa6_5_y4 = f_u_arrmul12_fa6_5_y4;
  assign f_u_arrmul12_fa7_5_y0 = f_u_arrmul12_fa7_5_f_u_arrmul12_and7_5_y0 ^ f_u_arrmul12_fa7_5_f_u_arrmul12_fa8_4_y2;
  assign f_u_arrmul12_fa7_5_y1 = f_u_arrmul12_fa7_5_f_u_arrmul12_and7_5_y0 & f_u_arrmul12_fa7_5_f_u_arrmul12_fa8_4_y2;
  assign f_u_arrmul12_fa7_5_y2 = f_u_arrmul12_fa7_5_y0 ^ f_u_arrmul12_fa7_5_f_u_arrmul12_fa6_5_y4;
  assign f_u_arrmul12_fa7_5_y3 = f_u_arrmul12_fa7_5_y0 & f_u_arrmul12_fa7_5_f_u_arrmul12_fa6_5_y4;
  assign f_u_arrmul12_fa7_5_y4 = f_u_arrmul12_fa7_5_y1 | f_u_arrmul12_fa7_5_y3;
  assign f_u_arrmul12_and8_5_a_8 = a_8;
  assign f_u_arrmul12_and8_5_b_5 = b_5;
  assign f_u_arrmul12_and8_5_y0 = f_u_arrmul12_and8_5_a_8 & f_u_arrmul12_and8_5_b_5;
  assign f_u_arrmul12_fa8_5_f_u_arrmul12_and8_5_y0 = f_u_arrmul12_and8_5_y0;
  assign f_u_arrmul12_fa8_5_f_u_arrmul12_fa9_4_y2 = f_u_arrmul12_fa9_4_y2;
  assign f_u_arrmul12_fa8_5_f_u_arrmul12_fa7_5_y4 = f_u_arrmul12_fa7_5_y4;
  assign f_u_arrmul12_fa8_5_y0 = f_u_arrmul12_fa8_5_f_u_arrmul12_and8_5_y0 ^ f_u_arrmul12_fa8_5_f_u_arrmul12_fa9_4_y2;
  assign f_u_arrmul12_fa8_5_y1 = f_u_arrmul12_fa8_5_f_u_arrmul12_and8_5_y0 & f_u_arrmul12_fa8_5_f_u_arrmul12_fa9_4_y2;
  assign f_u_arrmul12_fa8_5_y2 = f_u_arrmul12_fa8_5_y0 ^ f_u_arrmul12_fa8_5_f_u_arrmul12_fa7_5_y4;
  assign f_u_arrmul12_fa8_5_y3 = f_u_arrmul12_fa8_5_y0 & f_u_arrmul12_fa8_5_f_u_arrmul12_fa7_5_y4;
  assign f_u_arrmul12_fa8_5_y4 = f_u_arrmul12_fa8_5_y1 | f_u_arrmul12_fa8_5_y3;
  assign f_u_arrmul12_and9_5_a_9 = a_9;
  assign f_u_arrmul12_and9_5_b_5 = b_5;
  assign f_u_arrmul12_and9_5_y0 = f_u_arrmul12_and9_5_a_9 & f_u_arrmul12_and9_5_b_5;
  assign f_u_arrmul12_fa9_5_f_u_arrmul12_and9_5_y0 = f_u_arrmul12_and9_5_y0;
  assign f_u_arrmul12_fa9_5_f_u_arrmul12_fa10_4_y2 = f_u_arrmul12_fa10_4_y2;
  assign f_u_arrmul12_fa9_5_f_u_arrmul12_fa8_5_y4 = f_u_arrmul12_fa8_5_y4;
  assign f_u_arrmul12_fa9_5_y0 = f_u_arrmul12_fa9_5_f_u_arrmul12_and9_5_y0 ^ f_u_arrmul12_fa9_5_f_u_arrmul12_fa10_4_y2;
  assign f_u_arrmul12_fa9_5_y1 = f_u_arrmul12_fa9_5_f_u_arrmul12_and9_5_y0 & f_u_arrmul12_fa9_5_f_u_arrmul12_fa10_4_y2;
  assign f_u_arrmul12_fa9_5_y2 = f_u_arrmul12_fa9_5_y0 ^ f_u_arrmul12_fa9_5_f_u_arrmul12_fa8_5_y4;
  assign f_u_arrmul12_fa9_5_y3 = f_u_arrmul12_fa9_5_y0 & f_u_arrmul12_fa9_5_f_u_arrmul12_fa8_5_y4;
  assign f_u_arrmul12_fa9_5_y4 = f_u_arrmul12_fa9_5_y1 | f_u_arrmul12_fa9_5_y3;
  assign f_u_arrmul12_and10_5_a_10 = a_10;
  assign f_u_arrmul12_and10_5_b_5 = b_5;
  assign f_u_arrmul12_and10_5_y0 = f_u_arrmul12_and10_5_a_10 & f_u_arrmul12_and10_5_b_5;
  assign f_u_arrmul12_fa10_5_f_u_arrmul12_and10_5_y0 = f_u_arrmul12_and10_5_y0;
  assign f_u_arrmul12_fa10_5_f_u_arrmul12_fa11_4_y2 = f_u_arrmul12_fa11_4_y2;
  assign f_u_arrmul12_fa10_5_f_u_arrmul12_fa9_5_y4 = f_u_arrmul12_fa9_5_y4;
  assign f_u_arrmul12_fa10_5_y0 = f_u_arrmul12_fa10_5_f_u_arrmul12_and10_5_y0 ^ f_u_arrmul12_fa10_5_f_u_arrmul12_fa11_4_y2;
  assign f_u_arrmul12_fa10_5_y1 = f_u_arrmul12_fa10_5_f_u_arrmul12_and10_5_y0 & f_u_arrmul12_fa10_5_f_u_arrmul12_fa11_4_y2;
  assign f_u_arrmul12_fa10_5_y2 = f_u_arrmul12_fa10_5_y0 ^ f_u_arrmul12_fa10_5_f_u_arrmul12_fa9_5_y4;
  assign f_u_arrmul12_fa10_5_y3 = f_u_arrmul12_fa10_5_y0 & f_u_arrmul12_fa10_5_f_u_arrmul12_fa9_5_y4;
  assign f_u_arrmul12_fa10_5_y4 = f_u_arrmul12_fa10_5_y1 | f_u_arrmul12_fa10_5_y3;
  assign f_u_arrmul12_and11_5_a_11 = a_11;
  assign f_u_arrmul12_and11_5_b_5 = b_5;
  assign f_u_arrmul12_and11_5_y0 = f_u_arrmul12_and11_5_a_11 & f_u_arrmul12_and11_5_b_5;
  assign f_u_arrmul12_fa11_5_f_u_arrmul12_and11_5_y0 = f_u_arrmul12_and11_5_y0;
  assign f_u_arrmul12_fa11_5_f_u_arrmul12_fa11_4_y4 = f_u_arrmul12_fa11_4_y4;
  assign f_u_arrmul12_fa11_5_f_u_arrmul12_fa10_5_y4 = f_u_arrmul12_fa10_5_y4;
  assign f_u_arrmul12_fa11_5_y0 = f_u_arrmul12_fa11_5_f_u_arrmul12_and11_5_y0 ^ f_u_arrmul12_fa11_5_f_u_arrmul12_fa11_4_y4;
  assign f_u_arrmul12_fa11_5_y1 = f_u_arrmul12_fa11_5_f_u_arrmul12_and11_5_y0 & f_u_arrmul12_fa11_5_f_u_arrmul12_fa11_4_y4;
  assign f_u_arrmul12_fa11_5_y2 = f_u_arrmul12_fa11_5_y0 ^ f_u_arrmul12_fa11_5_f_u_arrmul12_fa10_5_y4;
  assign f_u_arrmul12_fa11_5_y3 = f_u_arrmul12_fa11_5_y0 & f_u_arrmul12_fa11_5_f_u_arrmul12_fa10_5_y4;
  assign f_u_arrmul12_fa11_5_y4 = f_u_arrmul12_fa11_5_y1 | f_u_arrmul12_fa11_5_y3;
  assign f_u_arrmul12_and0_6_a_0 = a_0;
  assign f_u_arrmul12_and0_6_b_6 = b_6;
  assign f_u_arrmul12_and0_6_y0 = f_u_arrmul12_and0_6_a_0 & f_u_arrmul12_and0_6_b_6;
  assign f_u_arrmul12_ha0_6_f_u_arrmul12_and0_6_y0 = f_u_arrmul12_and0_6_y0;
  assign f_u_arrmul12_ha0_6_f_u_arrmul12_fa1_5_y2 = f_u_arrmul12_fa1_5_y2;
  assign f_u_arrmul12_ha0_6_y0 = f_u_arrmul12_ha0_6_f_u_arrmul12_and0_6_y0 ^ f_u_arrmul12_ha0_6_f_u_arrmul12_fa1_5_y2;
  assign f_u_arrmul12_ha0_6_y1 = f_u_arrmul12_ha0_6_f_u_arrmul12_and0_6_y0 & f_u_arrmul12_ha0_6_f_u_arrmul12_fa1_5_y2;
  assign f_u_arrmul12_and1_6_a_1 = a_1;
  assign f_u_arrmul12_and1_6_b_6 = b_6;
  assign f_u_arrmul12_and1_6_y0 = f_u_arrmul12_and1_6_a_1 & f_u_arrmul12_and1_6_b_6;
  assign f_u_arrmul12_fa1_6_f_u_arrmul12_and1_6_y0 = f_u_arrmul12_and1_6_y0;
  assign f_u_arrmul12_fa1_6_f_u_arrmul12_fa2_5_y2 = f_u_arrmul12_fa2_5_y2;
  assign f_u_arrmul12_fa1_6_f_u_arrmul12_ha0_6_y1 = f_u_arrmul12_ha0_6_y1;
  assign f_u_arrmul12_fa1_6_y0 = f_u_arrmul12_fa1_6_f_u_arrmul12_and1_6_y0 ^ f_u_arrmul12_fa1_6_f_u_arrmul12_fa2_5_y2;
  assign f_u_arrmul12_fa1_6_y1 = f_u_arrmul12_fa1_6_f_u_arrmul12_and1_6_y0 & f_u_arrmul12_fa1_6_f_u_arrmul12_fa2_5_y2;
  assign f_u_arrmul12_fa1_6_y2 = f_u_arrmul12_fa1_6_y0 ^ f_u_arrmul12_fa1_6_f_u_arrmul12_ha0_6_y1;
  assign f_u_arrmul12_fa1_6_y3 = f_u_arrmul12_fa1_6_y0 & f_u_arrmul12_fa1_6_f_u_arrmul12_ha0_6_y1;
  assign f_u_arrmul12_fa1_6_y4 = f_u_arrmul12_fa1_6_y1 | f_u_arrmul12_fa1_6_y3;
  assign f_u_arrmul12_and2_6_a_2 = a_2;
  assign f_u_arrmul12_and2_6_b_6 = b_6;
  assign f_u_arrmul12_and2_6_y0 = f_u_arrmul12_and2_6_a_2 & f_u_arrmul12_and2_6_b_6;
  assign f_u_arrmul12_fa2_6_f_u_arrmul12_and2_6_y0 = f_u_arrmul12_and2_6_y0;
  assign f_u_arrmul12_fa2_6_f_u_arrmul12_fa3_5_y2 = f_u_arrmul12_fa3_5_y2;
  assign f_u_arrmul12_fa2_6_f_u_arrmul12_fa1_6_y4 = f_u_arrmul12_fa1_6_y4;
  assign f_u_arrmul12_fa2_6_y0 = f_u_arrmul12_fa2_6_f_u_arrmul12_and2_6_y0 ^ f_u_arrmul12_fa2_6_f_u_arrmul12_fa3_5_y2;
  assign f_u_arrmul12_fa2_6_y1 = f_u_arrmul12_fa2_6_f_u_arrmul12_and2_6_y0 & f_u_arrmul12_fa2_6_f_u_arrmul12_fa3_5_y2;
  assign f_u_arrmul12_fa2_6_y2 = f_u_arrmul12_fa2_6_y0 ^ f_u_arrmul12_fa2_6_f_u_arrmul12_fa1_6_y4;
  assign f_u_arrmul12_fa2_6_y3 = f_u_arrmul12_fa2_6_y0 & f_u_arrmul12_fa2_6_f_u_arrmul12_fa1_6_y4;
  assign f_u_arrmul12_fa2_6_y4 = f_u_arrmul12_fa2_6_y1 | f_u_arrmul12_fa2_6_y3;
  assign f_u_arrmul12_and3_6_a_3 = a_3;
  assign f_u_arrmul12_and3_6_b_6 = b_6;
  assign f_u_arrmul12_and3_6_y0 = f_u_arrmul12_and3_6_a_3 & f_u_arrmul12_and3_6_b_6;
  assign f_u_arrmul12_fa3_6_f_u_arrmul12_and3_6_y0 = f_u_arrmul12_and3_6_y0;
  assign f_u_arrmul12_fa3_6_f_u_arrmul12_fa4_5_y2 = f_u_arrmul12_fa4_5_y2;
  assign f_u_arrmul12_fa3_6_f_u_arrmul12_fa2_6_y4 = f_u_arrmul12_fa2_6_y4;
  assign f_u_arrmul12_fa3_6_y0 = f_u_arrmul12_fa3_6_f_u_arrmul12_and3_6_y0 ^ f_u_arrmul12_fa3_6_f_u_arrmul12_fa4_5_y2;
  assign f_u_arrmul12_fa3_6_y1 = f_u_arrmul12_fa3_6_f_u_arrmul12_and3_6_y0 & f_u_arrmul12_fa3_6_f_u_arrmul12_fa4_5_y2;
  assign f_u_arrmul12_fa3_6_y2 = f_u_arrmul12_fa3_6_y0 ^ f_u_arrmul12_fa3_6_f_u_arrmul12_fa2_6_y4;
  assign f_u_arrmul12_fa3_6_y3 = f_u_arrmul12_fa3_6_y0 & f_u_arrmul12_fa3_6_f_u_arrmul12_fa2_6_y4;
  assign f_u_arrmul12_fa3_6_y4 = f_u_arrmul12_fa3_6_y1 | f_u_arrmul12_fa3_6_y3;
  assign f_u_arrmul12_and4_6_a_4 = a_4;
  assign f_u_arrmul12_and4_6_b_6 = b_6;
  assign f_u_arrmul12_and4_6_y0 = f_u_arrmul12_and4_6_a_4 & f_u_arrmul12_and4_6_b_6;
  assign f_u_arrmul12_fa4_6_f_u_arrmul12_and4_6_y0 = f_u_arrmul12_and4_6_y0;
  assign f_u_arrmul12_fa4_6_f_u_arrmul12_fa5_5_y2 = f_u_arrmul12_fa5_5_y2;
  assign f_u_arrmul12_fa4_6_f_u_arrmul12_fa3_6_y4 = f_u_arrmul12_fa3_6_y4;
  assign f_u_arrmul12_fa4_6_y0 = f_u_arrmul12_fa4_6_f_u_arrmul12_and4_6_y0 ^ f_u_arrmul12_fa4_6_f_u_arrmul12_fa5_5_y2;
  assign f_u_arrmul12_fa4_6_y1 = f_u_arrmul12_fa4_6_f_u_arrmul12_and4_6_y0 & f_u_arrmul12_fa4_6_f_u_arrmul12_fa5_5_y2;
  assign f_u_arrmul12_fa4_6_y2 = f_u_arrmul12_fa4_6_y0 ^ f_u_arrmul12_fa4_6_f_u_arrmul12_fa3_6_y4;
  assign f_u_arrmul12_fa4_6_y3 = f_u_arrmul12_fa4_6_y0 & f_u_arrmul12_fa4_6_f_u_arrmul12_fa3_6_y4;
  assign f_u_arrmul12_fa4_6_y4 = f_u_arrmul12_fa4_6_y1 | f_u_arrmul12_fa4_6_y3;
  assign f_u_arrmul12_and5_6_a_5 = a_5;
  assign f_u_arrmul12_and5_6_b_6 = b_6;
  assign f_u_arrmul12_and5_6_y0 = f_u_arrmul12_and5_6_a_5 & f_u_arrmul12_and5_6_b_6;
  assign f_u_arrmul12_fa5_6_f_u_arrmul12_and5_6_y0 = f_u_arrmul12_and5_6_y0;
  assign f_u_arrmul12_fa5_6_f_u_arrmul12_fa6_5_y2 = f_u_arrmul12_fa6_5_y2;
  assign f_u_arrmul12_fa5_6_f_u_arrmul12_fa4_6_y4 = f_u_arrmul12_fa4_6_y4;
  assign f_u_arrmul12_fa5_6_y0 = f_u_arrmul12_fa5_6_f_u_arrmul12_and5_6_y0 ^ f_u_arrmul12_fa5_6_f_u_arrmul12_fa6_5_y2;
  assign f_u_arrmul12_fa5_6_y1 = f_u_arrmul12_fa5_6_f_u_arrmul12_and5_6_y0 & f_u_arrmul12_fa5_6_f_u_arrmul12_fa6_5_y2;
  assign f_u_arrmul12_fa5_6_y2 = f_u_arrmul12_fa5_6_y0 ^ f_u_arrmul12_fa5_6_f_u_arrmul12_fa4_6_y4;
  assign f_u_arrmul12_fa5_6_y3 = f_u_arrmul12_fa5_6_y0 & f_u_arrmul12_fa5_6_f_u_arrmul12_fa4_6_y4;
  assign f_u_arrmul12_fa5_6_y4 = f_u_arrmul12_fa5_6_y1 | f_u_arrmul12_fa5_6_y3;
  assign f_u_arrmul12_and6_6_a_6 = a_6;
  assign f_u_arrmul12_and6_6_b_6 = b_6;
  assign f_u_arrmul12_and6_6_y0 = f_u_arrmul12_and6_6_a_6 & f_u_arrmul12_and6_6_b_6;
  assign f_u_arrmul12_fa6_6_f_u_arrmul12_and6_6_y0 = f_u_arrmul12_and6_6_y0;
  assign f_u_arrmul12_fa6_6_f_u_arrmul12_fa7_5_y2 = f_u_arrmul12_fa7_5_y2;
  assign f_u_arrmul12_fa6_6_f_u_arrmul12_fa5_6_y4 = f_u_arrmul12_fa5_6_y4;
  assign f_u_arrmul12_fa6_6_y0 = f_u_arrmul12_fa6_6_f_u_arrmul12_and6_6_y0 ^ f_u_arrmul12_fa6_6_f_u_arrmul12_fa7_5_y2;
  assign f_u_arrmul12_fa6_6_y1 = f_u_arrmul12_fa6_6_f_u_arrmul12_and6_6_y0 & f_u_arrmul12_fa6_6_f_u_arrmul12_fa7_5_y2;
  assign f_u_arrmul12_fa6_6_y2 = f_u_arrmul12_fa6_6_y0 ^ f_u_arrmul12_fa6_6_f_u_arrmul12_fa5_6_y4;
  assign f_u_arrmul12_fa6_6_y3 = f_u_arrmul12_fa6_6_y0 & f_u_arrmul12_fa6_6_f_u_arrmul12_fa5_6_y4;
  assign f_u_arrmul12_fa6_6_y4 = f_u_arrmul12_fa6_6_y1 | f_u_arrmul12_fa6_6_y3;
  assign f_u_arrmul12_and7_6_a_7 = a_7;
  assign f_u_arrmul12_and7_6_b_6 = b_6;
  assign f_u_arrmul12_and7_6_y0 = f_u_arrmul12_and7_6_a_7 & f_u_arrmul12_and7_6_b_6;
  assign f_u_arrmul12_fa7_6_f_u_arrmul12_and7_6_y0 = f_u_arrmul12_and7_6_y0;
  assign f_u_arrmul12_fa7_6_f_u_arrmul12_fa8_5_y2 = f_u_arrmul12_fa8_5_y2;
  assign f_u_arrmul12_fa7_6_f_u_arrmul12_fa6_6_y4 = f_u_arrmul12_fa6_6_y4;
  assign f_u_arrmul12_fa7_6_y0 = f_u_arrmul12_fa7_6_f_u_arrmul12_and7_6_y0 ^ f_u_arrmul12_fa7_6_f_u_arrmul12_fa8_5_y2;
  assign f_u_arrmul12_fa7_6_y1 = f_u_arrmul12_fa7_6_f_u_arrmul12_and7_6_y0 & f_u_arrmul12_fa7_6_f_u_arrmul12_fa8_5_y2;
  assign f_u_arrmul12_fa7_6_y2 = f_u_arrmul12_fa7_6_y0 ^ f_u_arrmul12_fa7_6_f_u_arrmul12_fa6_6_y4;
  assign f_u_arrmul12_fa7_6_y3 = f_u_arrmul12_fa7_6_y0 & f_u_arrmul12_fa7_6_f_u_arrmul12_fa6_6_y4;
  assign f_u_arrmul12_fa7_6_y4 = f_u_arrmul12_fa7_6_y1 | f_u_arrmul12_fa7_6_y3;
  assign f_u_arrmul12_and8_6_a_8 = a_8;
  assign f_u_arrmul12_and8_6_b_6 = b_6;
  assign f_u_arrmul12_and8_6_y0 = f_u_arrmul12_and8_6_a_8 & f_u_arrmul12_and8_6_b_6;
  assign f_u_arrmul12_fa8_6_f_u_arrmul12_and8_6_y0 = f_u_arrmul12_and8_6_y0;
  assign f_u_arrmul12_fa8_6_f_u_arrmul12_fa9_5_y2 = f_u_arrmul12_fa9_5_y2;
  assign f_u_arrmul12_fa8_6_f_u_arrmul12_fa7_6_y4 = f_u_arrmul12_fa7_6_y4;
  assign f_u_arrmul12_fa8_6_y0 = f_u_arrmul12_fa8_6_f_u_arrmul12_and8_6_y0 ^ f_u_arrmul12_fa8_6_f_u_arrmul12_fa9_5_y2;
  assign f_u_arrmul12_fa8_6_y1 = f_u_arrmul12_fa8_6_f_u_arrmul12_and8_6_y0 & f_u_arrmul12_fa8_6_f_u_arrmul12_fa9_5_y2;
  assign f_u_arrmul12_fa8_6_y2 = f_u_arrmul12_fa8_6_y0 ^ f_u_arrmul12_fa8_6_f_u_arrmul12_fa7_6_y4;
  assign f_u_arrmul12_fa8_6_y3 = f_u_arrmul12_fa8_6_y0 & f_u_arrmul12_fa8_6_f_u_arrmul12_fa7_6_y4;
  assign f_u_arrmul12_fa8_6_y4 = f_u_arrmul12_fa8_6_y1 | f_u_arrmul12_fa8_6_y3;
  assign f_u_arrmul12_and9_6_a_9 = a_9;
  assign f_u_arrmul12_and9_6_b_6 = b_6;
  assign f_u_arrmul12_and9_6_y0 = f_u_arrmul12_and9_6_a_9 & f_u_arrmul12_and9_6_b_6;
  assign f_u_arrmul12_fa9_6_f_u_arrmul12_and9_6_y0 = f_u_arrmul12_and9_6_y0;
  assign f_u_arrmul12_fa9_6_f_u_arrmul12_fa10_5_y2 = f_u_arrmul12_fa10_5_y2;
  assign f_u_arrmul12_fa9_6_f_u_arrmul12_fa8_6_y4 = f_u_arrmul12_fa8_6_y4;
  assign f_u_arrmul12_fa9_6_y0 = f_u_arrmul12_fa9_6_f_u_arrmul12_and9_6_y0 ^ f_u_arrmul12_fa9_6_f_u_arrmul12_fa10_5_y2;
  assign f_u_arrmul12_fa9_6_y1 = f_u_arrmul12_fa9_6_f_u_arrmul12_and9_6_y0 & f_u_arrmul12_fa9_6_f_u_arrmul12_fa10_5_y2;
  assign f_u_arrmul12_fa9_6_y2 = f_u_arrmul12_fa9_6_y0 ^ f_u_arrmul12_fa9_6_f_u_arrmul12_fa8_6_y4;
  assign f_u_arrmul12_fa9_6_y3 = f_u_arrmul12_fa9_6_y0 & f_u_arrmul12_fa9_6_f_u_arrmul12_fa8_6_y4;
  assign f_u_arrmul12_fa9_6_y4 = f_u_arrmul12_fa9_6_y1 | f_u_arrmul12_fa9_6_y3;
  assign f_u_arrmul12_and10_6_a_10 = a_10;
  assign f_u_arrmul12_and10_6_b_6 = b_6;
  assign f_u_arrmul12_and10_6_y0 = f_u_arrmul12_and10_6_a_10 & f_u_arrmul12_and10_6_b_6;
  assign f_u_arrmul12_fa10_6_f_u_arrmul12_and10_6_y0 = f_u_arrmul12_and10_6_y0;
  assign f_u_arrmul12_fa10_6_f_u_arrmul12_fa11_5_y2 = f_u_arrmul12_fa11_5_y2;
  assign f_u_arrmul12_fa10_6_f_u_arrmul12_fa9_6_y4 = f_u_arrmul12_fa9_6_y4;
  assign f_u_arrmul12_fa10_6_y0 = f_u_arrmul12_fa10_6_f_u_arrmul12_and10_6_y0 ^ f_u_arrmul12_fa10_6_f_u_arrmul12_fa11_5_y2;
  assign f_u_arrmul12_fa10_6_y1 = f_u_arrmul12_fa10_6_f_u_arrmul12_and10_6_y0 & f_u_arrmul12_fa10_6_f_u_arrmul12_fa11_5_y2;
  assign f_u_arrmul12_fa10_6_y2 = f_u_arrmul12_fa10_6_y0 ^ f_u_arrmul12_fa10_6_f_u_arrmul12_fa9_6_y4;
  assign f_u_arrmul12_fa10_6_y3 = f_u_arrmul12_fa10_6_y0 & f_u_arrmul12_fa10_6_f_u_arrmul12_fa9_6_y4;
  assign f_u_arrmul12_fa10_6_y4 = f_u_arrmul12_fa10_6_y1 | f_u_arrmul12_fa10_6_y3;
  assign f_u_arrmul12_and11_6_a_11 = a_11;
  assign f_u_arrmul12_and11_6_b_6 = b_6;
  assign f_u_arrmul12_and11_6_y0 = f_u_arrmul12_and11_6_a_11 & f_u_arrmul12_and11_6_b_6;
  assign f_u_arrmul12_fa11_6_f_u_arrmul12_and11_6_y0 = f_u_arrmul12_and11_6_y0;
  assign f_u_arrmul12_fa11_6_f_u_arrmul12_fa11_5_y4 = f_u_arrmul12_fa11_5_y4;
  assign f_u_arrmul12_fa11_6_f_u_arrmul12_fa10_6_y4 = f_u_arrmul12_fa10_6_y4;
  assign f_u_arrmul12_fa11_6_y0 = f_u_arrmul12_fa11_6_f_u_arrmul12_and11_6_y0 ^ f_u_arrmul12_fa11_6_f_u_arrmul12_fa11_5_y4;
  assign f_u_arrmul12_fa11_6_y1 = f_u_arrmul12_fa11_6_f_u_arrmul12_and11_6_y0 & f_u_arrmul12_fa11_6_f_u_arrmul12_fa11_5_y4;
  assign f_u_arrmul12_fa11_6_y2 = f_u_arrmul12_fa11_6_y0 ^ f_u_arrmul12_fa11_6_f_u_arrmul12_fa10_6_y4;
  assign f_u_arrmul12_fa11_6_y3 = f_u_arrmul12_fa11_6_y0 & f_u_arrmul12_fa11_6_f_u_arrmul12_fa10_6_y4;
  assign f_u_arrmul12_fa11_6_y4 = f_u_arrmul12_fa11_6_y1 | f_u_arrmul12_fa11_6_y3;
  assign f_u_arrmul12_and0_7_a_0 = a_0;
  assign f_u_arrmul12_and0_7_b_7 = b_7;
  assign f_u_arrmul12_and0_7_y0 = f_u_arrmul12_and0_7_a_0 & f_u_arrmul12_and0_7_b_7;
  assign f_u_arrmul12_ha0_7_f_u_arrmul12_and0_7_y0 = f_u_arrmul12_and0_7_y0;
  assign f_u_arrmul12_ha0_7_f_u_arrmul12_fa1_6_y2 = f_u_arrmul12_fa1_6_y2;
  assign f_u_arrmul12_ha0_7_y0 = f_u_arrmul12_ha0_7_f_u_arrmul12_and0_7_y0 ^ f_u_arrmul12_ha0_7_f_u_arrmul12_fa1_6_y2;
  assign f_u_arrmul12_ha0_7_y1 = f_u_arrmul12_ha0_7_f_u_arrmul12_and0_7_y0 & f_u_arrmul12_ha0_7_f_u_arrmul12_fa1_6_y2;
  assign f_u_arrmul12_and1_7_a_1 = a_1;
  assign f_u_arrmul12_and1_7_b_7 = b_7;
  assign f_u_arrmul12_and1_7_y0 = f_u_arrmul12_and1_7_a_1 & f_u_arrmul12_and1_7_b_7;
  assign f_u_arrmul12_fa1_7_f_u_arrmul12_and1_7_y0 = f_u_arrmul12_and1_7_y0;
  assign f_u_arrmul12_fa1_7_f_u_arrmul12_fa2_6_y2 = f_u_arrmul12_fa2_6_y2;
  assign f_u_arrmul12_fa1_7_f_u_arrmul12_ha0_7_y1 = f_u_arrmul12_ha0_7_y1;
  assign f_u_arrmul12_fa1_7_y0 = f_u_arrmul12_fa1_7_f_u_arrmul12_and1_7_y0 ^ f_u_arrmul12_fa1_7_f_u_arrmul12_fa2_6_y2;
  assign f_u_arrmul12_fa1_7_y1 = f_u_arrmul12_fa1_7_f_u_arrmul12_and1_7_y0 & f_u_arrmul12_fa1_7_f_u_arrmul12_fa2_6_y2;
  assign f_u_arrmul12_fa1_7_y2 = f_u_arrmul12_fa1_7_y0 ^ f_u_arrmul12_fa1_7_f_u_arrmul12_ha0_7_y1;
  assign f_u_arrmul12_fa1_7_y3 = f_u_arrmul12_fa1_7_y0 & f_u_arrmul12_fa1_7_f_u_arrmul12_ha0_7_y1;
  assign f_u_arrmul12_fa1_7_y4 = f_u_arrmul12_fa1_7_y1 | f_u_arrmul12_fa1_7_y3;
  assign f_u_arrmul12_and2_7_a_2 = a_2;
  assign f_u_arrmul12_and2_7_b_7 = b_7;
  assign f_u_arrmul12_and2_7_y0 = f_u_arrmul12_and2_7_a_2 & f_u_arrmul12_and2_7_b_7;
  assign f_u_arrmul12_fa2_7_f_u_arrmul12_and2_7_y0 = f_u_arrmul12_and2_7_y0;
  assign f_u_arrmul12_fa2_7_f_u_arrmul12_fa3_6_y2 = f_u_arrmul12_fa3_6_y2;
  assign f_u_arrmul12_fa2_7_f_u_arrmul12_fa1_7_y4 = f_u_arrmul12_fa1_7_y4;
  assign f_u_arrmul12_fa2_7_y0 = f_u_arrmul12_fa2_7_f_u_arrmul12_and2_7_y0 ^ f_u_arrmul12_fa2_7_f_u_arrmul12_fa3_6_y2;
  assign f_u_arrmul12_fa2_7_y1 = f_u_arrmul12_fa2_7_f_u_arrmul12_and2_7_y0 & f_u_arrmul12_fa2_7_f_u_arrmul12_fa3_6_y2;
  assign f_u_arrmul12_fa2_7_y2 = f_u_arrmul12_fa2_7_y0 ^ f_u_arrmul12_fa2_7_f_u_arrmul12_fa1_7_y4;
  assign f_u_arrmul12_fa2_7_y3 = f_u_arrmul12_fa2_7_y0 & f_u_arrmul12_fa2_7_f_u_arrmul12_fa1_7_y4;
  assign f_u_arrmul12_fa2_7_y4 = f_u_arrmul12_fa2_7_y1 | f_u_arrmul12_fa2_7_y3;
  assign f_u_arrmul12_and3_7_a_3 = a_3;
  assign f_u_arrmul12_and3_7_b_7 = b_7;
  assign f_u_arrmul12_and3_7_y0 = f_u_arrmul12_and3_7_a_3 & f_u_arrmul12_and3_7_b_7;
  assign f_u_arrmul12_fa3_7_f_u_arrmul12_and3_7_y0 = f_u_arrmul12_and3_7_y0;
  assign f_u_arrmul12_fa3_7_f_u_arrmul12_fa4_6_y2 = f_u_arrmul12_fa4_6_y2;
  assign f_u_arrmul12_fa3_7_f_u_arrmul12_fa2_7_y4 = f_u_arrmul12_fa2_7_y4;
  assign f_u_arrmul12_fa3_7_y0 = f_u_arrmul12_fa3_7_f_u_arrmul12_and3_7_y0 ^ f_u_arrmul12_fa3_7_f_u_arrmul12_fa4_6_y2;
  assign f_u_arrmul12_fa3_7_y1 = f_u_arrmul12_fa3_7_f_u_arrmul12_and3_7_y0 & f_u_arrmul12_fa3_7_f_u_arrmul12_fa4_6_y2;
  assign f_u_arrmul12_fa3_7_y2 = f_u_arrmul12_fa3_7_y0 ^ f_u_arrmul12_fa3_7_f_u_arrmul12_fa2_7_y4;
  assign f_u_arrmul12_fa3_7_y3 = f_u_arrmul12_fa3_7_y0 & f_u_arrmul12_fa3_7_f_u_arrmul12_fa2_7_y4;
  assign f_u_arrmul12_fa3_7_y4 = f_u_arrmul12_fa3_7_y1 | f_u_arrmul12_fa3_7_y3;
  assign f_u_arrmul12_and4_7_a_4 = a_4;
  assign f_u_arrmul12_and4_7_b_7 = b_7;
  assign f_u_arrmul12_and4_7_y0 = f_u_arrmul12_and4_7_a_4 & f_u_arrmul12_and4_7_b_7;
  assign f_u_arrmul12_fa4_7_f_u_arrmul12_and4_7_y0 = f_u_arrmul12_and4_7_y0;
  assign f_u_arrmul12_fa4_7_f_u_arrmul12_fa5_6_y2 = f_u_arrmul12_fa5_6_y2;
  assign f_u_arrmul12_fa4_7_f_u_arrmul12_fa3_7_y4 = f_u_arrmul12_fa3_7_y4;
  assign f_u_arrmul12_fa4_7_y0 = f_u_arrmul12_fa4_7_f_u_arrmul12_and4_7_y0 ^ f_u_arrmul12_fa4_7_f_u_arrmul12_fa5_6_y2;
  assign f_u_arrmul12_fa4_7_y1 = f_u_arrmul12_fa4_7_f_u_arrmul12_and4_7_y0 & f_u_arrmul12_fa4_7_f_u_arrmul12_fa5_6_y2;
  assign f_u_arrmul12_fa4_7_y2 = f_u_arrmul12_fa4_7_y0 ^ f_u_arrmul12_fa4_7_f_u_arrmul12_fa3_7_y4;
  assign f_u_arrmul12_fa4_7_y3 = f_u_arrmul12_fa4_7_y0 & f_u_arrmul12_fa4_7_f_u_arrmul12_fa3_7_y4;
  assign f_u_arrmul12_fa4_7_y4 = f_u_arrmul12_fa4_7_y1 | f_u_arrmul12_fa4_7_y3;
  assign f_u_arrmul12_and5_7_a_5 = a_5;
  assign f_u_arrmul12_and5_7_b_7 = b_7;
  assign f_u_arrmul12_and5_7_y0 = f_u_arrmul12_and5_7_a_5 & f_u_arrmul12_and5_7_b_7;
  assign f_u_arrmul12_fa5_7_f_u_arrmul12_and5_7_y0 = f_u_arrmul12_and5_7_y0;
  assign f_u_arrmul12_fa5_7_f_u_arrmul12_fa6_6_y2 = f_u_arrmul12_fa6_6_y2;
  assign f_u_arrmul12_fa5_7_f_u_arrmul12_fa4_7_y4 = f_u_arrmul12_fa4_7_y4;
  assign f_u_arrmul12_fa5_7_y0 = f_u_arrmul12_fa5_7_f_u_arrmul12_and5_7_y0 ^ f_u_arrmul12_fa5_7_f_u_arrmul12_fa6_6_y2;
  assign f_u_arrmul12_fa5_7_y1 = f_u_arrmul12_fa5_7_f_u_arrmul12_and5_7_y0 & f_u_arrmul12_fa5_7_f_u_arrmul12_fa6_6_y2;
  assign f_u_arrmul12_fa5_7_y2 = f_u_arrmul12_fa5_7_y0 ^ f_u_arrmul12_fa5_7_f_u_arrmul12_fa4_7_y4;
  assign f_u_arrmul12_fa5_7_y3 = f_u_arrmul12_fa5_7_y0 & f_u_arrmul12_fa5_7_f_u_arrmul12_fa4_7_y4;
  assign f_u_arrmul12_fa5_7_y4 = f_u_arrmul12_fa5_7_y1 | f_u_arrmul12_fa5_7_y3;
  assign f_u_arrmul12_and6_7_a_6 = a_6;
  assign f_u_arrmul12_and6_7_b_7 = b_7;
  assign f_u_arrmul12_and6_7_y0 = f_u_arrmul12_and6_7_a_6 & f_u_arrmul12_and6_7_b_7;
  assign f_u_arrmul12_fa6_7_f_u_arrmul12_and6_7_y0 = f_u_arrmul12_and6_7_y0;
  assign f_u_arrmul12_fa6_7_f_u_arrmul12_fa7_6_y2 = f_u_arrmul12_fa7_6_y2;
  assign f_u_arrmul12_fa6_7_f_u_arrmul12_fa5_7_y4 = f_u_arrmul12_fa5_7_y4;
  assign f_u_arrmul12_fa6_7_y0 = f_u_arrmul12_fa6_7_f_u_arrmul12_and6_7_y0 ^ f_u_arrmul12_fa6_7_f_u_arrmul12_fa7_6_y2;
  assign f_u_arrmul12_fa6_7_y1 = f_u_arrmul12_fa6_7_f_u_arrmul12_and6_7_y0 & f_u_arrmul12_fa6_7_f_u_arrmul12_fa7_6_y2;
  assign f_u_arrmul12_fa6_7_y2 = f_u_arrmul12_fa6_7_y0 ^ f_u_arrmul12_fa6_7_f_u_arrmul12_fa5_7_y4;
  assign f_u_arrmul12_fa6_7_y3 = f_u_arrmul12_fa6_7_y0 & f_u_arrmul12_fa6_7_f_u_arrmul12_fa5_7_y4;
  assign f_u_arrmul12_fa6_7_y4 = f_u_arrmul12_fa6_7_y1 | f_u_arrmul12_fa6_7_y3;
  assign f_u_arrmul12_and7_7_a_7 = a_7;
  assign f_u_arrmul12_and7_7_b_7 = b_7;
  assign f_u_arrmul12_and7_7_y0 = f_u_arrmul12_and7_7_a_7 & f_u_arrmul12_and7_7_b_7;
  assign f_u_arrmul12_fa7_7_f_u_arrmul12_and7_7_y0 = f_u_arrmul12_and7_7_y0;
  assign f_u_arrmul12_fa7_7_f_u_arrmul12_fa8_6_y2 = f_u_arrmul12_fa8_6_y2;
  assign f_u_arrmul12_fa7_7_f_u_arrmul12_fa6_7_y4 = f_u_arrmul12_fa6_7_y4;
  assign f_u_arrmul12_fa7_7_y0 = f_u_arrmul12_fa7_7_f_u_arrmul12_and7_7_y0 ^ f_u_arrmul12_fa7_7_f_u_arrmul12_fa8_6_y2;
  assign f_u_arrmul12_fa7_7_y1 = f_u_arrmul12_fa7_7_f_u_arrmul12_and7_7_y0 & f_u_arrmul12_fa7_7_f_u_arrmul12_fa8_6_y2;
  assign f_u_arrmul12_fa7_7_y2 = f_u_arrmul12_fa7_7_y0 ^ f_u_arrmul12_fa7_7_f_u_arrmul12_fa6_7_y4;
  assign f_u_arrmul12_fa7_7_y3 = f_u_arrmul12_fa7_7_y0 & f_u_arrmul12_fa7_7_f_u_arrmul12_fa6_7_y4;
  assign f_u_arrmul12_fa7_7_y4 = f_u_arrmul12_fa7_7_y1 | f_u_arrmul12_fa7_7_y3;
  assign f_u_arrmul12_and8_7_a_8 = a_8;
  assign f_u_arrmul12_and8_7_b_7 = b_7;
  assign f_u_arrmul12_and8_7_y0 = f_u_arrmul12_and8_7_a_8 & f_u_arrmul12_and8_7_b_7;
  assign f_u_arrmul12_fa8_7_f_u_arrmul12_and8_7_y0 = f_u_arrmul12_and8_7_y0;
  assign f_u_arrmul12_fa8_7_f_u_arrmul12_fa9_6_y2 = f_u_arrmul12_fa9_6_y2;
  assign f_u_arrmul12_fa8_7_f_u_arrmul12_fa7_7_y4 = f_u_arrmul12_fa7_7_y4;
  assign f_u_arrmul12_fa8_7_y0 = f_u_arrmul12_fa8_7_f_u_arrmul12_and8_7_y0 ^ f_u_arrmul12_fa8_7_f_u_arrmul12_fa9_6_y2;
  assign f_u_arrmul12_fa8_7_y1 = f_u_arrmul12_fa8_7_f_u_arrmul12_and8_7_y0 & f_u_arrmul12_fa8_7_f_u_arrmul12_fa9_6_y2;
  assign f_u_arrmul12_fa8_7_y2 = f_u_arrmul12_fa8_7_y0 ^ f_u_arrmul12_fa8_7_f_u_arrmul12_fa7_7_y4;
  assign f_u_arrmul12_fa8_7_y3 = f_u_arrmul12_fa8_7_y0 & f_u_arrmul12_fa8_7_f_u_arrmul12_fa7_7_y4;
  assign f_u_arrmul12_fa8_7_y4 = f_u_arrmul12_fa8_7_y1 | f_u_arrmul12_fa8_7_y3;
  assign f_u_arrmul12_and9_7_a_9 = a_9;
  assign f_u_arrmul12_and9_7_b_7 = b_7;
  assign f_u_arrmul12_and9_7_y0 = f_u_arrmul12_and9_7_a_9 & f_u_arrmul12_and9_7_b_7;
  assign f_u_arrmul12_fa9_7_f_u_arrmul12_and9_7_y0 = f_u_arrmul12_and9_7_y0;
  assign f_u_arrmul12_fa9_7_f_u_arrmul12_fa10_6_y2 = f_u_arrmul12_fa10_6_y2;
  assign f_u_arrmul12_fa9_7_f_u_arrmul12_fa8_7_y4 = f_u_arrmul12_fa8_7_y4;
  assign f_u_arrmul12_fa9_7_y0 = f_u_arrmul12_fa9_7_f_u_arrmul12_and9_7_y0 ^ f_u_arrmul12_fa9_7_f_u_arrmul12_fa10_6_y2;
  assign f_u_arrmul12_fa9_7_y1 = f_u_arrmul12_fa9_7_f_u_arrmul12_and9_7_y0 & f_u_arrmul12_fa9_7_f_u_arrmul12_fa10_6_y2;
  assign f_u_arrmul12_fa9_7_y2 = f_u_arrmul12_fa9_7_y0 ^ f_u_arrmul12_fa9_7_f_u_arrmul12_fa8_7_y4;
  assign f_u_arrmul12_fa9_7_y3 = f_u_arrmul12_fa9_7_y0 & f_u_arrmul12_fa9_7_f_u_arrmul12_fa8_7_y4;
  assign f_u_arrmul12_fa9_7_y4 = f_u_arrmul12_fa9_7_y1 | f_u_arrmul12_fa9_7_y3;
  assign f_u_arrmul12_and10_7_a_10 = a_10;
  assign f_u_arrmul12_and10_7_b_7 = b_7;
  assign f_u_arrmul12_and10_7_y0 = f_u_arrmul12_and10_7_a_10 & f_u_arrmul12_and10_7_b_7;
  assign f_u_arrmul12_fa10_7_f_u_arrmul12_and10_7_y0 = f_u_arrmul12_and10_7_y0;
  assign f_u_arrmul12_fa10_7_f_u_arrmul12_fa11_6_y2 = f_u_arrmul12_fa11_6_y2;
  assign f_u_arrmul12_fa10_7_f_u_arrmul12_fa9_7_y4 = f_u_arrmul12_fa9_7_y4;
  assign f_u_arrmul12_fa10_7_y0 = f_u_arrmul12_fa10_7_f_u_arrmul12_and10_7_y0 ^ f_u_arrmul12_fa10_7_f_u_arrmul12_fa11_6_y2;
  assign f_u_arrmul12_fa10_7_y1 = f_u_arrmul12_fa10_7_f_u_arrmul12_and10_7_y0 & f_u_arrmul12_fa10_7_f_u_arrmul12_fa11_6_y2;
  assign f_u_arrmul12_fa10_7_y2 = f_u_arrmul12_fa10_7_y0 ^ f_u_arrmul12_fa10_7_f_u_arrmul12_fa9_7_y4;
  assign f_u_arrmul12_fa10_7_y3 = f_u_arrmul12_fa10_7_y0 & f_u_arrmul12_fa10_7_f_u_arrmul12_fa9_7_y4;
  assign f_u_arrmul12_fa10_7_y4 = f_u_arrmul12_fa10_7_y1 | f_u_arrmul12_fa10_7_y3;
  assign f_u_arrmul12_and11_7_a_11 = a_11;
  assign f_u_arrmul12_and11_7_b_7 = b_7;
  assign f_u_arrmul12_and11_7_y0 = f_u_arrmul12_and11_7_a_11 & f_u_arrmul12_and11_7_b_7;
  assign f_u_arrmul12_fa11_7_f_u_arrmul12_and11_7_y0 = f_u_arrmul12_and11_7_y0;
  assign f_u_arrmul12_fa11_7_f_u_arrmul12_fa11_6_y4 = f_u_arrmul12_fa11_6_y4;
  assign f_u_arrmul12_fa11_7_f_u_arrmul12_fa10_7_y4 = f_u_arrmul12_fa10_7_y4;
  assign f_u_arrmul12_fa11_7_y0 = f_u_arrmul12_fa11_7_f_u_arrmul12_and11_7_y0 ^ f_u_arrmul12_fa11_7_f_u_arrmul12_fa11_6_y4;
  assign f_u_arrmul12_fa11_7_y1 = f_u_arrmul12_fa11_7_f_u_arrmul12_and11_7_y0 & f_u_arrmul12_fa11_7_f_u_arrmul12_fa11_6_y4;
  assign f_u_arrmul12_fa11_7_y2 = f_u_arrmul12_fa11_7_y0 ^ f_u_arrmul12_fa11_7_f_u_arrmul12_fa10_7_y4;
  assign f_u_arrmul12_fa11_7_y3 = f_u_arrmul12_fa11_7_y0 & f_u_arrmul12_fa11_7_f_u_arrmul12_fa10_7_y4;
  assign f_u_arrmul12_fa11_7_y4 = f_u_arrmul12_fa11_7_y1 | f_u_arrmul12_fa11_7_y3;
  assign f_u_arrmul12_and0_8_a_0 = a_0;
  assign f_u_arrmul12_and0_8_b_8 = b_8;
  assign f_u_arrmul12_and0_8_y0 = f_u_arrmul12_and0_8_a_0 & f_u_arrmul12_and0_8_b_8;
  assign f_u_arrmul12_ha0_8_f_u_arrmul12_and0_8_y0 = f_u_arrmul12_and0_8_y0;
  assign f_u_arrmul12_ha0_8_f_u_arrmul12_fa1_7_y2 = f_u_arrmul12_fa1_7_y2;
  assign f_u_arrmul12_ha0_8_y0 = f_u_arrmul12_ha0_8_f_u_arrmul12_and0_8_y0 ^ f_u_arrmul12_ha0_8_f_u_arrmul12_fa1_7_y2;
  assign f_u_arrmul12_ha0_8_y1 = f_u_arrmul12_ha0_8_f_u_arrmul12_and0_8_y0 & f_u_arrmul12_ha0_8_f_u_arrmul12_fa1_7_y2;
  assign f_u_arrmul12_and1_8_a_1 = a_1;
  assign f_u_arrmul12_and1_8_b_8 = b_8;
  assign f_u_arrmul12_and1_8_y0 = f_u_arrmul12_and1_8_a_1 & f_u_arrmul12_and1_8_b_8;
  assign f_u_arrmul12_fa1_8_f_u_arrmul12_and1_8_y0 = f_u_arrmul12_and1_8_y0;
  assign f_u_arrmul12_fa1_8_f_u_arrmul12_fa2_7_y2 = f_u_arrmul12_fa2_7_y2;
  assign f_u_arrmul12_fa1_8_f_u_arrmul12_ha0_8_y1 = f_u_arrmul12_ha0_8_y1;
  assign f_u_arrmul12_fa1_8_y0 = f_u_arrmul12_fa1_8_f_u_arrmul12_and1_8_y0 ^ f_u_arrmul12_fa1_8_f_u_arrmul12_fa2_7_y2;
  assign f_u_arrmul12_fa1_8_y1 = f_u_arrmul12_fa1_8_f_u_arrmul12_and1_8_y0 & f_u_arrmul12_fa1_8_f_u_arrmul12_fa2_7_y2;
  assign f_u_arrmul12_fa1_8_y2 = f_u_arrmul12_fa1_8_y0 ^ f_u_arrmul12_fa1_8_f_u_arrmul12_ha0_8_y1;
  assign f_u_arrmul12_fa1_8_y3 = f_u_arrmul12_fa1_8_y0 & f_u_arrmul12_fa1_8_f_u_arrmul12_ha0_8_y1;
  assign f_u_arrmul12_fa1_8_y4 = f_u_arrmul12_fa1_8_y1 | f_u_arrmul12_fa1_8_y3;
  assign f_u_arrmul12_and2_8_a_2 = a_2;
  assign f_u_arrmul12_and2_8_b_8 = b_8;
  assign f_u_arrmul12_and2_8_y0 = f_u_arrmul12_and2_8_a_2 & f_u_arrmul12_and2_8_b_8;
  assign f_u_arrmul12_fa2_8_f_u_arrmul12_and2_8_y0 = f_u_arrmul12_and2_8_y0;
  assign f_u_arrmul12_fa2_8_f_u_arrmul12_fa3_7_y2 = f_u_arrmul12_fa3_7_y2;
  assign f_u_arrmul12_fa2_8_f_u_arrmul12_fa1_8_y4 = f_u_arrmul12_fa1_8_y4;
  assign f_u_arrmul12_fa2_8_y0 = f_u_arrmul12_fa2_8_f_u_arrmul12_and2_8_y0 ^ f_u_arrmul12_fa2_8_f_u_arrmul12_fa3_7_y2;
  assign f_u_arrmul12_fa2_8_y1 = f_u_arrmul12_fa2_8_f_u_arrmul12_and2_8_y0 & f_u_arrmul12_fa2_8_f_u_arrmul12_fa3_7_y2;
  assign f_u_arrmul12_fa2_8_y2 = f_u_arrmul12_fa2_8_y0 ^ f_u_arrmul12_fa2_8_f_u_arrmul12_fa1_8_y4;
  assign f_u_arrmul12_fa2_8_y3 = f_u_arrmul12_fa2_8_y0 & f_u_arrmul12_fa2_8_f_u_arrmul12_fa1_8_y4;
  assign f_u_arrmul12_fa2_8_y4 = f_u_arrmul12_fa2_8_y1 | f_u_arrmul12_fa2_8_y3;
  assign f_u_arrmul12_and3_8_a_3 = a_3;
  assign f_u_arrmul12_and3_8_b_8 = b_8;
  assign f_u_arrmul12_and3_8_y0 = f_u_arrmul12_and3_8_a_3 & f_u_arrmul12_and3_8_b_8;
  assign f_u_arrmul12_fa3_8_f_u_arrmul12_and3_8_y0 = f_u_arrmul12_and3_8_y0;
  assign f_u_arrmul12_fa3_8_f_u_arrmul12_fa4_7_y2 = f_u_arrmul12_fa4_7_y2;
  assign f_u_arrmul12_fa3_8_f_u_arrmul12_fa2_8_y4 = f_u_arrmul12_fa2_8_y4;
  assign f_u_arrmul12_fa3_8_y0 = f_u_arrmul12_fa3_8_f_u_arrmul12_and3_8_y0 ^ f_u_arrmul12_fa3_8_f_u_arrmul12_fa4_7_y2;
  assign f_u_arrmul12_fa3_8_y1 = f_u_arrmul12_fa3_8_f_u_arrmul12_and3_8_y0 & f_u_arrmul12_fa3_8_f_u_arrmul12_fa4_7_y2;
  assign f_u_arrmul12_fa3_8_y2 = f_u_arrmul12_fa3_8_y0 ^ f_u_arrmul12_fa3_8_f_u_arrmul12_fa2_8_y4;
  assign f_u_arrmul12_fa3_8_y3 = f_u_arrmul12_fa3_8_y0 & f_u_arrmul12_fa3_8_f_u_arrmul12_fa2_8_y4;
  assign f_u_arrmul12_fa3_8_y4 = f_u_arrmul12_fa3_8_y1 | f_u_arrmul12_fa3_8_y3;
  assign f_u_arrmul12_and4_8_a_4 = a_4;
  assign f_u_arrmul12_and4_8_b_8 = b_8;
  assign f_u_arrmul12_and4_8_y0 = f_u_arrmul12_and4_8_a_4 & f_u_arrmul12_and4_8_b_8;
  assign f_u_arrmul12_fa4_8_f_u_arrmul12_and4_8_y0 = f_u_arrmul12_and4_8_y0;
  assign f_u_arrmul12_fa4_8_f_u_arrmul12_fa5_7_y2 = f_u_arrmul12_fa5_7_y2;
  assign f_u_arrmul12_fa4_8_f_u_arrmul12_fa3_8_y4 = f_u_arrmul12_fa3_8_y4;
  assign f_u_arrmul12_fa4_8_y0 = f_u_arrmul12_fa4_8_f_u_arrmul12_and4_8_y0 ^ f_u_arrmul12_fa4_8_f_u_arrmul12_fa5_7_y2;
  assign f_u_arrmul12_fa4_8_y1 = f_u_arrmul12_fa4_8_f_u_arrmul12_and4_8_y0 & f_u_arrmul12_fa4_8_f_u_arrmul12_fa5_7_y2;
  assign f_u_arrmul12_fa4_8_y2 = f_u_arrmul12_fa4_8_y0 ^ f_u_arrmul12_fa4_8_f_u_arrmul12_fa3_8_y4;
  assign f_u_arrmul12_fa4_8_y3 = f_u_arrmul12_fa4_8_y0 & f_u_arrmul12_fa4_8_f_u_arrmul12_fa3_8_y4;
  assign f_u_arrmul12_fa4_8_y4 = f_u_arrmul12_fa4_8_y1 | f_u_arrmul12_fa4_8_y3;
  assign f_u_arrmul12_and5_8_a_5 = a_5;
  assign f_u_arrmul12_and5_8_b_8 = b_8;
  assign f_u_arrmul12_and5_8_y0 = f_u_arrmul12_and5_8_a_5 & f_u_arrmul12_and5_8_b_8;
  assign f_u_arrmul12_fa5_8_f_u_arrmul12_and5_8_y0 = f_u_arrmul12_and5_8_y0;
  assign f_u_arrmul12_fa5_8_f_u_arrmul12_fa6_7_y2 = f_u_arrmul12_fa6_7_y2;
  assign f_u_arrmul12_fa5_8_f_u_arrmul12_fa4_8_y4 = f_u_arrmul12_fa4_8_y4;
  assign f_u_arrmul12_fa5_8_y0 = f_u_arrmul12_fa5_8_f_u_arrmul12_and5_8_y0 ^ f_u_arrmul12_fa5_8_f_u_arrmul12_fa6_7_y2;
  assign f_u_arrmul12_fa5_8_y1 = f_u_arrmul12_fa5_8_f_u_arrmul12_and5_8_y0 & f_u_arrmul12_fa5_8_f_u_arrmul12_fa6_7_y2;
  assign f_u_arrmul12_fa5_8_y2 = f_u_arrmul12_fa5_8_y0 ^ f_u_arrmul12_fa5_8_f_u_arrmul12_fa4_8_y4;
  assign f_u_arrmul12_fa5_8_y3 = f_u_arrmul12_fa5_8_y0 & f_u_arrmul12_fa5_8_f_u_arrmul12_fa4_8_y4;
  assign f_u_arrmul12_fa5_8_y4 = f_u_arrmul12_fa5_8_y1 | f_u_arrmul12_fa5_8_y3;
  assign f_u_arrmul12_and6_8_a_6 = a_6;
  assign f_u_arrmul12_and6_8_b_8 = b_8;
  assign f_u_arrmul12_and6_8_y0 = f_u_arrmul12_and6_8_a_6 & f_u_arrmul12_and6_8_b_8;
  assign f_u_arrmul12_fa6_8_f_u_arrmul12_and6_8_y0 = f_u_arrmul12_and6_8_y0;
  assign f_u_arrmul12_fa6_8_f_u_arrmul12_fa7_7_y2 = f_u_arrmul12_fa7_7_y2;
  assign f_u_arrmul12_fa6_8_f_u_arrmul12_fa5_8_y4 = f_u_arrmul12_fa5_8_y4;
  assign f_u_arrmul12_fa6_8_y0 = f_u_arrmul12_fa6_8_f_u_arrmul12_and6_8_y0 ^ f_u_arrmul12_fa6_8_f_u_arrmul12_fa7_7_y2;
  assign f_u_arrmul12_fa6_8_y1 = f_u_arrmul12_fa6_8_f_u_arrmul12_and6_8_y0 & f_u_arrmul12_fa6_8_f_u_arrmul12_fa7_7_y2;
  assign f_u_arrmul12_fa6_8_y2 = f_u_arrmul12_fa6_8_y0 ^ f_u_arrmul12_fa6_8_f_u_arrmul12_fa5_8_y4;
  assign f_u_arrmul12_fa6_8_y3 = f_u_arrmul12_fa6_8_y0 & f_u_arrmul12_fa6_8_f_u_arrmul12_fa5_8_y4;
  assign f_u_arrmul12_fa6_8_y4 = f_u_arrmul12_fa6_8_y1 | f_u_arrmul12_fa6_8_y3;
  assign f_u_arrmul12_and7_8_a_7 = a_7;
  assign f_u_arrmul12_and7_8_b_8 = b_8;
  assign f_u_arrmul12_and7_8_y0 = f_u_arrmul12_and7_8_a_7 & f_u_arrmul12_and7_8_b_8;
  assign f_u_arrmul12_fa7_8_f_u_arrmul12_and7_8_y0 = f_u_arrmul12_and7_8_y0;
  assign f_u_arrmul12_fa7_8_f_u_arrmul12_fa8_7_y2 = f_u_arrmul12_fa8_7_y2;
  assign f_u_arrmul12_fa7_8_f_u_arrmul12_fa6_8_y4 = f_u_arrmul12_fa6_8_y4;
  assign f_u_arrmul12_fa7_8_y0 = f_u_arrmul12_fa7_8_f_u_arrmul12_and7_8_y0 ^ f_u_arrmul12_fa7_8_f_u_arrmul12_fa8_7_y2;
  assign f_u_arrmul12_fa7_8_y1 = f_u_arrmul12_fa7_8_f_u_arrmul12_and7_8_y0 & f_u_arrmul12_fa7_8_f_u_arrmul12_fa8_7_y2;
  assign f_u_arrmul12_fa7_8_y2 = f_u_arrmul12_fa7_8_y0 ^ f_u_arrmul12_fa7_8_f_u_arrmul12_fa6_8_y4;
  assign f_u_arrmul12_fa7_8_y3 = f_u_arrmul12_fa7_8_y0 & f_u_arrmul12_fa7_8_f_u_arrmul12_fa6_8_y4;
  assign f_u_arrmul12_fa7_8_y4 = f_u_arrmul12_fa7_8_y1 | f_u_arrmul12_fa7_8_y3;
  assign f_u_arrmul12_and8_8_a_8 = a_8;
  assign f_u_arrmul12_and8_8_b_8 = b_8;
  assign f_u_arrmul12_and8_8_y0 = f_u_arrmul12_and8_8_a_8 & f_u_arrmul12_and8_8_b_8;
  assign f_u_arrmul12_fa8_8_f_u_arrmul12_and8_8_y0 = f_u_arrmul12_and8_8_y0;
  assign f_u_arrmul12_fa8_8_f_u_arrmul12_fa9_7_y2 = f_u_arrmul12_fa9_7_y2;
  assign f_u_arrmul12_fa8_8_f_u_arrmul12_fa7_8_y4 = f_u_arrmul12_fa7_8_y4;
  assign f_u_arrmul12_fa8_8_y0 = f_u_arrmul12_fa8_8_f_u_arrmul12_and8_8_y0 ^ f_u_arrmul12_fa8_8_f_u_arrmul12_fa9_7_y2;
  assign f_u_arrmul12_fa8_8_y1 = f_u_arrmul12_fa8_8_f_u_arrmul12_and8_8_y0 & f_u_arrmul12_fa8_8_f_u_arrmul12_fa9_7_y2;
  assign f_u_arrmul12_fa8_8_y2 = f_u_arrmul12_fa8_8_y0 ^ f_u_arrmul12_fa8_8_f_u_arrmul12_fa7_8_y4;
  assign f_u_arrmul12_fa8_8_y3 = f_u_arrmul12_fa8_8_y0 & f_u_arrmul12_fa8_8_f_u_arrmul12_fa7_8_y4;
  assign f_u_arrmul12_fa8_8_y4 = f_u_arrmul12_fa8_8_y1 | f_u_arrmul12_fa8_8_y3;
  assign f_u_arrmul12_and9_8_a_9 = a_9;
  assign f_u_arrmul12_and9_8_b_8 = b_8;
  assign f_u_arrmul12_and9_8_y0 = f_u_arrmul12_and9_8_a_9 & f_u_arrmul12_and9_8_b_8;
  assign f_u_arrmul12_fa9_8_f_u_arrmul12_and9_8_y0 = f_u_arrmul12_and9_8_y0;
  assign f_u_arrmul12_fa9_8_f_u_arrmul12_fa10_7_y2 = f_u_arrmul12_fa10_7_y2;
  assign f_u_arrmul12_fa9_8_f_u_arrmul12_fa8_8_y4 = f_u_arrmul12_fa8_8_y4;
  assign f_u_arrmul12_fa9_8_y0 = f_u_arrmul12_fa9_8_f_u_arrmul12_and9_8_y0 ^ f_u_arrmul12_fa9_8_f_u_arrmul12_fa10_7_y2;
  assign f_u_arrmul12_fa9_8_y1 = f_u_arrmul12_fa9_8_f_u_arrmul12_and9_8_y0 & f_u_arrmul12_fa9_8_f_u_arrmul12_fa10_7_y2;
  assign f_u_arrmul12_fa9_8_y2 = f_u_arrmul12_fa9_8_y0 ^ f_u_arrmul12_fa9_8_f_u_arrmul12_fa8_8_y4;
  assign f_u_arrmul12_fa9_8_y3 = f_u_arrmul12_fa9_8_y0 & f_u_arrmul12_fa9_8_f_u_arrmul12_fa8_8_y4;
  assign f_u_arrmul12_fa9_8_y4 = f_u_arrmul12_fa9_8_y1 | f_u_arrmul12_fa9_8_y3;
  assign f_u_arrmul12_and10_8_a_10 = a_10;
  assign f_u_arrmul12_and10_8_b_8 = b_8;
  assign f_u_arrmul12_and10_8_y0 = f_u_arrmul12_and10_8_a_10 & f_u_arrmul12_and10_8_b_8;
  assign f_u_arrmul12_fa10_8_f_u_arrmul12_and10_8_y0 = f_u_arrmul12_and10_8_y0;
  assign f_u_arrmul12_fa10_8_f_u_arrmul12_fa11_7_y2 = f_u_arrmul12_fa11_7_y2;
  assign f_u_arrmul12_fa10_8_f_u_arrmul12_fa9_8_y4 = f_u_arrmul12_fa9_8_y4;
  assign f_u_arrmul12_fa10_8_y0 = f_u_arrmul12_fa10_8_f_u_arrmul12_and10_8_y0 ^ f_u_arrmul12_fa10_8_f_u_arrmul12_fa11_7_y2;
  assign f_u_arrmul12_fa10_8_y1 = f_u_arrmul12_fa10_8_f_u_arrmul12_and10_8_y0 & f_u_arrmul12_fa10_8_f_u_arrmul12_fa11_7_y2;
  assign f_u_arrmul12_fa10_8_y2 = f_u_arrmul12_fa10_8_y0 ^ f_u_arrmul12_fa10_8_f_u_arrmul12_fa9_8_y4;
  assign f_u_arrmul12_fa10_8_y3 = f_u_arrmul12_fa10_8_y0 & f_u_arrmul12_fa10_8_f_u_arrmul12_fa9_8_y4;
  assign f_u_arrmul12_fa10_8_y4 = f_u_arrmul12_fa10_8_y1 | f_u_arrmul12_fa10_8_y3;
  assign f_u_arrmul12_and11_8_a_11 = a_11;
  assign f_u_arrmul12_and11_8_b_8 = b_8;
  assign f_u_arrmul12_and11_8_y0 = f_u_arrmul12_and11_8_a_11 & f_u_arrmul12_and11_8_b_8;
  assign f_u_arrmul12_fa11_8_f_u_arrmul12_and11_8_y0 = f_u_arrmul12_and11_8_y0;
  assign f_u_arrmul12_fa11_8_f_u_arrmul12_fa11_7_y4 = f_u_arrmul12_fa11_7_y4;
  assign f_u_arrmul12_fa11_8_f_u_arrmul12_fa10_8_y4 = f_u_arrmul12_fa10_8_y4;
  assign f_u_arrmul12_fa11_8_y0 = f_u_arrmul12_fa11_8_f_u_arrmul12_and11_8_y0 ^ f_u_arrmul12_fa11_8_f_u_arrmul12_fa11_7_y4;
  assign f_u_arrmul12_fa11_8_y1 = f_u_arrmul12_fa11_8_f_u_arrmul12_and11_8_y0 & f_u_arrmul12_fa11_8_f_u_arrmul12_fa11_7_y4;
  assign f_u_arrmul12_fa11_8_y2 = f_u_arrmul12_fa11_8_y0 ^ f_u_arrmul12_fa11_8_f_u_arrmul12_fa10_8_y4;
  assign f_u_arrmul12_fa11_8_y3 = f_u_arrmul12_fa11_8_y0 & f_u_arrmul12_fa11_8_f_u_arrmul12_fa10_8_y4;
  assign f_u_arrmul12_fa11_8_y4 = f_u_arrmul12_fa11_8_y1 | f_u_arrmul12_fa11_8_y3;
  assign f_u_arrmul12_and0_9_a_0 = a_0;
  assign f_u_arrmul12_and0_9_b_9 = b_9;
  assign f_u_arrmul12_and0_9_y0 = f_u_arrmul12_and0_9_a_0 & f_u_arrmul12_and0_9_b_9;
  assign f_u_arrmul12_ha0_9_f_u_arrmul12_and0_9_y0 = f_u_arrmul12_and0_9_y0;
  assign f_u_arrmul12_ha0_9_f_u_arrmul12_fa1_8_y2 = f_u_arrmul12_fa1_8_y2;
  assign f_u_arrmul12_ha0_9_y0 = f_u_arrmul12_ha0_9_f_u_arrmul12_and0_9_y0 ^ f_u_arrmul12_ha0_9_f_u_arrmul12_fa1_8_y2;
  assign f_u_arrmul12_ha0_9_y1 = f_u_arrmul12_ha0_9_f_u_arrmul12_and0_9_y0 & f_u_arrmul12_ha0_9_f_u_arrmul12_fa1_8_y2;
  assign f_u_arrmul12_and1_9_a_1 = a_1;
  assign f_u_arrmul12_and1_9_b_9 = b_9;
  assign f_u_arrmul12_and1_9_y0 = f_u_arrmul12_and1_9_a_1 & f_u_arrmul12_and1_9_b_9;
  assign f_u_arrmul12_fa1_9_f_u_arrmul12_and1_9_y0 = f_u_arrmul12_and1_9_y0;
  assign f_u_arrmul12_fa1_9_f_u_arrmul12_fa2_8_y2 = f_u_arrmul12_fa2_8_y2;
  assign f_u_arrmul12_fa1_9_f_u_arrmul12_ha0_9_y1 = f_u_arrmul12_ha0_9_y1;
  assign f_u_arrmul12_fa1_9_y0 = f_u_arrmul12_fa1_9_f_u_arrmul12_and1_9_y0 ^ f_u_arrmul12_fa1_9_f_u_arrmul12_fa2_8_y2;
  assign f_u_arrmul12_fa1_9_y1 = f_u_arrmul12_fa1_9_f_u_arrmul12_and1_9_y0 & f_u_arrmul12_fa1_9_f_u_arrmul12_fa2_8_y2;
  assign f_u_arrmul12_fa1_9_y2 = f_u_arrmul12_fa1_9_y0 ^ f_u_arrmul12_fa1_9_f_u_arrmul12_ha0_9_y1;
  assign f_u_arrmul12_fa1_9_y3 = f_u_arrmul12_fa1_9_y0 & f_u_arrmul12_fa1_9_f_u_arrmul12_ha0_9_y1;
  assign f_u_arrmul12_fa1_9_y4 = f_u_arrmul12_fa1_9_y1 | f_u_arrmul12_fa1_9_y3;
  assign f_u_arrmul12_and2_9_a_2 = a_2;
  assign f_u_arrmul12_and2_9_b_9 = b_9;
  assign f_u_arrmul12_and2_9_y0 = f_u_arrmul12_and2_9_a_2 & f_u_arrmul12_and2_9_b_9;
  assign f_u_arrmul12_fa2_9_f_u_arrmul12_and2_9_y0 = f_u_arrmul12_and2_9_y0;
  assign f_u_arrmul12_fa2_9_f_u_arrmul12_fa3_8_y2 = f_u_arrmul12_fa3_8_y2;
  assign f_u_arrmul12_fa2_9_f_u_arrmul12_fa1_9_y4 = f_u_arrmul12_fa1_9_y4;
  assign f_u_arrmul12_fa2_9_y0 = f_u_arrmul12_fa2_9_f_u_arrmul12_and2_9_y0 ^ f_u_arrmul12_fa2_9_f_u_arrmul12_fa3_8_y2;
  assign f_u_arrmul12_fa2_9_y1 = f_u_arrmul12_fa2_9_f_u_arrmul12_and2_9_y0 & f_u_arrmul12_fa2_9_f_u_arrmul12_fa3_8_y2;
  assign f_u_arrmul12_fa2_9_y2 = f_u_arrmul12_fa2_9_y0 ^ f_u_arrmul12_fa2_9_f_u_arrmul12_fa1_9_y4;
  assign f_u_arrmul12_fa2_9_y3 = f_u_arrmul12_fa2_9_y0 & f_u_arrmul12_fa2_9_f_u_arrmul12_fa1_9_y4;
  assign f_u_arrmul12_fa2_9_y4 = f_u_arrmul12_fa2_9_y1 | f_u_arrmul12_fa2_9_y3;
  assign f_u_arrmul12_and3_9_a_3 = a_3;
  assign f_u_arrmul12_and3_9_b_9 = b_9;
  assign f_u_arrmul12_and3_9_y0 = f_u_arrmul12_and3_9_a_3 & f_u_arrmul12_and3_9_b_9;
  assign f_u_arrmul12_fa3_9_f_u_arrmul12_and3_9_y0 = f_u_arrmul12_and3_9_y0;
  assign f_u_arrmul12_fa3_9_f_u_arrmul12_fa4_8_y2 = f_u_arrmul12_fa4_8_y2;
  assign f_u_arrmul12_fa3_9_f_u_arrmul12_fa2_9_y4 = f_u_arrmul12_fa2_9_y4;
  assign f_u_arrmul12_fa3_9_y0 = f_u_arrmul12_fa3_9_f_u_arrmul12_and3_9_y0 ^ f_u_arrmul12_fa3_9_f_u_arrmul12_fa4_8_y2;
  assign f_u_arrmul12_fa3_9_y1 = f_u_arrmul12_fa3_9_f_u_arrmul12_and3_9_y0 & f_u_arrmul12_fa3_9_f_u_arrmul12_fa4_8_y2;
  assign f_u_arrmul12_fa3_9_y2 = f_u_arrmul12_fa3_9_y0 ^ f_u_arrmul12_fa3_9_f_u_arrmul12_fa2_9_y4;
  assign f_u_arrmul12_fa3_9_y3 = f_u_arrmul12_fa3_9_y0 & f_u_arrmul12_fa3_9_f_u_arrmul12_fa2_9_y4;
  assign f_u_arrmul12_fa3_9_y4 = f_u_arrmul12_fa3_9_y1 | f_u_arrmul12_fa3_9_y3;
  assign f_u_arrmul12_and4_9_a_4 = a_4;
  assign f_u_arrmul12_and4_9_b_9 = b_9;
  assign f_u_arrmul12_and4_9_y0 = f_u_arrmul12_and4_9_a_4 & f_u_arrmul12_and4_9_b_9;
  assign f_u_arrmul12_fa4_9_f_u_arrmul12_and4_9_y0 = f_u_arrmul12_and4_9_y0;
  assign f_u_arrmul12_fa4_9_f_u_arrmul12_fa5_8_y2 = f_u_arrmul12_fa5_8_y2;
  assign f_u_arrmul12_fa4_9_f_u_arrmul12_fa3_9_y4 = f_u_arrmul12_fa3_9_y4;
  assign f_u_arrmul12_fa4_9_y0 = f_u_arrmul12_fa4_9_f_u_arrmul12_and4_9_y0 ^ f_u_arrmul12_fa4_9_f_u_arrmul12_fa5_8_y2;
  assign f_u_arrmul12_fa4_9_y1 = f_u_arrmul12_fa4_9_f_u_arrmul12_and4_9_y0 & f_u_arrmul12_fa4_9_f_u_arrmul12_fa5_8_y2;
  assign f_u_arrmul12_fa4_9_y2 = f_u_arrmul12_fa4_9_y0 ^ f_u_arrmul12_fa4_9_f_u_arrmul12_fa3_9_y4;
  assign f_u_arrmul12_fa4_9_y3 = f_u_arrmul12_fa4_9_y0 & f_u_arrmul12_fa4_9_f_u_arrmul12_fa3_9_y4;
  assign f_u_arrmul12_fa4_9_y4 = f_u_arrmul12_fa4_9_y1 | f_u_arrmul12_fa4_9_y3;
  assign f_u_arrmul12_and5_9_a_5 = a_5;
  assign f_u_arrmul12_and5_9_b_9 = b_9;
  assign f_u_arrmul12_and5_9_y0 = f_u_arrmul12_and5_9_a_5 & f_u_arrmul12_and5_9_b_9;
  assign f_u_arrmul12_fa5_9_f_u_arrmul12_and5_9_y0 = f_u_arrmul12_and5_9_y0;
  assign f_u_arrmul12_fa5_9_f_u_arrmul12_fa6_8_y2 = f_u_arrmul12_fa6_8_y2;
  assign f_u_arrmul12_fa5_9_f_u_arrmul12_fa4_9_y4 = f_u_arrmul12_fa4_9_y4;
  assign f_u_arrmul12_fa5_9_y0 = f_u_arrmul12_fa5_9_f_u_arrmul12_and5_9_y0 ^ f_u_arrmul12_fa5_9_f_u_arrmul12_fa6_8_y2;
  assign f_u_arrmul12_fa5_9_y1 = f_u_arrmul12_fa5_9_f_u_arrmul12_and5_9_y0 & f_u_arrmul12_fa5_9_f_u_arrmul12_fa6_8_y2;
  assign f_u_arrmul12_fa5_9_y2 = f_u_arrmul12_fa5_9_y0 ^ f_u_arrmul12_fa5_9_f_u_arrmul12_fa4_9_y4;
  assign f_u_arrmul12_fa5_9_y3 = f_u_arrmul12_fa5_9_y0 & f_u_arrmul12_fa5_9_f_u_arrmul12_fa4_9_y4;
  assign f_u_arrmul12_fa5_9_y4 = f_u_arrmul12_fa5_9_y1 | f_u_arrmul12_fa5_9_y3;
  assign f_u_arrmul12_and6_9_a_6 = a_6;
  assign f_u_arrmul12_and6_9_b_9 = b_9;
  assign f_u_arrmul12_and6_9_y0 = f_u_arrmul12_and6_9_a_6 & f_u_arrmul12_and6_9_b_9;
  assign f_u_arrmul12_fa6_9_f_u_arrmul12_and6_9_y0 = f_u_arrmul12_and6_9_y0;
  assign f_u_arrmul12_fa6_9_f_u_arrmul12_fa7_8_y2 = f_u_arrmul12_fa7_8_y2;
  assign f_u_arrmul12_fa6_9_f_u_arrmul12_fa5_9_y4 = f_u_arrmul12_fa5_9_y4;
  assign f_u_arrmul12_fa6_9_y0 = f_u_arrmul12_fa6_9_f_u_arrmul12_and6_9_y0 ^ f_u_arrmul12_fa6_9_f_u_arrmul12_fa7_8_y2;
  assign f_u_arrmul12_fa6_9_y1 = f_u_arrmul12_fa6_9_f_u_arrmul12_and6_9_y0 & f_u_arrmul12_fa6_9_f_u_arrmul12_fa7_8_y2;
  assign f_u_arrmul12_fa6_9_y2 = f_u_arrmul12_fa6_9_y0 ^ f_u_arrmul12_fa6_9_f_u_arrmul12_fa5_9_y4;
  assign f_u_arrmul12_fa6_9_y3 = f_u_arrmul12_fa6_9_y0 & f_u_arrmul12_fa6_9_f_u_arrmul12_fa5_9_y4;
  assign f_u_arrmul12_fa6_9_y4 = f_u_arrmul12_fa6_9_y1 | f_u_arrmul12_fa6_9_y3;
  assign f_u_arrmul12_and7_9_a_7 = a_7;
  assign f_u_arrmul12_and7_9_b_9 = b_9;
  assign f_u_arrmul12_and7_9_y0 = f_u_arrmul12_and7_9_a_7 & f_u_arrmul12_and7_9_b_9;
  assign f_u_arrmul12_fa7_9_f_u_arrmul12_and7_9_y0 = f_u_arrmul12_and7_9_y0;
  assign f_u_arrmul12_fa7_9_f_u_arrmul12_fa8_8_y2 = f_u_arrmul12_fa8_8_y2;
  assign f_u_arrmul12_fa7_9_f_u_arrmul12_fa6_9_y4 = f_u_arrmul12_fa6_9_y4;
  assign f_u_arrmul12_fa7_9_y0 = f_u_arrmul12_fa7_9_f_u_arrmul12_and7_9_y0 ^ f_u_arrmul12_fa7_9_f_u_arrmul12_fa8_8_y2;
  assign f_u_arrmul12_fa7_9_y1 = f_u_arrmul12_fa7_9_f_u_arrmul12_and7_9_y0 & f_u_arrmul12_fa7_9_f_u_arrmul12_fa8_8_y2;
  assign f_u_arrmul12_fa7_9_y2 = f_u_arrmul12_fa7_9_y0 ^ f_u_arrmul12_fa7_9_f_u_arrmul12_fa6_9_y4;
  assign f_u_arrmul12_fa7_9_y3 = f_u_arrmul12_fa7_9_y0 & f_u_arrmul12_fa7_9_f_u_arrmul12_fa6_9_y4;
  assign f_u_arrmul12_fa7_9_y4 = f_u_arrmul12_fa7_9_y1 | f_u_arrmul12_fa7_9_y3;
  assign f_u_arrmul12_and8_9_a_8 = a_8;
  assign f_u_arrmul12_and8_9_b_9 = b_9;
  assign f_u_arrmul12_and8_9_y0 = f_u_arrmul12_and8_9_a_8 & f_u_arrmul12_and8_9_b_9;
  assign f_u_arrmul12_fa8_9_f_u_arrmul12_and8_9_y0 = f_u_arrmul12_and8_9_y0;
  assign f_u_arrmul12_fa8_9_f_u_arrmul12_fa9_8_y2 = f_u_arrmul12_fa9_8_y2;
  assign f_u_arrmul12_fa8_9_f_u_arrmul12_fa7_9_y4 = f_u_arrmul12_fa7_9_y4;
  assign f_u_arrmul12_fa8_9_y0 = f_u_arrmul12_fa8_9_f_u_arrmul12_and8_9_y0 ^ f_u_arrmul12_fa8_9_f_u_arrmul12_fa9_8_y2;
  assign f_u_arrmul12_fa8_9_y1 = f_u_arrmul12_fa8_9_f_u_arrmul12_and8_9_y0 & f_u_arrmul12_fa8_9_f_u_arrmul12_fa9_8_y2;
  assign f_u_arrmul12_fa8_9_y2 = f_u_arrmul12_fa8_9_y0 ^ f_u_arrmul12_fa8_9_f_u_arrmul12_fa7_9_y4;
  assign f_u_arrmul12_fa8_9_y3 = f_u_arrmul12_fa8_9_y0 & f_u_arrmul12_fa8_9_f_u_arrmul12_fa7_9_y4;
  assign f_u_arrmul12_fa8_9_y4 = f_u_arrmul12_fa8_9_y1 | f_u_arrmul12_fa8_9_y3;
  assign f_u_arrmul12_and9_9_a_9 = a_9;
  assign f_u_arrmul12_and9_9_b_9 = b_9;
  assign f_u_arrmul12_and9_9_y0 = f_u_arrmul12_and9_9_a_9 & f_u_arrmul12_and9_9_b_9;
  assign f_u_arrmul12_fa9_9_f_u_arrmul12_and9_9_y0 = f_u_arrmul12_and9_9_y0;
  assign f_u_arrmul12_fa9_9_f_u_arrmul12_fa10_8_y2 = f_u_arrmul12_fa10_8_y2;
  assign f_u_arrmul12_fa9_9_f_u_arrmul12_fa8_9_y4 = f_u_arrmul12_fa8_9_y4;
  assign f_u_arrmul12_fa9_9_y0 = f_u_arrmul12_fa9_9_f_u_arrmul12_and9_9_y0 ^ f_u_arrmul12_fa9_9_f_u_arrmul12_fa10_8_y2;
  assign f_u_arrmul12_fa9_9_y1 = f_u_arrmul12_fa9_9_f_u_arrmul12_and9_9_y0 & f_u_arrmul12_fa9_9_f_u_arrmul12_fa10_8_y2;
  assign f_u_arrmul12_fa9_9_y2 = f_u_arrmul12_fa9_9_y0 ^ f_u_arrmul12_fa9_9_f_u_arrmul12_fa8_9_y4;
  assign f_u_arrmul12_fa9_9_y3 = f_u_arrmul12_fa9_9_y0 & f_u_arrmul12_fa9_9_f_u_arrmul12_fa8_9_y4;
  assign f_u_arrmul12_fa9_9_y4 = f_u_arrmul12_fa9_9_y1 | f_u_arrmul12_fa9_9_y3;
  assign f_u_arrmul12_and10_9_a_10 = a_10;
  assign f_u_arrmul12_and10_9_b_9 = b_9;
  assign f_u_arrmul12_and10_9_y0 = f_u_arrmul12_and10_9_a_10 & f_u_arrmul12_and10_9_b_9;
  assign f_u_arrmul12_fa10_9_f_u_arrmul12_and10_9_y0 = f_u_arrmul12_and10_9_y0;
  assign f_u_arrmul12_fa10_9_f_u_arrmul12_fa11_8_y2 = f_u_arrmul12_fa11_8_y2;
  assign f_u_arrmul12_fa10_9_f_u_arrmul12_fa9_9_y4 = f_u_arrmul12_fa9_9_y4;
  assign f_u_arrmul12_fa10_9_y0 = f_u_arrmul12_fa10_9_f_u_arrmul12_and10_9_y0 ^ f_u_arrmul12_fa10_9_f_u_arrmul12_fa11_8_y2;
  assign f_u_arrmul12_fa10_9_y1 = f_u_arrmul12_fa10_9_f_u_arrmul12_and10_9_y0 & f_u_arrmul12_fa10_9_f_u_arrmul12_fa11_8_y2;
  assign f_u_arrmul12_fa10_9_y2 = f_u_arrmul12_fa10_9_y0 ^ f_u_arrmul12_fa10_9_f_u_arrmul12_fa9_9_y4;
  assign f_u_arrmul12_fa10_9_y3 = f_u_arrmul12_fa10_9_y0 & f_u_arrmul12_fa10_9_f_u_arrmul12_fa9_9_y4;
  assign f_u_arrmul12_fa10_9_y4 = f_u_arrmul12_fa10_9_y1 | f_u_arrmul12_fa10_9_y3;
  assign f_u_arrmul12_and11_9_a_11 = a_11;
  assign f_u_arrmul12_and11_9_b_9 = b_9;
  assign f_u_arrmul12_and11_9_y0 = f_u_arrmul12_and11_9_a_11 & f_u_arrmul12_and11_9_b_9;
  assign f_u_arrmul12_fa11_9_f_u_arrmul12_and11_9_y0 = f_u_arrmul12_and11_9_y0;
  assign f_u_arrmul12_fa11_9_f_u_arrmul12_fa11_8_y4 = f_u_arrmul12_fa11_8_y4;
  assign f_u_arrmul12_fa11_9_f_u_arrmul12_fa10_9_y4 = f_u_arrmul12_fa10_9_y4;
  assign f_u_arrmul12_fa11_9_y0 = f_u_arrmul12_fa11_9_f_u_arrmul12_and11_9_y0 ^ f_u_arrmul12_fa11_9_f_u_arrmul12_fa11_8_y4;
  assign f_u_arrmul12_fa11_9_y1 = f_u_arrmul12_fa11_9_f_u_arrmul12_and11_9_y0 & f_u_arrmul12_fa11_9_f_u_arrmul12_fa11_8_y4;
  assign f_u_arrmul12_fa11_9_y2 = f_u_arrmul12_fa11_9_y0 ^ f_u_arrmul12_fa11_9_f_u_arrmul12_fa10_9_y4;
  assign f_u_arrmul12_fa11_9_y3 = f_u_arrmul12_fa11_9_y0 & f_u_arrmul12_fa11_9_f_u_arrmul12_fa10_9_y4;
  assign f_u_arrmul12_fa11_9_y4 = f_u_arrmul12_fa11_9_y1 | f_u_arrmul12_fa11_9_y3;
  assign f_u_arrmul12_and0_10_a_0 = a_0;
  assign f_u_arrmul12_and0_10_b_10 = b_10;
  assign f_u_arrmul12_and0_10_y0 = f_u_arrmul12_and0_10_a_0 & f_u_arrmul12_and0_10_b_10;
  assign f_u_arrmul12_ha0_10_f_u_arrmul12_and0_10_y0 = f_u_arrmul12_and0_10_y0;
  assign f_u_arrmul12_ha0_10_f_u_arrmul12_fa1_9_y2 = f_u_arrmul12_fa1_9_y2;
  assign f_u_arrmul12_ha0_10_y0 = f_u_arrmul12_ha0_10_f_u_arrmul12_and0_10_y0 ^ f_u_arrmul12_ha0_10_f_u_arrmul12_fa1_9_y2;
  assign f_u_arrmul12_ha0_10_y1 = f_u_arrmul12_ha0_10_f_u_arrmul12_and0_10_y0 & f_u_arrmul12_ha0_10_f_u_arrmul12_fa1_9_y2;
  assign f_u_arrmul12_and1_10_a_1 = a_1;
  assign f_u_arrmul12_and1_10_b_10 = b_10;
  assign f_u_arrmul12_and1_10_y0 = f_u_arrmul12_and1_10_a_1 & f_u_arrmul12_and1_10_b_10;
  assign f_u_arrmul12_fa1_10_f_u_arrmul12_and1_10_y0 = f_u_arrmul12_and1_10_y0;
  assign f_u_arrmul12_fa1_10_f_u_arrmul12_fa2_9_y2 = f_u_arrmul12_fa2_9_y2;
  assign f_u_arrmul12_fa1_10_f_u_arrmul12_ha0_10_y1 = f_u_arrmul12_ha0_10_y1;
  assign f_u_arrmul12_fa1_10_y0 = f_u_arrmul12_fa1_10_f_u_arrmul12_and1_10_y0 ^ f_u_arrmul12_fa1_10_f_u_arrmul12_fa2_9_y2;
  assign f_u_arrmul12_fa1_10_y1 = f_u_arrmul12_fa1_10_f_u_arrmul12_and1_10_y0 & f_u_arrmul12_fa1_10_f_u_arrmul12_fa2_9_y2;
  assign f_u_arrmul12_fa1_10_y2 = f_u_arrmul12_fa1_10_y0 ^ f_u_arrmul12_fa1_10_f_u_arrmul12_ha0_10_y1;
  assign f_u_arrmul12_fa1_10_y3 = f_u_arrmul12_fa1_10_y0 & f_u_arrmul12_fa1_10_f_u_arrmul12_ha0_10_y1;
  assign f_u_arrmul12_fa1_10_y4 = f_u_arrmul12_fa1_10_y1 | f_u_arrmul12_fa1_10_y3;
  assign f_u_arrmul12_and2_10_a_2 = a_2;
  assign f_u_arrmul12_and2_10_b_10 = b_10;
  assign f_u_arrmul12_and2_10_y0 = f_u_arrmul12_and2_10_a_2 & f_u_arrmul12_and2_10_b_10;
  assign f_u_arrmul12_fa2_10_f_u_arrmul12_and2_10_y0 = f_u_arrmul12_and2_10_y0;
  assign f_u_arrmul12_fa2_10_f_u_arrmul12_fa3_9_y2 = f_u_arrmul12_fa3_9_y2;
  assign f_u_arrmul12_fa2_10_f_u_arrmul12_fa1_10_y4 = f_u_arrmul12_fa1_10_y4;
  assign f_u_arrmul12_fa2_10_y0 = f_u_arrmul12_fa2_10_f_u_arrmul12_and2_10_y0 ^ f_u_arrmul12_fa2_10_f_u_arrmul12_fa3_9_y2;
  assign f_u_arrmul12_fa2_10_y1 = f_u_arrmul12_fa2_10_f_u_arrmul12_and2_10_y0 & f_u_arrmul12_fa2_10_f_u_arrmul12_fa3_9_y2;
  assign f_u_arrmul12_fa2_10_y2 = f_u_arrmul12_fa2_10_y0 ^ f_u_arrmul12_fa2_10_f_u_arrmul12_fa1_10_y4;
  assign f_u_arrmul12_fa2_10_y3 = f_u_arrmul12_fa2_10_y0 & f_u_arrmul12_fa2_10_f_u_arrmul12_fa1_10_y4;
  assign f_u_arrmul12_fa2_10_y4 = f_u_arrmul12_fa2_10_y1 | f_u_arrmul12_fa2_10_y3;
  assign f_u_arrmul12_and3_10_a_3 = a_3;
  assign f_u_arrmul12_and3_10_b_10 = b_10;
  assign f_u_arrmul12_and3_10_y0 = f_u_arrmul12_and3_10_a_3 & f_u_arrmul12_and3_10_b_10;
  assign f_u_arrmul12_fa3_10_f_u_arrmul12_and3_10_y0 = f_u_arrmul12_and3_10_y0;
  assign f_u_arrmul12_fa3_10_f_u_arrmul12_fa4_9_y2 = f_u_arrmul12_fa4_9_y2;
  assign f_u_arrmul12_fa3_10_f_u_arrmul12_fa2_10_y4 = f_u_arrmul12_fa2_10_y4;
  assign f_u_arrmul12_fa3_10_y0 = f_u_arrmul12_fa3_10_f_u_arrmul12_and3_10_y0 ^ f_u_arrmul12_fa3_10_f_u_arrmul12_fa4_9_y2;
  assign f_u_arrmul12_fa3_10_y1 = f_u_arrmul12_fa3_10_f_u_arrmul12_and3_10_y0 & f_u_arrmul12_fa3_10_f_u_arrmul12_fa4_9_y2;
  assign f_u_arrmul12_fa3_10_y2 = f_u_arrmul12_fa3_10_y0 ^ f_u_arrmul12_fa3_10_f_u_arrmul12_fa2_10_y4;
  assign f_u_arrmul12_fa3_10_y3 = f_u_arrmul12_fa3_10_y0 & f_u_arrmul12_fa3_10_f_u_arrmul12_fa2_10_y4;
  assign f_u_arrmul12_fa3_10_y4 = f_u_arrmul12_fa3_10_y1 | f_u_arrmul12_fa3_10_y3;
  assign f_u_arrmul12_and4_10_a_4 = a_4;
  assign f_u_arrmul12_and4_10_b_10 = b_10;
  assign f_u_arrmul12_and4_10_y0 = f_u_arrmul12_and4_10_a_4 & f_u_arrmul12_and4_10_b_10;
  assign f_u_arrmul12_fa4_10_f_u_arrmul12_and4_10_y0 = f_u_arrmul12_and4_10_y0;
  assign f_u_arrmul12_fa4_10_f_u_arrmul12_fa5_9_y2 = f_u_arrmul12_fa5_9_y2;
  assign f_u_arrmul12_fa4_10_f_u_arrmul12_fa3_10_y4 = f_u_arrmul12_fa3_10_y4;
  assign f_u_arrmul12_fa4_10_y0 = f_u_arrmul12_fa4_10_f_u_arrmul12_and4_10_y0 ^ f_u_arrmul12_fa4_10_f_u_arrmul12_fa5_9_y2;
  assign f_u_arrmul12_fa4_10_y1 = f_u_arrmul12_fa4_10_f_u_arrmul12_and4_10_y0 & f_u_arrmul12_fa4_10_f_u_arrmul12_fa5_9_y2;
  assign f_u_arrmul12_fa4_10_y2 = f_u_arrmul12_fa4_10_y0 ^ f_u_arrmul12_fa4_10_f_u_arrmul12_fa3_10_y4;
  assign f_u_arrmul12_fa4_10_y3 = f_u_arrmul12_fa4_10_y0 & f_u_arrmul12_fa4_10_f_u_arrmul12_fa3_10_y4;
  assign f_u_arrmul12_fa4_10_y4 = f_u_arrmul12_fa4_10_y1 | f_u_arrmul12_fa4_10_y3;
  assign f_u_arrmul12_and5_10_a_5 = a_5;
  assign f_u_arrmul12_and5_10_b_10 = b_10;
  assign f_u_arrmul12_and5_10_y0 = f_u_arrmul12_and5_10_a_5 & f_u_arrmul12_and5_10_b_10;
  assign f_u_arrmul12_fa5_10_f_u_arrmul12_and5_10_y0 = f_u_arrmul12_and5_10_y0;
  assign f_u_arrmul12_fa5_10_f_u_arrmul12_fa6_9_y2 = f_u_arrmul12_fa6_9_y2;
  assign f_u_arrmul12_fa5_10_f_u_arrmul12_fa4_10_y4 = f_u_arrmul12_fa4_10_y4;
  assign f_u_arrmul12_fa5_10_y0 = f_u_arrmul12_fa5_10_f_u_arrmul12_and5_10_y0 ^ f_u_arrmul12_fa5_10_f_u_arrmul12_fa6_9_y2;
  assign f_u_arrmul12_fa5_10_y1 = f_u_arrmul12_fa5_10_f_u_arrmul12_and5_10_y0 & f_u_arrmul12_fa5_10_f_u_arrmul12_fa6_9_y2;
  assign f_u_arrmul12_fa5_10_y2 = f_u_arrmul12_fa5_10_y0 ^ f_u_arrmul12_fa5_10_f_u_arrmul12_fa4_10_y4;
  assign f_u_arrmul12_fa5_10_y3 = f_u_arrmul12_fa5_10_y0 & f_u_arrmul12_fa5_10_f_u_arrmul12_fa4_10_y4;
  assign f_u_arrmul12_fa5_10_y4 = f_u_arrmul12_fa5_10_y1 | f_u_arrmul12_fa5_10_y3;
  assign f_u_arrmul12_and6_10_a_6 = a_6;
  assign f_u_arrmul12_and6_10_b_10 = b_10;
  assign f_u_arrmul12_and6_10_y0 = f_u_arrmul12_and6_10_a_6 & f_u_arrmul12_and6_10_b_10;
  assign f_u_arrmul12_fa6_10_f_u_arrmul12_and6_10_y0 = f_u_arrmul12_and6_10_y0;
  assign f_u_arrmul12_fa6_10_f_u_arrmul12_fa7_9_y2 = f_u_arrmul12_fa7_9_y2;
  assign f_u_arrmul12_fa6_10_f_u_arrmul12_fa5_10_y4 = f_u_arrmul12_fa5_10_y4;
  assign f_u_arrmul12_fa6_10_y0 = f_u_arrmul12_fa6_10_f_u_arrmul12_and6_10_y0 ^ f_u_arrmul12_fa6_10_f_u_arrmul12_fa7_9_y2;
  assign f_u_arrmul12_fa6_10_y1 = f_u_arrmul12_fa6_10_f_u_arrmul12_and6_10_y0 & f_u_arrmul12_fa6_10_f_u_arrmul12_fa7_9_y2;
  assign f_u_arrmul12_fa6_10_y2 = f_u_arrmul12_fa6_10_y0 ^ f_u_arrmul12_fa6_10_f_u_arrmul12_fa5_10_y4;
  assign f_u_arrmul12_fa6_10_y3 = f_u_arrmul12_fa6_10_y0 & f_u_arrmul12_fa6_10_f_u_arrmul12_fa5_10_y4;
  assign f_u_arrmul12_fa6_10_y4 = f_u_arrmul12_fa6_10_y1 | f_u_arrmul12_fa6_10_y3;
  assign f_u_arrmul12_and7_10_a_7 = a_7;
  assign f_u_arrmul12_and7_10_b_10 = b_10;
  assign f_u_arrmul12_and7_10_y0 = f_u_arrmul12_and7_10_a_7 & f_u_arrmul12_and7_10_b_10;
  assign f_u_arrmul12_fa7_10_f_u_arrmul12_and7_10_y0 = f_u_arrmul12_and7_10_y0;
  assign f_u_arrmul12_fa7_10_f_u_arrmul12_fa8_9_y2 = f_u_arrmul12_fa8_9_y2;
  assign f_u_arrmul12_fa7_10_f_u_arrmul12_fa6_10_y4 = f_u_arrmul12_fa6_10_y4;
  assign f_u_arrmul12_fa7_10_y0 = f_u_arrmul12_fa7_10_f_u_arrmul12_and7_10_y0 ^ f_u_arrmul12_fa7_10_f_u_arrmul12_fa8_9_y2;
  assign f_u_arrmul12_fa7_10_y1 = f_u_arrmul12_fa7_10_f_u_arrmul12_and7_10_y0 & f_u_arrmul12_fa7_10_f_u_arrmul12_fa8_9_y2;
  assign f_u_arrmul12_fa7_10_y2 = f_u_arrmul12_fa7_10_y0 ^ f_u_arrmul12_fa7_10_f_u_arrmul12_fa6_10_y4;
  assign f_u_arrmul12_fa7_10_y3 = f_u_arrmul12_fa7_10_y0 & f_u_arrmul12_fa7_10_f_u_arrmul12_fa6_10_y4;
  assign f_u_arrmul12_fa7_10_y4 = f_u_arrmul12_fa7_10_y1 | f_u_arrmul12_fa7_10_y3;
  assign f_u_arrmul12_and8_10_a_8 = a_8;
  assign f_u_arrmul12_and8_10_b_10 = b_10;
  assign f_u_arrmul12_and8_10_y0 = f_u_arrmul12_and8_10_a_8 & f_u_arrmul12_and8_10_b_10;
  assign f_u_arrmul12_fa8_10_f_u_arrmul12_and8_10_y0 = f_u_arrmul12_and8_10_y0;
  assign f_u_arrmul12_fa8_10_f_u_arrmul12_fa9_9_y2 = f_u_arrmul12_fa9_9_y2;
  assign f_u_arrmul12_fa8_10_f_u_arrmul12_fa7_10_y4 = f_u_arrmul12_fa7_10_y4;
  assign f_u_arrmul12_fa8_10_y0 = f_u_arrmul12_fa8_10_f_u_arrmul12_and8_10_y0 ^ f_u_arrmul12_fa8_10_f_u_arrmul12_fa9_9_y2;
  assign f_u_arrmul12_fa8_10_y1 = f_u_arrmul12_fa8_10_f_u_arrmul12_and8_10_y0 & f_u_arrmul12_fa8_10_f_u_arrmul12_fa9_9_y2;
  assign f_u_arrmul12_fa8_10_y2 = f_u_arrmul12_fa8_10_y0 ^ f_u_arrmul12_fa8_10_f_u_arrmul12_fa7_10_y4;
  assign f_u_arrmul12_fa8_10_y3 = f_u_arrmul12_fa8_10_y0 & f_u_arrmul12_fa8_10_f_u_arrmul12_fa7_10_y4;
  assign f_u_arrmul12_fa8_10_y4 = f_u_arrmul12_fa8_10_y1 | f_u_arrmul12_fa8_10_y3;
  assign f_u_arrmul12_and9_10_a_9 = a_9;
  assign f_u_arrmul12_and9_10_b_10 = b_10;
  assign f_u_arrmul12_and9_10_y0 = f_u_arrmul12_and9_10_a_9 & f_u_arrmul12_and9_10_b_10;
  assign f_u_arrmul12_fa9_10_f_u_arrmul12_and9_10_y0 = f_u_arrmul12_and9_10_y0;
  assign f_u_arrmul12_fa9_10_f_u_arrmul12_fa10_9_y2 = f_u_arrmul12_fa10_9_y2;
  assign f_u_arrmul12_fa9_10_f_u_arrmul12_fa8_10_y4 = f_u_arrmul12_fa8_10_y4;
  assign f_u_arrmul12_fa9_10_y0 = f_u_arrmul12_fa9_10_f_u_arrmul12_and9_10_y0 ^ f_u_arrmul12_fa9_10_f_u_arrmul12_fa10_9_y2;
  assign f_u_arrmul12_fa9_10_y1 = f_u_arrmul12_fa9_10_f_u_arrmul12_and9_10_y0 & f_u_arrmul12_fa9_10_f_u_arrmul12_fa10_9_y2;
  assign f_u_arrmul12_fa9_10_y2 = f_u_arrmul12_fa9_10_y0 ^ f_u_arrmul12_fa9_10_f_u_arrmul12_fa8_10_y4;
  assign f_u_arrmul12_fa9_10_y3 = f_u_arrmul12_fa9_10_y0 & f_u_arrmul12_fa9_10_f_u_arrmul12_fa8_10_y4;
  assign f_u_arrmul12_fa9_10_y4 = f_u_arrmul12_fa9_10_y1 | f_u_arrmul12_fa9_10_y3;
  assign f_u_arrmul12_and10_10_a_10 = a_10;
  assign f_u_arrmul12_and10_10_b_10 = b_10;
  assign f_u_arrmul12_and10_10_y0 = f_u_arrmul12_and10_10_a_10 & f_u_arrmul12_and10_10_b_10;
  assign f_u_arrmul12_fa10_10_f_u_arrmul12_and10_10_y0 = f_u_arrmul12_and10_10_y0;
  assign f_u_arrmul12_fa10_10_f_u_arrmul12_fa11_9_y2 = f_u_arrmul12_fa11_9_y2;
  assign f_u_arrmul12_fa10_10_f_u_arrmul12_fa9_10_y4 = f_u_arrmul12_fa9_10_y4;
  assign f_u_arrmul12_fa10_10_y0 = f_u_arrmul12_fa10_10_f_u_arrmul12_and10_10_y0 ^ f_u_arrmul12_fa10_10_f_u_arrmul12_fa11_9_y2;
  assign f_u_arrmul12_fa10_10_y1 = f_u_arrmul12_fa10_10_f_u_arrmul12_and10_10_y0 & f_u_arrmul12_fa10_10_f_u_arrmul12_fa11_9_y2;
  assign f_u_arrmul12_fa10_10_y2 = f_u_arrmul12_fa10_10_y0 ^ f_u_arrmul12_fa10_10_f_u_arrmul12_fa9_10_y4;
  assign f_u_arrmul12_fa10_10_y3 = f_u_arrmul12_fa10_10_y0 & f_u_arrmul12_fa10_10_f_u_arrmul12_fa9_10_y4;
  assign f_u_arrmul12_fa10_10_y4 = f_u_arrmul12_fa10_10_y1 | f_u_arrmul12_fa10_10_y3;
  assign f_u_arrmul12_and11_10_a_11 = a_11;
  assign f_u_arrmul12_and11_10_b_10 = b_10;
  assign f_u_arrmul12_and11_10_y0 = f_u_arrmul12_and11_10_a_11 & f_u_arrmul12_and11_10_b_10;
  assign f_u_arrmul12_fa11_10_f_u_arrmul12_and11_10_y0 = f_u_arrmul12_and11_10_y0;
  assign f_u_arrmul12_fa11_10_f_u_arrmul12_fa11_9_y4 = f_u_arrmul12_fa11_9_y4;
  assign f_u_arrmul12_fa11_10_f_u_arrmul12_fa10_10_y4 = f_u_arrmul12_fa10_10_y4;
  assign f_u_arrmul12_fa11_10_y0 = f_u_arrmul12_fa11_10_f_u_arrmul12_and11_10_y0 ^ f_u_arrmul12_fa11_10_f_u_arrmul12_fa11_9_y4;
  assign f_u_arrmul12_fa11_10_y1 = f_u_arrmul12_fa11_10_f_u_arrmul12_and11_10_y0 & f_u_arrmul12_fa11_10_f_u_arrmul12_fa11_9_y4;
  assign f_u_arrmul12_fa11_10_y2 = f_u_arrmul12_fa11_10_y0 ^ f_u_arrmul12_fa11_10_f_u_arrmul12_fa10_10_y4;
  assign f_u_arrmul12_fa11_10_y3 = f_u_arrmul12_fa11_10_y0 & f_u_arrmul12_fa11_10_f_u_arrmul12_fa10_10_y4;
  assign f_u_arrmul12_fa11_10_y4 = f_u_arrmul12_fa11_10_y1 | f_u_arrmul12_fa11_10_y3;
  assign f_u_arrmul12_and0_11_a_0 = a_0;
  assign f_u_arrmul12_and0_11_b_11 = b_11;
  assign f_u_arrmul12_and0_11_y0 = f_u_arrmul12_and0_11_a_0 & f_u_arrmul12_and0_11_b_11;
  assign f_u_arrmul12_ha0_11_f_u_arrmul12_and0_11_y0 = f_u_arrmul12_and0_11_y0;
  assign f_u_arrmul12_ha0_11_f_u_arrmul12_fa1_10_y2 = f_u_arrmul12_fa1_10_y2;
  assign f_u_arrmul12_ha0_11_y0 = f_u_arrmul12_ha0_11_f_u_arrmul12_and0_11_y0 ^ f_u_arrmul12_ha0_11_f_u_arrmul12_fa1_10_y2;
  assign f_u_arrmul12_ha0_11_y1 = f_u_arrmul12_ha0_11_f_u_arrmul12_and0_11_y0 & f_u_arrmul12_ha0_11_f_u_arrmul12_fa1_10_y2;
  assign f_u_arrmul12_and1_11_a_1 = a_1;
  assign f_u_arrmul12_and1_11_b_11 = b_11;
  assign f_u_arrmul12_and1_11_y0 = f_u_arrmul12_and1_11_a_1 & f_u_arrmul12_and1_11_b_11;
  assign f_u_arrmul12_fa1_11_f_u_arrmul12_and1_11_y0 = f_u_arrmul12_and1_11_y0;
  assign f_u_arrmul12_fa1_11_f_u_arrmul12_fa2_10_y2 = f_u_arrmul12_fa2_10_y2;
  assign f_u_arrmul12_fa1_11_f_u_arrmul12_ha0_11_y1 = f_u_arrmul12_ha0_11_y1;
  assign f_u_arrmul12_fa1_11_y0 = f_u_arrmul12_fa1_11_f_u_arrmul12_and1_11_y0 ^ f_u_arrmul12_fa1_11_f_u_arrmul12_fa2_10_y2;
  assign f_u_arrmul12_fa1_11_y1 = f_u_arrmul12_fa1_11_f_u_arrmul12_and1_11_y0 & f_u_arrmul12_fa1_11_f_u_arrmul12_fa2_10_y2;
  assign f_u_arrmul12_fa1_11_y2 = f_u_arrmul12_fa1_11_y0 ^ f_u_arrmul12_fa1_11_f_u_arrmul12_ha0_11_y1;
  assign f_u_arrmul12_fa1_11_y3 = f_u_arrmul12_fa1_11_y0 & f_u_arrmul12_fa1_11_f_u_arrmul12_ha0_11_y1;
  assign f_u_arrmul12_fa1_11_y4 = f_u_arrmul12_fa1_11_y1 | f_u_arrmul12_fa1_11_y3;
  assign f_u_arrmul12_and2_11_a_2 = a_2;
  assign f_u_arrmul12_and2_11_b_11 = b_11;
  assign f_u_arrmul12_and2_11_y0 = f_u_arrmul12_and2_11_a_2 & f_u_arrmul12_and2_11_b_11;
  assign f_u_arrmul12_fa2_11_f_u_arrmul12_and2_11_y0 = f_u_arrmul12_and2_11_y0;
  assign f_u_arrmul12_fa2_11_f_u_arrmul12_fa3_10_y2 = f_u_arrmul12_fa3_10_y2;
  assign f_u_arrmul12_fa2_11_f_u_arrmul12_fa1_11_y4 = f_u_arrmul12_fa1_11_y4;
  assign f_u_arrmul12_fa2_11_y0 = f_u_arrmul12_fa2_11_f_u_arrmul12_and2_11_y0 ^ f_u_arrmul12_fa2_11_f_u_arrmul12_fa3_10_y2;
  assign f_u_arrmul12_fa2_11_y1 = f_u_arrmul12_fa2_11_f_u_arrmul12_and2_11_y0 & f_u_arrmul12_fa2_11_f_u_arrmul12_fa3_10_y2;
  assign f_u_arrmul12_fa2_11_y2 = f_u_arrmul12_fa2_11_y0 ^ f_u_arrmul12_fa2_11_f_u_arrmul12_fa1_11_y4;
  assign f_u_arrmul12_fa2_11_y3 = f_u_arrmul12_fa2_11_y0 & f_u_arrmul12_fa2_11_f_u_arrmul12_fa1_11_y4;
  assign f_u_arrmul12_fa2_11_y4 = f_u_arrmul12_fa2_11_y1 | f_u_arrmul12_fa2_11_y3;
  assign f_u_arrmul12_and3_11_a_3 = a_3;
  assign f_u_arrmul12_and3_11_b_11 = b_11;
  assign f_u_arrmul12_and3_11_y0 = f_u_arrmul12_and3_11_a_3 & f_u_arrmul12_and3_11_b_11;
  assign f_u_arrmul12_fa3_11_f_u_arrmul12_and3_11_y0 = f_u_arrmul12_and3_11_y0;
  assign f_u_arrmul12_fa3_11_f_u_arrmul12_fa4_10_y2 = f_u_arrmul12_fa4_10_y2;
  assign f_u_arrmul12_fa3_11_f_u_arrmul12_fa2_11_y4 = f_u_arrmul12_fa2_11_y4;
  assign f_u_arrmul12_fa3_11_y0 = f_u_arrmul12_fa3_11_f_u_arrmul12_and3_11_y0 ^ f_u_arrmul12_fa3_11_f_u_arrmul12_fa4_10_y2;
  assign f_u_arrmul12_fa3_11_y1 = f_u_arrmul12_fa3_11_f_u_arrmul12_and3_11_y0 & f_u_arrmul12_fa3_11_f_u_arrmul12_fa4_10_y2;
  assign f_u_arrmul12_fa3_11_y2 = f_u_arrmul12_fa3_11_y0 ^ f_u_arrmul12_fa3_11_f_u_arrmul12_fa2_11_y4;
  assign f_u_arrmul12_fa3_11_y3 = f_u_arrmul12_fa3_11_y0 & f_u_arrmul12_fa3_11_f_u_arrmul12_fa2_11_y4;
  assign f_u_arrmul12_fa3_11_y4 = f_u_arrmul12_fa3_11_y1 | f_u_arrmul12_fa3_11_y3;
  assign f_u_arrmul12_and4_11_a_4 = a_4;
  assign f_u_arrmul12_and4_11_b_11 = b_11;
  assign f_u_arrmul12_and4_11_y0 = f_u_arrmul12_and4_11_a_4 & f_u_arrmul12_and4_11_b_11;
  assign f_u_arrmul12_fa4_11_f_u_arrmul12_and4_11_y0 = f_u_arrmul12_and4_11_y0;
  assign f_u_arrmul12_fa4_11_f_u_arrmul12_fa5_10_y2 = f_u_arrmul12_fa5_10_y2;
  assign f_u_arrmul12_fa4_11_f_u_arrmul12_fa3_11_y4 = f_u_arrmul12_fa3_11_y4;
  assign f_u_arrmul12_fa4_11_y0 = f_u_arrmul12_fa4_11_f_u_arrmul12_and4_11_y0 ^ f_u_arrmul12_fa4_11_f_u_arrmul12_fa5_10_y2;
  assign f_u_arrmul12_fa4_11_y1 = f_u_arrmul12_fa4_11_f_u_arrmul12_and4_11_y0 & f_u_arrmul12_fa4_11_f_u_arrmul12_fa5_10_y2;
  assign f_u_arrmul12_fa4_11_y2 = f_u_arrmul12_fa4_11_y0 ^ f_u_arrmul12_fa4_11_f_u_arrmul12_fa3_11_y4;
  assign f_u_arrmul12_fa4_11_y3 = f_u_arrmul12_fa4_11_y0 & f_u_arrmul12_fa4_11_f_u_arrmul12_fa3_11_y4;
  assign f_u_arrmul12_fa4_11_y4 = f_u_arrmul12_fa4_11_y1 | f_u_arrmul12_fa4_11_y3;
  assign f_u_arrmul12_and5_11_a_5 = a_5;
  assign f_u_arrmul12_and5_11_b_11 = b_11;
  assign f_u_arrmul12_and5_11_y0 = f_u_arrmul12_and5_11_a_5 & f_u_arrmul12_and5_11_b_11;
  assign f_u_arrmul12_fa5_11_f_u_arrmul12_and5_11_y0 = f_u_arrmul12_and5_11_y0;
  assign f_u_arrmul12_fa5_11_f_u_arrmul12_fa6_10_y2 = f_u_arrmul12_fa6_10_y2;
  assign f_u_arrmul12_fa5_11_f_u_arrmul12_fa4_11_y4 = f_u_arrmul12_fa4_11_y4;
  assign f_u_arrmul12_fa5_11_y0 = f_u_arrmul12_fa5_11_f_u_arrmul12_and5_11_y0 ^ f_u_arrmul12_fa5_11_f_u_arrmul12_fa6_10_y2;
  assign f_u_arrmul12_fa5_11_y1 = f_u_arrmul12_fa5_11_f_u_arrmul12_and5_11_y0 & f_u_arrmul12_fa5_11_f_u_arrmul12_fa6_10_y2;
  assign f_u_arrmul12_fa5_11_y2 = f_u_arrmul12_fa5_11_y0 ^ f_u_arrmul12_fa5_11_f_u_arrmul12_fa4_11_y4;
  assign f_u_arrmul12_fa5_11_y3 = f_u_arrmul12_fa5_11_y0 & f_u_arrmul12_fa5_11_f_u_arrmul12_fa4_11_y4;
  assign f_u_arrmul12_fa5_11_y4 = f_u_arrmul12_fa5_11_y1 | f_u_arrmul12_fa5_11_y3;
  assign f_u_arrmul12_and6_11_a_6 = a_6;
  assign f_u_arrmul12_and6_11_b_11 = b_11;
  assign f_u_arrmul12_and6_11_y0 = f_u_arrmul12_and6_11_a_6 & f_u_arrmul12_and6_11_b_11;
  assign f_u_arrmul12_fa6_11_f_u_arrmul12_and6_11_y0 = f_u_arrmul12_and6_11_y0;
  assign f_u_arrmul12_fa6_11_f_u_arrmul12_fa7_10_y2 = f_u_arrmul12_fa7_10_y2;
  assign f_u_arrmul12_fa6_11_f_u_arrmul12_fa5_11_y4 = f_u_arrmul12_fa5_11_y4;
  assign f_u_arrmul12_fa6_11_y0 = f_u_arrmul12_fa6_11_f_u_arrmul12_and6_11_y0 ^ f_u_arrmul12_fa6_11_f_u_arrmul12_fa7_10_y2;
  assign f_u_arrmul12_fa6_11_y1 = f_u_arrmul12_fa6_11_f_u_arrmul12_and6_11_y0 & f_u_arrmul12_fa6_11_f_u_arrmul12_fa7_10_y2;
  assign f_u_arrmul12_fa6_11_y2 = f_u_arrmul12_fa6_11_y0 ^ f_u_arrmul12_fa6_11_f_u_arrmul12_fa5_11_y4;
  assign f_u_arrmul12_fa6_11_y3 = f_u_arrmul12_fa6_11_y0 & f_u_arrmul12_fa6_11_f_u_arrmul12_fa5_11_y4;
  assign f_u_arrmul12_fa6_11_y4 = f_u_arrmul12_fa6_11_y1 | f_u_arrmul12_fa6_11_y3;
  assign f_u_arrmul12_and7_11_a_7 = a_7;
  assign f_u_arrmul12_and7_11_b_11 = b_11;
  assign f_u_arrmul12_and7_11_y0 = f_u_arrmul12_and7_11_a_7 & f_u_arrmul12_and7_11_b_11;
  assign f_u_arrmul12_fa7_11_f_u_arrmul12_and7_11_y0 = f_u_arrmul12_and7_11_y0;
  assign f_u_arrmul12_fa7_11_f_u_arrmul12_fa8_10_y2 = f_u_arrmul12_fa8_10_y2;
  assign f_u_arrmul12_fa7_11_f_u_arrmul12_fa6_11_y4 = f_u_arrmul12_fa6_11_y4;
  assign f_u_arrmul12_fa7_11_y0 = f_u_arrmul12_fa7_11_f_u_arrmul12_and7_11_y0 ^ f_u_arrmul12_fa7_11_f_u_arrmul12_fa8_10_y2;
  assign f_u_arrmul12_fa7_11_y1 = f_u_arrmul12_fa7_11_f_u_arrmul12_and7_11_y0 & f_u_arrmul12_fa7_11_f_u_arrmul12_fa8_10_y2;
  assign f_u_arrmul12_fa7_11_y2 = f_u_arrmul12_fa7_11_y0 ^ f_u_arrmul12_fa7_11_f_u_arrmul12_fa6_11_y4;
  assign f_u_arrmul12_fa7_11_y3 = f_u_arrmul12_fa7_11_y0 & f_u_arrmul12_fa7_11_f_u_arrmul12_fa6_11_y4;
  assign f_u_arrmul12_fa7_11_y4 = f_u_arrmul12_fa7_11_y1 | f_u_arrmul12_fa7_11_y3;
  assign f_u_arrmul12_and8_11_a_8 = a_8;
  assign f_u_arrmul12_and8_11_b_11 = b_11;
  assign f_u_arrmul12_and8_11_y0 = f_u_arrmul12_and8_11_a_8 & f_u_arrmul12_and8_11_b_11;
  assign f_u_arrmul12_fa8_11_f_u_arrmul12_and8_11_y0 = f_u_arrmul12_and8_11_y0;
  assign f_u_arrmul12_fa8_11_f_u_arrmul12_fa9_10_y2 = f_u_arrmul12_fa9_10_y2;
  assign f_u_arrmul12_fa8_11_f_u_arrmul12_fa7_11_y4 = f_u_arrmul12_fa7_11_y4;
  assign f_u_arrmul12_fa8_11_y0 = f_u_arrmul12_fa8_11_f_u_arrmul12_and8_11_y0 ^ f_u_arrmul12_fa8_11_f_u_arrmul12_fa9_10_y2;
  assign f_u_arrmul12_fa8_11_y1 = f_u_arrmul12_fa8_11_f_u_arrmul12_and8_11_y0 & f_u_arrmul12_fa8_11_f_u_arrmul12_fa9_10_y2;
  assign f_u_arrmul12_fa8_11_y2 = f_u_arrmul12_fa8_11_y0 ^ f_u_arrmul12_fa8_11_f_u_arrmul12_fa7_11_y4;
  assign f_u_arrmul12_fa8_11_y3 = f_u_arrmul12_fa8_11_y0 & f_u_arrmul12_fa8_11_f_u_arrmul12_fa7_11_y4;
  assign f_u_arrmul12_fa8_11_y4 = f_u_arrmul12_fa8_11_y1 | f_u_arrmul12_fa8_11_y3;
  assign f_u_arrmul12_and9_11_a_9 = a_9;
  assign f_u_arrmul12_and9_11_b_11 = b_11;
  assign f_u_arrmul12_and9_11_y0 = f_u_arrmul12_and9_11_a_9 & f_u_arrmul12_and9_11_b_11;
  assign f_u_arrmul12_fa9_11_f_u_arrmul12_and9_11_y0 = f_u_arrmul12_and9_11_y0;
  assign f_u_arrmul12_fa9_11_f_u_arrmul12_fa10_10_y2 = f_u_arrmul12_fa10_10_y2;
  assign f_u_arrmul12_fa9_11_f_u_arrmul12_fa8_11_y4 = f_u_arrmul12_fa8_11_y4;
  assign f_u_arrmul12_fa9_11_y0 = f_u_arrmul12_fa9_11_f_u_arrmul12_and9_11_y0 ^ f_u_arrmul12_fa9_11_f_u_arrmul12_fa10_10_y2;
  assign f_u_arrmul12_fa9_11_y1 = f_u_arrmul12_fa9_11_f_u_arrmul12_and9_11_y0 & f_u_arrmul12_fa9_11_f_u_arrmul12_fa10_10_y2;
  assign f_u_arrmul12_fa9_11_y2 = f_u_arrmul12_fa9_11_y0 ^ f_u_arrmul12_fa9_11_f_u_arrmul12_fa8_11_y4;
  assign f_u_arrmul12_fa9_11_y3 = f_u_arrmul12_fa9_11_y0 & f_u_arrmul12_fa9_11_f_u_arrmul12_fa8_11_y4;
  assign f_u_arrmul12_fa9_11_y4 = f_u_arrmul12_fa9_11_y1 | f_u_arrmul12_fa9_11_y3;
  assign f_u_arrmul12_and10_11_a_10 = a_10;
  assign f_u_arrmul12_and10_11_b_11 = b_11;
  assign f_u_arrmul12_and10_11_y0 = f_u_arrmul12_and10_11_a_10 & f_u_arrmul12_and10_11_b_11;
  assign f_u_arrmul12_fa10_11_f_u_arrmul12_and10_11_y0 = f_u_arrmul12_and10_11_y0;
  assign f_u_arrmul12_fa10_11_f_u_arrmul12_fa11_10_y2 = f_u_arrmul12_fa11_10_y2;
  assign f_u_arrmul12_fa10_11_f_u_arrmul12_fa9_11_y4 = f_u_arrmul12_fa9_11_y4;
  assign f_u_arrmul12_fa10_11_y0 = f_u_arrmul12_fa10_11_f_u_arrmul12_and10_11_y0 ^ f_u_arrmul12_fa10_11_f_u_arrmul12_fa11_10_y2;
  assign f_u_arrmul12_fa10_11_y1 = f_u_arrmul12_fa10_11_f_u_arrmul12_and10_11_y0 & f_u_arrmul12_fa10_11_f_u_arrmul12_fa11_10_y2;
  assign f_u_arrmul12_fa10_11_y2 = f_u_arrmul12_fa10_11_y0 ^ f_u_arrmul12_fa10_11_f_u_arrmul12_fa9_11_y4;
  assign f_u_arrmul12_fa10_11_y3 = f_u_arrmul12_fa10_11_y0 & f_u_arrmul12_fa10_11_f_u_arrmul12_fa9_11_y4;
  assign f_u_arrmul12_fa10_11_y4 = f_u_arrmul12_fa10_11_y1 | f_u_arrmul12_fa10_11_y3;
  assign f_u_arrmul12_and11_11_a_11 = a_11;
  assign f_u_arrmul12_and11_11_b_11 = b_11;
  assign f_u_arrmul12_and11_11_y0 = f_u_arrmul12_and11_11_a_11 & f_u_arrmul12_and11_11_b_11;
  assign f_u_arrmul12_fa11_11_f_u_arrmul12_and11_11_y0 = f_u_arrmul12_and11_11_y0;
  assign f_u_arrmul12_fa11_11_f_u_arrmul12_fa11_10_y4 = f_u_arrmul12_fa11_10_y4;
  assign f_u_arrmul12_fa11_11_f_u_arrmul12_fa10_11_y4 = f_u_arrmul12_fa10_11_y4;
  assign f_u_arrmul12_fa11_11_y0 = f_u_arrmul12_fa11_11_f_u_arrmul12_and11_11_y0 ^ f_u_arrmul12_fa11_11_f_u_arrmul12_fa11_10_y4;
  assign f_u_arrmul12_fa11_11_y1 = f_u_arrmul12_fa11_11_f_u_arrmul12_and11_11_y0 & f_u_arrmul12_fa11_11_f_u_arrmul12_fa11_10_y4;
  assign f_u_arrmul12_fa11_11_y2 = f_u_arrmul12_fa11_11_y0 ^ f_u_arrmul12_fa11_11_f_u_arrmul12_fa10_11_y4;
  assign f_u_arrmul12_fa11_11_y3 = f_u_arrmul12_fa11_11_y0 & f_u_arrmul12_fa11_11_f_u_arrmul12_fa10_11_y4;
  assign f_u_arrmul12_fa11_11_y4 = f_u_arrmul12_fa11_11_y1 | f_u_arrmul12_fa11_11_y3;

  assign out[0] = f_u_arrmul12_and0_0_y0;
  assign out[1] = f_u_arrmul12_ha0_1_y0;
  assign out[2] = f_u_arrmul12_ha0_2_y0;
  assign out[3] = f_u_arrmul12_ha0_3_y0;
  assign out[4] = f_u_arrmul12_ha0_4_y0;
  assign out[5] = f_u_arrmul12_ha0_5_y0;
  assign out[6] = f_u_arrmul12_ha0_6_y0;
  assign out[7] = f_u_arrmul12_ha0_7_y0;
  assign out[8] = f_u_arrmul12_ha0_8_y0;
  assign out[9] = f_u_arrmul12_ha0_9_y0;
  assign out[10] = f_u_arrmul12_ha0_10_y0;
  assign out[11] = f_u_arrmul12_ha0_11_y0;
  assign out[12] = f_u_arrmul12_fa1_11_y2;
  assign out[13] = f_u_arrmul12_fa2_11_y2;
  assign out[14] = f_u_arrmul12_fa3_11_y2;
  assign out[15] = f_u_arrmul12_fa4_11_y2;
  assign out[16] = f_u_arrmul12_fa5_11_y2;
  assign out[17] = f_u_arrmul12_fa6_11_y2;
  assign out[18] = f_u_arrmul12_fa7_11_y2;
  assign out[19] = f_u_arrmul12_fa8_11_y2;
  assign out[20] = f_u_arrmul12_fa9_11_y2;
  assign out[21] = f_u_arrmul12_fa10_11_y2;
  assign out[22] = f_u_arrmul12_fa11_11_y2;
  assign out[23] = f_u_arrmul12_fa11_11_y4;
endmodule