module or_gate(input a, input b, output or_gate);
  assign or_gate = a | b;
endmodule