module xor_gate(input a, input b, output xor_gate);
  assign xor_gate = a ^ b;
endmodule