module u_rca4(input [3:0] a, input [3:0] b, output [4:0] u_rca4_out);
  wire u_rca4_ha_xor0;
  wire u_rca4_ha_and0;
  wire u_rca4_fa1_xor0;
  wire u_rca4_fa1_and0;
  wire u_rca4_fa1_xor1;
  wire u_rca4_fa1_and1;
  wire u_rca4_fa1_or0;
  wire u_rca4_fa2_xor0;
  wire u_rca4_fa2_and0;
  wire u_rca4_fa2_xor1;
  wire u_rca4_fa2_and1;
  wire u_rca4_fa2_or0;
  wire u_rca4_fa3_xor0;
  wire u_rca4_fa3_and0;
  wire u_rca4_fa3_xor1;
  wire u_rca4_fa3_and1;
  wire u_rca4_fa3_or0;

  assign u_rca4_ha_xor0 = a[0] ^ b[0];
  assign u_rca4_ha_and0 = a[0] & b[0];
  assign u_rca4_fa1_xor0 = a[1] ^ b[1];
  assign u_rca4_fa1_and0 = a[1] & b[1];
  assign u_rca4_fa1_xor1 = u_rca4_fa1_xor0 ^ u_rca4_ha_and0;
  assign u_rca4_fa1_and1 = u_rca4_fa1_xor0 & u_rca4_ha_and0;
  assign u_rca4_fa1_or0 = u_rca4_fa1_and0 | u_rca4_fa1_and1;
  assign u_rca4_fa2_xor0 = a[2] ^ b[2];
  assign u_rca4_fa2_and0 = a[2] & b[2];
  assign u_rca4_fa2_xor1 = u_rca4_fa2_xor0 ^ u_rca4_fa1_or0;
  assign u_rca4_fa2_and1 = u_rca4_fa2_xor0 & u_rca4_fa1_or0;
  assign u_rca4_fa2_or0 = u_rca4_fa2_and0 | u_rca4_fa2_and1;
  assign u_rca4_fa3_xor0 = a[3] ^ b[3];
  assign u_rca4_fa3_and0 = a[3] & b[3];
  assign u_rca4_fa3_xor1 = u_rca4_fa3_xor0 ^ u_rca4_fa2_or0;
  assign u_rca4_fa3_and1 = u_rca4_fa3_xor0 & u_rca4_fa2_or0;
  assign u_rca4_fa3_or0 = u_rca4_fa3_and0 | u_rca4_fa3_and1;

  assign u_rca4_out[0] = u_rca4_ha_xor0;
  assign u_rca4_out[1] = u_rca4_fa1_xor1;
  assign u_rca4_out[2] = u_rca4_fa2_xor1;
  assign u_rca4_out[3] = u_rca4_fa3_xor1;
  assign u_rca4_out[4] = u_rca4_fa3_or0;
endmodule