module _not_gate(input _a, output _y0);
  assign _y0 =  ~_a;
endmodule